`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iMNrs/xGUapAQqnTpsnLPCXUJ51ycUqRibMxluSlWyB4sGVAcCp/ILcZQfgi+JhR2CNq48kyZX1L
mH/vf7Kprg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
H7Z3IB1v3drLp3rDBCLqQjQmFK6J4MRSgGqazHH7W1T71FHW+dZ/CBfsCeP6t/uw1+viCHeYpiHx
Ts0hK/qUX+An4SPp4kqE46H6ObKf9crqnnGOhxhng1dPdEUKSsk/8MHfmqpT03zFHLoUEzGAihye
3amKH29QDLPcCRkaLBw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J+pPV7pcY4Frgq3lWOlY9UHMtz5gA+vrh6UEYfQgFMw/5FMP+YkKz6SNUgSIvfeoyO7C/N8YwIHt
o510Zx+PTek07+e6HG5/SAugUDEN9T0O4Dc+gNlTEcx9xxoppkRigIMOWaTn1qiaqCFBzkIqjiwt
AqIL4jv53/jaxlNn56cIn49CyVZoiw3Sca4HJoppPdpfWxxpehoVrM11UlnWXWPDoVmnaihVAsqt
XrhrYbHbd/eGhvyZ+YA3MoBVdKb12qcPEoiSUxt10/i37LMPNk3zeJNksedA+MxwR6VDDnPPctBI
8VIYG26fh9c+2yro989k49Yxv8UnMbJp/aTx8Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zOyj522533FuS4Dhk8EUvy8HWZPAcGO72EdDgsNS9UbFW7UcT7F2oT35Gtlmy3ZJWkJ+PsGoQIxn
MaSVerZMjOxGPmhLx1rUWk2CkTxjonEuoM+GL1zTeSaL/bajGb+SyXfh2XjYNqL8DTy6eQaJsO3a
BesrzIGgRt6J5OsfRSg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kPXbYUW0nftXjyLFl8kOO+siwO2qim0AenLBtzM7kBzb98F6JQYWX4WPpVsWnySQFapPpyUPgPgd
b41JJGid7kQU3QSuH5nxgCj7a5k8Zjg+6hfpM9eHrCluIHZWYYZ40B6kctSXOFA/EdIruSavnNTK
BNa3wU1BrF3Xxe/3+pOUbVhiVpEAqtEogWNb5u6vuRJTDU8KMOmfyGpNGlDqT37UZrO++ljGkc2q
1rVIXufoYQIi/E4ACedXsZraxPnY773JmwAhumUzg9DsvPM9jhOc69eUhR7OmSvdzSVSMwcm9O8N
HEetPWFYKG5KpJaeOjrP3YrPUAndtYADpefBfQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HeONVLbck70+T3lUDee+OJI3960XbNMkfPLjCjAIeJEQUNGjYdy2cTx8TK5gFIm1Szw7lYhxL2E9
YbrqbEsord1TReD53Kw6IZbGcc4QtQ5weq0gv6AWLIBjMw1m/qtENMRyh+DaJYaZRvbG39WqwSv9
RKdyxcegQjSx0Wi9Mkw5ukKUO1SNBlzYjZZoCNQrh7K1KFjCs5o+icQwipAdSx3UEX++1/NPTSsr
z+uZW+pfTKM2BwcOcvUXBstmUIi/8loExiVnke9pDvlKyTCB/1onLpaA2jRpuUE62vHJcTz9m32n
uh5OTObd4uPX8Mi2u5vV+Q/TsdiI86XA8c8evA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13632)
`protect data_block
m31p4DvPR0Op1Hr3mLHwzfsD73KREP/fJkbLzTxgfb68WDLCagDoUVoClZYF7HCu+9MppRWvanHn
nNoLoxJ6FG4PvtUyX7xJiXcIBQR8PQhzcTEZg9Lf+cWumFS3791mUYunHkaR1NzDetOV9Ixv0xNM
ubPBPwAmeDZ5AWC+RZ/nfRWQzMoWmypoOO9WnwbtE98dh85fARs581uimWdgYkLX5AFqhOFC5bap
QSBvXuJbAtD2OzySaukKZsHmNJR61v2q/GfSClokq/jf8M02W19X2pVjaZFlOy5Kph4D4ePPjLq8
mkE6x1pErtJAfXA9OZV9y6/AOJs5450yT+FQA1aHir5f/fl9WToi2dbKloCkZNyAPDiLY/yaFIKw
b5e/ed+Rm9sF4d5s9ffcrf0ugw7Fm77CFiCuhK0Jgdyea39kVEASb2KvvtX/zKQiahuVtNsKyaZe
f/QtmMQVUMbqgSJ4HyqNaJkjpbGqLLwuiorUI9klpQ91RKyVBvomDx5rany/O8C1tEnI1Qs5L2Y8
jAcOZmU086p7h+RUu1d2B/hqrvObpnmJL2l7eag1GjveS1rRLcRp+OAmn+PBhqALQ6hk2XDttiXV
DoiwzD1vg5YyjZvopsxbkcMe3JuRKhqqVw1lIYHywho68cRICGXF6VLm3WaSH+KbJ1h7Fvubs2gf
t045TuFOjUzusXxx6j9sXBi/0qXayNRf5kc4p5fMgDZC1znjdMYMXxGRflufonV8V8miheoCFIHs
NpKivtEQC05rYqJFEFHmCAY71VLs7+/kTi7BLJ8+60sin43mD0ThGn9ahG/w3+J/gZlPuouW1YDt
DnZKWNMgM9MAd0aXJupWecow9vFa3qus0vypBssHrhRCvMJ9Un4R0xJK1WJ9ja8tkDHuEKkrlut3
FP0b4CMS4F27fBTmnQ/NXHcrRHM9tkZXpzBwLOO2QBbgWv6IE7Xk67KpwEM21AZPQxQR0sLPpo0g
ASVog4gXtGXmYnQleyZLiO69UEZ/aQexXLxcU0C5N9DnxFiGAeg58wAQJv0YeNYvCfPsVPkCLVWJ
05mCR3aonq4OuVnWDuzK23h/DqdRKmUlGAC0qsRjvHdYmAHlyzDFSLI3lFnfSm5+mcmuOge1RFRG
ZQsuEmYeXA4iQ8gkI6Q/Vrh32d3koJMkTNxs1b/dlmsi22Pcx3yTsGb38LtxAeQG9THIH/JLnn4i
n0BsUN1qokTwsAOdYACCB24BXBquZ9jvkK+kklvH63gDyXMX1/MbFWB1pBzzPX4exEWQ6vzPX5wr
oaAZ8nspDZTDb2uhe4Dj3lBWPinPYusqXNsW0mHMTdFThEL5MlnxIqPRHfobZjsihAw2jQahQRNn
bzYWL1Mb/6ig/AOG8jcO/OPT8GnDcU9na9r3Anhwb+7gzzUluAn40bo3Sq+dd159GMhhahzyN8G0
SIcpU1kR0ci5DJi+9ENQ4g5mh/SyJB8yJ/Xp7KDa4mthq7jzktVnPOEsdJ8qejzsSgouKZIskkH9
9gdMew2BZQAoq0vW3APaa1sRFGnjYzmbQ6ctvkTV5Jifhx98iEJFBQe+ZjRTLQ9y/CTvlvf5Wahn
H+ffEFu81GYE3Lnb/92mVmNXaUo0uDbaiv5anq8t9JbtGf9bQplgLmu9rr8ED2o/VjRUT4GtEzOR
GC3nDCeDCMvWJLnvml0lolD/qQdyPiLfiFbpBSZPUw4dFiZjnCRp7EOJqXLKP5UjkPXSW6ej2p3f
UZ6iGuIEvajThAhdfr1fWI7BPngEp32fzu44O0/K9BKpOQH6oiwfttycqGGoNbzCHoTkHwdvnaCb
d6OJ7Y3ap5YMP5WaX0Wqvqu+PJ8M4bNIGxwLbwkEyIuOHrzuTvLHHiYpPmv+1GeFdl0AqOY1gKer
sj8JaqTuAs3kmxOfSpuB7e8Sd4TVCrxYCHZlQZtByWQqMRjB1fP7lDssdkHMp9rOhEoejFKz9brf
imujI4qBjMjfQLY+a5ELsWOmOeg+A9Wyp6fnpff9Xhz8vFhw48M3HCFlKvDyPrBA6Nambjni3ZUi
3I6L+F4rntNZpdvkw4t4zU7FPbTJqYTAE16ExsExpTKX1f7Pckcz+T8AowconBL/c4NirAR7m7fR
LSNbt/n6e0nRk5yZq/7zDS1hqbpUOi7ro4zd+TGnAs00dvrIZSjf5Ylw6sHnQcm9YX++Ig8P8Gli
YDBjm6UhDatdlTx07pfNmsqcbQO5rOAi86mHjVg6MU5rZnrY2OVHEvwfeKtZFd4IfjNR+Ef7tAAO
6bXuINkDQSGdqkIJrMTGS3CPx1FdhWuCjibI706/bQHvX2cIkMpcqCiIN/C6CxZSoUZzEV5Fv67j
gkFORCGtrTXRtbY4gvzSprUv7e0Hk2sgHVL/q3AFNd+lq3aL73IXeydn1IBAfEzZ0z3BgGa/fdun
tpgUb37lfegDOCiUCxMZLnAoPnCVKy8nGImJWgbIJ90vuOIUIAma0iJHQcZI6wywsbBqOdWDW6Us
VM1hfm+w1ETpkMuFqUc08kxlQG0CsEBx2RA+NA1FHghRNLs8xWhIMMkRO2yx71vCt1p1+qPThm/z
SH76zk6AQze+Hhlj0Hf0FAONz9iKODGRcFWTnrkPMzeYtG3JVF1ajpxdEYbJmk4fzt8Ll3g7ilZo
dbVQJsQdC8FNz1Lvcr8V3pPop6V+IegRg9wfmVYd04X+ZR0KW96C0nnbCW08mKSUQJ4JFbP0AA7v
XZiJACxJQtC8UZScZN1GdW6cadFqmxsLCI3Z9Eta3JdIYjfKZ/Scnrv44m1Kz04KHkyYCyXWwkUb
lksmYD41k7nMDa+lvojU41tsBAWruZf2P+zhHFY9VcznqRw16/3gvYcO2eIs8XDu3fxDMPWv1z2o
4/vAS5fn5/GNMHRoGT1tTiOQcJS33d/g4zVcjz1rE8Q8JYSle4YTWsbz7h6zKDnu6zm4M17Z3iie
wY9kjonMzJEEhb/lAonJhMCL9herCpYdSEib3FHjZSTg4suyUvemn7YS/feHli8F059s9J3rJ8dT
/w1YNf/Xb+F+OCIvh+HZFWSp8KsDNanYznPpPVNXqvoR4ZWbnY8iN+r4X2JtVa0fKpFsTFZwE4Wh
r3xGTCxY8QVQs5VfdRWhYbp6PyAsSOi5nTt5+rNNdhJQMFPlkE48wkJvk9pV5bgUrXpKN0ApFGCd
cxsLRPKcR6F2/9eCE/c75pwc6V8ngF4SQWH0i0XNEl6Kbd5WfkFvZl2RZA6RpdD7MQbVYEGT95p6
mgpx341n+StwkY8IjEN53rEOGDtbVz9l3krC55l5dawUlzjDvz1U4ixevoYTceYClHHR+T4r76S+
twTo/Gzz5Ml62MYtaAlBgQMJ7Fot5gC0DID+f1nZnhfnpsaXjKwiAXVJ0zk6NHPmHGNJXPH2xW5x
F4wCnY/eeiZvhZty/X4wDwBCdhBwfCc4owWgDQP1Th2GDsSJIW7JiSTv4E5+qjHsYJ9J4VcB8tsv
yMeigu4VqZnvIwvJHDiEa3uPh/+fgZEnm+L3Q3I8d5Z9Rp9awq5XpP4RBCescsO5x1YL1FRZ4L2v
OqP9f8pjGb5oKevszstgznUCTmxL4WWzZqt+pkg1Ighubwp3rrluMkf+rpD/s/kB/jvhgb3I81ko
YPwa6gSQe/gCmM2wI0+/OQO40Ov3ixaFe1XwKL5duin21zQKeyFtt24Q9g3rHAF967H+vuF3QiSu
L0d1oAvyIwkGIkePerMdiI7zTyhyqDyNX6uoCoOLgykKW1pW3aN/MHoKFMqpg5yih7bWXXrOLQMT
p8u703SgFoaAKfVQOCUmC2fbT6IVb1Lmw+LqxLBu0Zh2ZOTUbG4VW/F6OL9PlqbyFYTOvaoWfoaV
tca2BVqY6e6dCgqDibC7I8WKorRzg0D8JAfEg1a0t7d5KpXOp8WoH2qGiAB4tKRpxmWTtHb2vR9T
INycPWihaLqihW8Umys8GhyvwHbyNrK1Wv3nFNA7WMuuE8wICRdnWDNO5TVQ/MPB3CwILEyX7E65
oQpMZ9/7DsAOVUvuDKEi/1pHrEzSgj6X5MtjxEOYyqg5YBEMlHOviodsZSduLJ3PK0ckah7Ahv+w
eOxE+K5LRttRVvFizsH2JsympU/S/zcXwHFU5GppTB5JpG8L3+S695J1Z0kvkyC/2neMypMmG8bn
qUzOzcHi2CNxV5nqlf7k/iGhGdmNgRTskn80ba3UnairsVthsJAOLQeuZX4tFmm2qbLh6vrtpo+X
EipIdy51k9oPjsfDlP3YwNVJc65t/6cKRykGfCJ0ku8fAGSY59/zffXpULwBa96cXPvWl767OqPY
42uKamu1tncbpOCYjP8DxerNLDRhoLfPnAkBcg1H7j1c2psXRPiD9MPv3peRNd/gN9sQBLMLORDQ
XviOVgScnIoKl2N1cIpQSt/84Xd+2H4H+FN/XPBzONPKq6okvcHK0UaArK8g72c3XlQhja+p/vlo
ANpahlmTingyfUGbK64Fw7iT9k81T+1n9mAJ3CfM+XNNkIpUt4n6UJpKQMZi4LRB4vgImZQnAlZs
21KWY0K0lIkFC69LyO/YT6V7f7Ud/NE0h0p94i3PmRlYmsgviRcwPhybM99t7W8gDdIu2ebSN8Q9
Biu4dJcJyWVJXJ18a6CNaTaQQVdF5T5QHv1N4OAYIvFEQyi4f4lCh79EnhAx7FvVFlr1v84yXum1
XJb6gddw9qlmNAVQA/3AzI/lgEFzjngs7dPfQJqx4tI8DWYL9EUtEnE/vrdt7Jh6x3IAfevM0vrw
7IINGJmZuAzsSnB/zDpJtlMl8BprpCp/SPh91VxWBRLvh294ag0agzmKXohiNGwVvb9CVeHiO/sK
ag2nNMXGMAkKbfU/d8q32BYDZtccFWHsINAvt/fJgeWWE67KLufuL8qrUEjFRq4MMHmv3eBoWDOw
yaGO7rqcYbFQCWlvWX9wXXYQ0o37GpzENUvyhRw6LGbGwhv0zWO5ExL8rnTvQAm/xLpUG5XNNW3A
2DLFDmr7d6VKgKMZaxi9Ov99l40GbhG1G6kC+t3cSdSP5fyhvdC9q5iYygiHFcQxr9yT8o0ThC9F
liaIt/JUs2GxFJZ4XR1EDrd6j3WUOQkAWiBswLu5MKqK1Dstlib3OCIwlsnAW66C7GBXbEPGDbzp
koLP19cBryzTj8bi6hkvM0CT4OPJrKFsqA8cx0FLeJ7jFUH75HzuuY4NgtYIV0afOUWLt6pdQ+33
Vq03pAmYKRqb939qyOJgr9UqkKYKQ8suehAN0VUh6x4hw3nZpz0qatI95OkgSg6PPdgppnUPgADB
91HyUgvYkasabSRy6sGr+H4g/tyGwC0XJakyUjKVE/8D68iYA++ja+DUfRqqLK9cvsyPZPwyJsLn
vXSXzb872IVxvPUMq6ipn7ZqoUKL6SvrN7gG9OSNPC7qv3rgNmf/o5pFI4skqXmULLgOJLmBTZea
xGgMwvQVKhfBA0NA5i6hfHthoVDkNpD40F8PT4+q7W4gBmlGkRei+PfMrtXX6x/ruJ1flXqJNIjZ
By3y5wI2w2ssTIPCV5+CLfSxzY1fimvY7Xclfo2+Dch9Moq6rrruI0ODIqXqbDVCXjU41HcPATep
We3jUGlikhLXbAZmLV2xtvsNi+W/+Q8qHBoKbCgeJLLVnZL73D0nspKs4Iq3j1RjiJ1d0mDLpdXL
Zav4EI4AxIZIrUQAqrApINMeexfI+tPqud/eK+mWn1dWQLnOM76yDF9G6nxgf2f64kf6T3WRzotG
OQwkhgYYrBRFbN/lxlsO3PAvxyoQJn7YpahN8Mo3bdRnadGxXXoQ27u98lkRsbU48cSX2p9suk3A
5NlEtjrTxUPYgHmLd6qYrLU+/ALzywdK9cK3pZueadDrhCEqhiB4InB8TBXkxndVVc3JwJtWqsIW
HmQ36btFDMt4mdK79hIEJLK2kLM7Mf74JEAAq3Fp7mLuojEOXYyID4Kzs11R9G4/BouK6cG5eAC0
b7ONC8RTXMMjPBbGRPQwhIwhzpnCnpC0LdF2KIGrs/KOf9K45zl3Ij1vhd0eSf80ranhzlO2SM1p
BgOsv1IjTUET3CYzlTVrVaNMC+c2zLxMANh7j1X9U11SijerN+N9agmRICE4xfTnA7E2lhyH8nyC
TrqtHPRyXXBkqf8d5nMxAa78Po7QqodTkUamF+CD6dw1ueqCDma0w96PVusuPDr+LdoF1zPmOHU2
AOGS3mFTmJCg+XPl2C22atWHyM4BC58D6HsKeVIA7bytFGqNkEDQ04cUyvifyp3crOU0xgV22CoA
X58kQl5ATQnz+J5nAaHDQFY/UcEi+H/046JcxBCwarydkBtE5UJyEGA2aVVTWHcqwKll+w91L8Vh
9nrHy6ToZ3AohtFsB8yff68uDff7b96sphVlJWKbJ3xpxpMEGGPbyr9W/TvsNv+uzA2jGYTz9evr
wnPtMLPMQPNW1jte4lgUYdjteSKqQoFS4BtwtnH1d7BLrkGRYSpDPHdc2fj105evlyWvL8f4oWvw
A9/VrswEE3jceD+mOGEeALXrSvNkU8T5QjBqfAo9x2vFVTgz4rkuHM/de2UIKJJutO/vbfMxgxeA
+VNHaBnoiLbkp5kLLQJvAKfownZ4+KNm7LWMIdHQ2xGZ57Sa0seukABFL/HeRUqJLz8oV1pmmHNN
tMqmKNzMlbkVO5KO+86oUKYaJR0o70eESIL8k5fpt8RfOqyIel/vQ7+aL2YouagJvlMnMIPfNYiZ
FJRnSse74MOh2PUxYtv7S5sS0/XMn0/+KoSjDhKa3adByGiJ/VrUmo38SkgjH1NdydzKZZir0Uz0
ANBc0DwVwEcotKZirkTUA5uhKiNnflEZTweoevW16gSW0vSeSJrR8cOA2XdmwGcqOwq9KfEUFiFj
YcwQzvYezqBwW/nuQRFhl6gCaIA3S0jwMZ8OOoHcP4YtlEtk7zvCBViuANkxzJi0wCxfYT7zCEDo
LQzpVo5VBHNwDfzbUO2+kwsvwilecg29wpcALzRld35I7TU98ZJJ0DPhXQPgfbdrYdIJo8EQNkt2
qx9mwTk8ny1xJduzoaZhS7qJs7gZMW9pzbdDtjSN5qT+++s2+ysPhCR0YVSvbVpqeRtkeGx1OEyr
z8ZLAMUG3e7q54OhR9zPMmdIBwBegcwg5hMT2kBtnnz8s1b/BGHRK23tY8aR6/MKCqs5c6EZMugZ
KFUXACcY7SyUxCk1OVDMO3dxn9/fTRdSEEObmKyeX2jOjgWqbMVrMP0WdIbyYAwSL6C3FXieCFTx
J2qqqOA97QjLZr6rrnvPymRxAKIAEVInhObu8rdiLxYludQcGxQSSb/pmbGvpgsnaaw5mkCcN2Y9
PLgt5q1u+n9ew0U9ObPhC2pYuY0Z00a+IsGwP1DGC6fmmveZBGdCsFhB1gf2NDnj8qynps8sAtUY
Y3NUBm1FeAy6JOJdwEWj3d5cr7T7bYoCIqFnSxNBOvUiE+kZz7kGJIKhA61TC+KSc14w/DepuTei
G9UdcaXWIdI/FcGT8Y4k+iRgsXkiY6OA3MYOD12QHHJmNUywVKAHeR5oBEB+cJUPmM5E+qyRipSc
WOkCJK8bKleK/aoMrpZxHwKW8t+FRNb4sRhgqPFNbPCXEyw7owW37ukciPcJi72jNwMxkSifrToB
MQ+BYvOoCakROAFp11EuGukyK9+Rxxrp+0hSaQJrWX64u4siEKjPhIa+bu5xeVdvNxYnj74R2oRc
1u+jRzFBeHxUXoIhQNV+aiUBLCnkIjSdbDvVgR4XWEXJ9JT/W+AZ4sVeCPRSnvunUfnkTzXSfQSi
GsV3MfH4fjxn6Zgx3XqEse/MByNvQDCMwY4YoYQ2YTNyvcQHWrqCNN2vzjx0sbiHc5JzMegPPKZH
v/alg3Uj2VjR6+UNRNfHOlRFmOER5X6M2mi1ShmSYKQSH3CCUL8yMHMdAaJHujlTdEynUMt9nhGF
5iCzk01I5H90nZHZYsJm+EL66ZDhAHUtq7pgPDhisQjpZWfrLu9gajY32M8yB8xRp4/wonejSsNZ
J3Z9QDzIEggddFx57fqo+EneLVgzYvWCsPorOAQD/EpdcknNmlpEoV+HcZfP4BhuzAtgUX6K4q3u
+plJ+4r8QTdA1rBH/TQZcAXKBhKk4eOrQ0WZKjN/1hUW14b1A3RyBEUjYvWI9lc95h6vyHoCtfDG
Bfsbai5+0MSXYzq5NAGnY9cQLfH+lPfVm3Pb1uNJzIZke2t7BWRpk79+fDlqItRvIO/59A+gevhx
YwfSoMR8yx7pf1L6bE7TfbIv15rYojLztxgqINkmhZPNpIrjWeqkpHFIiPlSCZcBh6aktC/y2gI3
/J3zk26Kponcu2bOgIPDgGN3svleae+pdU5RvJH4opsTqgq5LUS2fJoiEnGnQGspPC3yHwJeQ+N1
WAzoSbwtiUlsFkw8Qz2tm9Fndt5dhcLYSu3AxG2YxKWtvg/ZzpnEJ0BUNa8U442j1Xo+YSU1VCoD
L0YnrHuMR+0AYZvoM15uLI27M6nwa21rskDePJ3koXmGw/kAUCV9kln+JPN/Tfeca8i8PqZEoqXD
uCjxveTTmYGhx7pmFTLYDXWP+s8ig+8MuaNw7eSudSBrg+3cQlhZMmG0Hl+4YWUHkU4iFgVLmJPA
d5/TJ2o3b8j+prSdQZYn7nWFNxH4A8Ev7+AkQn9MUAl8Clc39qFdEg+4mAO/swSanM0VT3Iu76yi
grnlbdfyu0U8WM3ezXeRe+qLdVPA/Jv7jp1JUSJO0RkUV9s1cEenZ0xibPfFq9s/+zwMKyiF6FR7
o2rM0cxTCf2flcPMhZhG1We/B73TAYuM8Llh6zIepCowu66pAq8iGTMHxRJgMeJg84R2vyCL2lI/
VZ/p3ps0urQECGFitSxNT3ugTV7y7Tdq+JTkAkUlXCrEtBliMnJKQ9WJ3VzyB4mPI1rNAX3qxtfC
s8GN+GXG4x/fjX2kY5R2EJHKW1/TWwmYDHCG9tAMI1b2x1k40IX9WAWNJ+EvLiw2AEY8ANXw74F6
BIzx18cthpZm4VLTu+7p5KuPX+eGv6iLCGXAlvZSqbTJeBIB2F/+EB1Y522j3K+A2It90pKScONw
6sDDxh8jlTMh4ZkuJgsxwT7eObvYr2WlkPDoL/vhkHs9RXRN2gEP+MxB1uPaMmXjEIQ9yhVPepg2
7R7K9YyDkIHltVc1fJl36mLABBlrhObN8M7Hwgt8vdvddbAw7ZDo/Ftt53zmHXQ5bCzaccPxRPIp
QZ5MHIfHovx8euwbzZb88fxS+NDfyWfnvBMN1HSlVSuCeLbHBk5w9zOl3q/GGhjwpFHo4BP1K/j/
xfh5NAUIo6Q5CeQy2AL0Wk1l5AB2BfchqHKBZ0HA0aQhavEpVhjpSp36fH/M0oZ+Dxg+7rFsF3rS
FLF7zCjDU7CYoq6gxT39msyuHQY7n33tmNk+tACjQ5HU68re2UihbkI0Dsnv1lRkKIxnPto5LQj1
2hUQLVMVGFHMpf7RxgFYbDo961whFwAhEoEmM8ZhUBJf1Me2XGC6rpw7+W1s9Dd7D88xIPazvbdX
TWDxYuDQOmdjGj5p0k7DvKxbVGseWJanuP+2QxPUUeH6h94mRKwy4QuvOGh+D3XXDFl4FVY8B6A9
O0jJG2eRzoHVjAuHSaH11J9ORartv/J7R6s1WGTvlbDcJ0kbI0TBsQ55upIt3dPQ4SDaPxVzEJ5q
tgCJNjugs0yk7F6xpdVEb8tI/vzBqZ8H7jPZ18fE3jAT374kQ3nxcsmBog8SIQ2gl6BRteMZfwDH
c4skhvIja1caVwqo+ZN/KVObuAXJ8fv61elG47Ws/2B3pQn7GTzPDOkWEDUEQ/n3Ti8cuTK+lj4D
JxDZfu1JkRJDGKzKgVE1qZGpbIpKoy/WiycOl+sCXqpYdjEBR1Kb+podS7PWKXOhfxXMH/2+rk1z
OLlB1h8X2LbTHcenKkUFBDm+oV9NDmB1rX057C3ukHrTpDkyxZuUc8Ec/wLve+NnKmYPJHDdrhUG
5vdhFyAl/gCWj4Y0Enl66HCw7YPWNeOTs3zh2L0FnFY7NLnm18dYMuzcP/8QqKshmpIJ/e2uz7uD
DRChMbcrxepGKNmRhRhOVCcq4gZAXble8tNJi8ciBj4t49L6lfCtX1n4Yn1CJzvCloqdxJBeb8dG
ZIB2KmLvlGjTiYs3NK2HC6RUaaahZhmoRC1I44acwUvrIuhbqo9gS9fg1+/ZbYktjxYkBNXNd9MR
Ph68mQtir1DkPCPa2Z5HTq6ChIoze5W5G2m4JgRg4SvWcHL4QhEsAob4PQGT3dnVTWZ/njAQ2ReG
47dCA8+MxuFJSPFKs1k8s6GsBQ5AcjVQ1dTcZG+9vxN6RXF3qBITZ1ZD1gWMCVu9c1sKwza4rAyD
Np/lCvzmG6ZIjlWXXce6veBx+Bql1cl0hrrBNkpEVVgMFa/5D/B8XAPY3bSOvjP1pFZU/ip9Fh8l
jjhL+TmWHpsWBTfs/TVvepZ0MpUEj5DM14F8RI5KXmNIBtzkH6L+8g4pbIhd4zbi8StAm3Qk/A7c
nElQ/ueOC9BCtycV5tDJA1Sg/ZZyW/F2MAYp+qcqdmxYZVV0v6e019TeufFClzLlf5UA99fw+j6s
2wzFuwapPVImBIkW+ztXnjSA962ouNImmKbTjY36l3pK1TNZVUihXY1kZQK2cZIW2INfIPKz/j2J
V3ABMcOTPZUCMV3uRocS5R+EdwlYQMTjwWid/Ccl+P8JDxXSbbNO0YcTGw6xooldWMTsbYHThKPl
/Ai/bbKzJPCxvVPOglXU3A6HRoxqeGXH5tCsTT8WHF5Y8/QcT4mhcLL9nuP7NHFER5rsRmVbdlB3
pFou8faLQRGejzwJ5qEpNPLEIOYCY80JQ7X1hrHKpylghXipfPjcbtpFniSOnxlKQr8/C29G+/n+
F6SjwM3Cx+Mr/GldD6QZyNlpHsNtBQSpk+ujTSicMWrFRsWmMowqbEAERgphf8jMOJGezpcN9uwq
pBVSWMG74UXQhDT+gms+uoFl7k0I+WiWPWw9QXQHgw/8UMrUCNF4HCMhx1oHRaVbJv2PkEiDFw/x
vLg4en1GHNWnbUQawOgyAUh9UqPVs6W45RTBnqWT/HUdp1t1f18P3fRR6x5nu7aZIfAVGIJnqNxA
PevpqXBqt86e+836plrDgKJlgc6TUk/CYhkl26t2QkNuSyCsNtQeDaRfOKZ5tuPF+SqgjKOZtsyO
2hgVuIA6xS4+caizN5/llWcbQtVnPu87x/DE1rp42wt4MumhSFPRUQQ2P2Ik65jxpEc79kOppZvQ
Gb6iVL3IYDkVLIjei0/rjE2bM1jde6HkWWgZ5DB28QPcTZdXhA/uwFJA8CW05JL+2ImPO7Ei8w0F
Om2ywlLaIrnOucMc35jl3LO6iMKJjOCrEzBsw87d0AS4AUu+E6ZM5MqA0XdhtHxOsjzGIFZ11g/b
32S6i8UDGH/Ocb8f0HlsCbrkABYrV5NhOwnV2f9WamwcgF7KGkArp4+1cJTwzTSKL9RamMqRKijO
kNFXa81eXzIl2Il1l9OBe4tU5M0av39GtL9c4972kr+PnEEyo8l/FTtu7kB6n5RWkVZq/Hq00KA0
EEKXmawAH7reblt9FTrrgNnjwUt6U27ixrUGu+DcAXQlC7cWm4koOBFDQdSq43KUkKQ9WICVfR4Q
55DSUHxHNDM2XQlCEi8bby1BKx1EiBuY9bvfd9wXVyHs/tpmrlURZ+FrxnU+BnQxxnAPzr88qyQ4
RqNqLUqTlxzv7XJOCNmQ5NRrurh+6h4SnwS6IkEF976nno7v0GcEAn3anoCT/mDBmRG00EOJoBwX
diIGdyP3WL0u2KxfnTwoKGVjCLXB9NKR816X4Rl+MPU2ugLq0FvozAyWrvySs/N5xVdRfuR/sZct
55MSgDB7X4U5J/2YZ5mGBi5ntzroEDbat+DpImixWBsr0iE/73Np8OiCfdTAtq5JXJF3dmCB5e9W
6XXrOPW5NqsDgCdhohmDpvolonWJMvhjUAygnytGXx/AGKiPUhisnqUKvFJPUTUxKtqzaQUjYde9
SQg61cv4AqkcjtgZ1IFPImAKodb1sxYYlU0fv+WruvCdoVBNce/epkNk8HpTDfnJmQeMcT1mX+Qo
IaYli2SjpV4W9vPuBkHMv9pA9Ziae1oN1C6Ic/K+vIha2ZpVaYrC8rja0HU1pl6aMP6gn/zmGvRm
/FXxVhfmN6Cn2Vk40EPT6p2Km92L4/mv/9SEIpbG0zG+M682V7oRBfEZAvt6WVw62ZRIOhaoTni1
FMoPeikiXESNHXp5Ns6niRnhbZYfK869Ds8EYF9/H7zClPGidWHaWXL7T6Jn20WOE9ue2dVf2/LJ
PeoP6QRrH3aer+Vgfg+7XGB6rL/ruaOsuuwkafXBuUbE3Z1pSroDlEP+FKJl3K50RtfLmyxALD/k
RuWCq7AIacaQ6b6ddzE1SvtS8tx5RJw85q3avp0JSfpZUgF8CnIUd0hs/UrQfcwvoeN0+QCBiI2t
N+j3/E5Sr1gZ/MKwbjrrnjWO47UrSd9mmhraYrBauZidGisvYVvnxhJut26VkpmS02JdVCuSIMD7
hNs/U8+h0V2LCOIVtYrcNnAoW7khst7oOyYMf01j9pdgO9shfH7Utn8x1N0hwJ079c0MTqwPHoP3
Fa6FmUeqnRwMFMdNji6Wt35R25AEm1TME/hzxxTq+KaJ/AIk4efq9sjo/0YYknRfdoqASWWlYKUc
S0yOFyz52T0NmDVd/g/U75clwMeoR6Fyp2u7ZeScIWTfSSOlhD593Lxw97QapuPGKLEf83t+QDEG
bsgx9k6BNkyE34NqsebDCe6sRnudZlmdycBgk8bSrYbt8HPSH6ywR9eUSkhiwB1FeRD7/Ih+dNO6
jghEoY3IWfGm2W55n2+8leDf7XLMUn58P4huklYCR3WxU0xG66Sb+V+iGMh0UQPNVLzcEyvZTxeb
BPgTqL1totJVy4TCdWWsnoWLSyA88uFGBjwMKKfAdU05Ifwo9Yl56F+TPwIoEuhszq4tYKjEL167
8+e32fSoJltNKzgfQWJFk/t6YQvaENKTESj+2nbIh7wOGo3pQFOOooz8AX1OiKGsPAARVm8kvig3
cX06acOncSNxLwvkroxG81/is9tj5FErbcedXpbjWMAJHxXmr+GPtkasfU7vDjEB/2HFKQQZI8zf
oI4uIJhAgO8vBEy3ftRAdvhhf3G0JKApoNnOWbghx6INoEvkgKPodeshp5Axb2bW6t/DEwqmMsPS
kcNsQOVPeQR+ikDeNtyoYFF42GuXZIpEi0Ggd6Jh24JRjEAzqf74/IOEDJL9f5eNAMdDEnOVchlv
FeKD86cT07rYyL1uAm3N9fqB6hOAl3UNze3hHc31JuiW4KtSOFcbvnpE8ROCEhZX9rC3J7ZMp82J
+Y4sOli4VdCYo4/TKjVNO0iogXFm+RK1PgOO5HQ/6kzmvmtChy2FbG/7hlPLFiYuoom+23VMmz9O
+DZYP8modfB7kbSavwbQvLlA23zTOzv6hxtsusNT/ph43yfwXcQB4x/vtfy9Z7ilCB6iDm8KSwWm
KYuuzGSj3LZdardWxq/GNkOUCNZbv54h518lXznSkURcgtAj+XAuvF9gTRw7+LPCNwpjtToqcCYo
T/aUQtWKsIP4j+19/erskjTKEcKRiR4OVcBubWjghOr10RaGs+RPyx/61UIQlm5/efNggjJe5WDD
1YKXVhzdUTYjvZ0wg3n8WSje3VGloktFDW/2YodjrWMjdBgOj0bJuwM2DfY3eZtwp98gBsYm4+7J
a1yBHEekqrzidoTaB92rtemCcPpeKN/BbGdINkWuvAWoZr/p2R+zD99qZuAgt80nyD1gb+amnaJ/
aKuinYLrc+57y2x9h/7II4z6TycMAeO9rzuYSfA73uowkxWVHoryF+6u/8FJUz18zdryljNyZaNQ
gTAhMr72q+r+viV3se14vhZg8IM9XQQjBbm0GC+QJVodlfSBoV+QGyIoqlw2Jg7JYqvcmmMfFcR1
M2FN4kmtLhRX6PenIZgq2C8R1IqX6SYvEOoykYjqut194JXQlx9h2TIHeLewhGyWU3uaQx4D3fO3
XyEmG5xl3FdaVi4RBrf83UVZPcaOzdnmhuaRQ6fFbi+KsgSixyjtw442FiO0AKFjXY1yJoQgIqGJ
s7ljIiDgFGz6XDjRS0AWFL7BH2v+5JnrGAu/C8giIMiU3xzrK05gOKUg87aEYWMqAycQkTAnyuV0
c1/E4zTW+WYnA5oZtumaeE1zOXNK4B33ya5Drn5k6Pyrgr4jpQ4UgrN/niLo8UFct/IjG4a3L3tQ
kDbkTskvKKJNkk5WkGf6pkhNn3el4+cTQm7PeSpn9KWdvACbW2meuLVa6lu/hbLPbhE8NGxCAJnY
T6dFVx1ViW77nsWUmEJLaW5hMtDBZ8TvLs1FIUPaGysLw1mr45Q1M8JlMaiMpI3AQEgMckzQ94Ep
iwp7Hs2Wx2E8CcsoSUH3gJ4CvW97Dp3mo7abmymDGLbqsfJRQbq/VVanPz6zpOSL4TelM3JZIGBD
aiO4NwpqOX7nVoHfhELcGqwws5Idn21wUH1q60fcQrcu/L3HNzvnm9a1t32e29YBi4wZQWStBuqz
tY1XTNoecuB6y5qGjnyey/UJx8pAF08VVU/u6bD4BX4QB0u+Nt5WjjUKWqTQDO7i2XF4sESZVLoV
1nnF0Oj+PYX3FfZxImpJAmJqX2SqrI+4vgDfSeisVzxmiwUf+QQODRuePPdQHUMb25PjY2IZaX/5
We6ICYM5pxRZpRSU/NFWRY9oyOJepwzekwzd+/ORzd/XnVFx2hjo6KJDrpYFBR1SIIRm8Zy9bM1I
mafrYgZcrysl96S+/+zRMHBjQpoMplsh0GkmPDZdPqMpheHD2LpgMxocaPbzI4aWdIeQOrT8qhqg
ntzY6y88R0Qa9LF9tAIFvCJsATIuFbJhAQSnjuapLJDmWDeTH2z2O5tW8KH8AS8VwDRGEsZll1lq
yL/AMOqF7KSwCrkG2kZ0sT9nkC7ersZnNTrDPjLn9kpRp8uTVmFYadL3eJ6UCwRPiaOdeEmERUld
Yt1+WHVEAYTgvh4Xwvp+MD1ykCNm8xIBvP5VyDPNHr6vyUTI0+18oMltW0YnWrAR/GkDMkjNlj+N
cFhm6FfPzKTe143JscJjKXQISsJVmTZyIdm7TWSJBLjHNMKR/mZl/H5Eq3mTyKQLgHYcanKO53pD
9TBOHvERGHBOVd9+TyiCb9oEk0bIGoAG+63VEgKhrlAXxOAi2t9nTtmf84tv8XeoEnQPGSS5sGUQ
appxm9mahBQIRQwoiavjjPBxihn7xY/0BVair8nCQprArmH8A3lqDzk5poUrUEoC/dIhxVVkEGYL
lmWyIrFT7QlXVKceayIyerm3DY6pjOPr+9Zs+hk7wLqATkW4/3+4w1+UIPgZi4+AZzxmU0BPycLp
SBFjs8/emArhmvWsVrSslp2EBltpqkvLDDmKaxIFbxj1vskCHlAtUrEfb6x+FRSP+vVIkKtH4dkn
1l6/iMiqhOqDJSyO663tTJXbozCfhMi7YXSuTpcey6RInRIO6O1/VB1sMuH4wDJFFQsR4sd0t5cm
W7aXvfDDvhQwPG30nRWj99WXxPMNtC0bPX+gtojxbETqMf18Sta3YnTbXg8JMjQ54kMr6I6Ek4ej
mX2GlGSx0gniB+7WJdWpAsJrwJUNr5+Gljc+GM8rzjzKBXAXqlVXHe/xPNeM2YaC7W2v3hJ/BZ6R
vCWUk/Wpo2Laihc5tt5vJLkoYazActgFoBgjvdth50meKqiajgkkIDcZu+USDlYh4XFkXLjqJ7W/
EwgcrvXga7yHfA/44Jj/HMjRbiuZ9qtJXvQhqA3N7iLLEP8XA7ZrIAFU8FgaaFfVoFxw6lfsT14L
ciuP64br9H5u6GHHkxBfpGgVhlZ5RS/c2woPU9IqjO47jL5pUOqjZMyE9i6zP7nZnUxLWbDhd/Mo
/gGbubRW4ijqrATP4gWWvOpsBo479zbS3LSZnanHanWxkKh6/uabLr+tbQX0g7VDt4dL9sUdQw3u
HgQajh+8K5/DzCctor8K3cKZxeKSSg81fTqPQe8vUTMal6nq2hb3OwAD/RG3fG+4fSKLRZ92sh0m
wLEHkoV98VMHmbSDoj3YY6hnLcEfx2DC48O5HT9IdbKKEtMjXVeZ6uSv7/9E5F+gti1MazaRHvF0
pHQmwRYjr/SnUH1SQciCoJFqwQiDUFmvfrrLRNAJ1bh7+S9Vq91Z5QcmcC4ij2UNpTRB25dWB/gu
M4fuXbpwgoDy7L/zZsW44rcAtystfieWoNIDVxfdwu951MKHtag2aKv8NdWuK0vvfPITIRg+JFqv
98p4ZQEYL3KJ18WXnBhsw4cVbVX7iM+mxfC4tx4axZ0Sew/lkH3ScTieAcR9WTcjF3qxPFJ5gmy/
VOURchHkQOxbfwLmDoILiVjgCzodSfVu9LuuhmBkOQphLMHzEZ5LR0TNArYDVkcHcgTQfnR+intX
P5YdBdGHy8S/mRPSmKW7LeVM6cOrrwK4S3R6jQHJxY99xIYCIVyx53zmFhH+BKgaoI+9EW3Q3wSe
Jekt+WwiT6SM0kqfBxLnUjrZzlyCXVm4EvHc7nmYP5Exqkqs76Q3u5MgAqytnaLGUI+QN1RLqt+g
ay0Lrzqo3bnnEFI1ZuK1SJGf0z0SMCXHzFYSnJerL6MjFjtrei0U3+0dkMSTNdPd4nDAm+hO5N6N
3ky4BKafjmHhASdcF72YY4y0fNfl6TQzz5sXCpqw4yU6pKntklNMbAEFKWkPVjaGNCnyUMHacFOA
0pqqueGtmHfdDro+No+I5Z24nqpvYpwU3JvD/k6BuvzAM5CLul1Oi9sn7qNRc2wAXXSDWsLKe0PP
w7w2x0O7XhN6/ZlwNE0OvXRj2gRyv9SRlzkcp+DljSo/SgUX5lPVpCh3i2rCz8iZhSqxr+hTMFgC
GXbU8TmBtrQZcapq0iWqBuMTFTSNJirXvaUkJe1+nhaq4RGh633myxl5pWHKKbn1rCisMVeRKmmz
9roCdGD7Qp8iF8gTMW6yhdjgRPvx+BXRfksFBohpIoylT1zlvDHFrP9SP8NjiBWUoTtB6M67j0Bm
GrM995Y/dHRt06snR7DtiKB6xGIu/73TZRs0VJFXqzoNf/bZKrkfgUiMojZlT2hURF3P0pbYGTmY
sez4KtCebci/Gdy3DmcXEnOUJNTQFhMXY1+mIq09xhMSRXA00KkrCN56O7CMSnmlZic1gk5tnDrD
OxNj1ht6ZzoNdwAJFKqlkZH63n+nn/MEjMElhLtb4N2xUYRoAEPItSR8W/tNe6ItKD9gdZUIWUSs
wgSnV0OpWiiqtIBkgXCifRmNAS6oOzkBiZgWkmFssFmGQB1t8c7qSMjn0yohLVXaYLkJGHAb5n84
dlZ8YlfREo3roX9hgP3UufJP9PyeaXtWZevIATypP6MTPE7fV3WiSYd9IpAP2n6zpvlVwYl6leHi
Zy+kcoHzu/ZJFl6n5yPG90ntJWfEbJ/1O9rdBmOVh/LWJ2muzimtZyjJ9oX1ZoeES6D7CDdZQLzu
mx76mEqs62cPNYzFsRNjTheXrbx4QuVzWUlFO4VQCBf4LXqvPIqxU7YldQkb6zNA6eGNLsi0CHx5
PvhG70L8DmiwrRIMsg0PQzM3El3zSwW+Hq3cNX6s5mwMKfgJQYvEcShiyb1bpPib25jrjJxfrrzd
2h5DNQL1jph/in13sbaCnP5cSnSEc5PABy9Pd4BX9TCa19ng0KtXQueZhTmxa1FsIYnsBrt9ZHsS
JGw4DeZXc0Fp+ZjRWRet9+QIAQH1/hUDtx+4rYuugMD4RvGmI3d374SpthtlfRKMwLWPc1+L6Ew1
qN4br1M+Yz1rodzvbvfh+Z+a0Hb0Z+i7axCO0sKQozG9DOEGB2QuP5T/4IFTbyh70/0ehmiP8YCj
XDA24wvfdIjyIhWTu3sqZ1hxdGVKC/sVCaIMoFksk+6zrgqmrenwJWYQctQfJcphaSoiX/abyYAb
gf4aDe5S57HyLgPScC4ZzeS5TrlaEmLWFElVuj4lM15ca2p/H/y6bYMkCy9FUMyvl+eRhen71fsz
+bRQqy1TAwCC
`protect end_protected
