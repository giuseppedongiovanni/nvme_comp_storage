`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EIJPO9OSDMvMNdOLRjwQaF6UWoBQGuoL9zzQDGu35ZPwlaCEsuX2/bXZpi1PYJWx1fIV4fCHJ2uv
SGI9TaOoYQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jR96W/xy6IU1CwVZ4OWs9uQHbt8MxEY6OnhSFsNtb0hYTN1DbC1Q7k1rAopY5R85kliEBsNMYuT4
cKz3DR/nTb0Q1MQjXvFgtNYTIJn+x3l/oYgzda29/A8PpsBi6sz8KIglPS1mIVYa6RurRv4LkYKw
EaTHjYSLD9yqzkfqJaQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l+dRl/KQgn5YC8NdqXiuF3uROWLYUXnJ8JxZFU5L4rAPmX7kzGUXJZnRPvSDiahmvJuv8ANZs5gh
xs5LoEmDF0CFompV5QwULgbR2Q6qtwhrEPfg6MLWV0rRtc667uYFE9KTsFf9JZKKO4/H6DzzAdIP
WLVbf01tBroj4IeWcXlkzK/313rQETBKihcoZIo95c6hdiOI/cthsmWnNjsjRy0+PSU4464xZnC5
TEcE7sJSPGR/fWSbLVlBZxn3OEvlbOzvjiNR8+/H97sx/ei8Vj94gc3yWS1QgQO+AcvptL0n+FEy
JyLr8oQ6zAVfPaFj40vg/JebO/peHp+yKYPY5w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KHbON44TPSwtGlB38csZ+aUEMwCA8EA+f07XdNfbRNzHCWdzgmAoOb7uBfu7KxgTm9Dt8IjH0z68
A8EQUItPb1xEcce3WQRQmtBL+94WCLdFalg3R9madXc+OvDU9lJ30/cmMgJzC7ZqYcKNxsY+MltP
9DTs2k9PQ9HK8xPytpE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wBWhADcN+GmDp1YCpVhIm6ehHfqFBS6YvXzYJFLy6Hbtd4ICJ88jM6iQIHo3AmpIauawmkob48i5
njLAuUbhiO3pjbjswXm9m5ULq7P4Zl16GePbc8+NzBZSqwO0mIMB8wKnwW++E2Rn+Nns6sn6MC2x
zonzzsSzqRzajp9fUDbbOq2tS/NGomoy1+X36PLd7Cy5AliI6CDkRHdS0IOLAwKKtEXzMUbjOg7H
Dtr1NedDgP/xgl72/c9xLklOb+LA3hVkJJO16GJEccChdA/9ulSyPIsSQmXX2bub6jXFEifZQ/8t
ihBzhm2r0HZ75QWpj/gbGRQxM/9gTCkKkqLwzg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WEJsl//nwwFukI7AawNtPva4Okhp5BPPbpvcOrHU2WhmmE+kpe4aQOMO547NxOMlZwGZ/nioOZpi
LrmS2pTou7semtJjuwLmE1hUNq1JnXEjxFJO4V4nyJ54enCYSCvNZDfgVzETNMWgvh00LJlZjybK
m78e6vo4JdsWwhR2Egwd030HGF+WhpCBmJqVrWwK5tEGZIr/dG0JtSC4lyLT4TI0WhfArNiIuILg
4hItSA/a2fFSiFfuPJXYSodzb/CpnIKOqjTcK004JEGCZJcglHRpZxK5ieOzXEV5LQE3Ouc6ACbl
rwBw6NkW9ODG4U4PpNFnPhbwmmQLP3dpSXp4+A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 65248)
`protect data_block
bMfPX2R1tFs2k3nA+qlwsKoJziUZOwPs6DjXY9eXJxQc0uYM+CDAUpiUG6V+TMR2PH6ijTgCb6B7
pMdc5/pDtb2YVPqF9LhiTeT7x8zKqx0AuDMtUiYsaO9reuGcYhltSdOUxhRM5Oa7MwfI24R38I//
xvI73Y3knWzqvIm5U/S6lmzGiJZ6Jayeft38z0veeVMMJ63DPaqQtRaAqtYndrlmC6GSEc+hpdWc
2LC+hPSyC9dNUhKrbD5rxhyPaV5j8Todz1U/YupkRZ/4sxll4oDltMJjulXYkQS4qlLD5Y74KeI/
ABPQ1HgNly4+UW+GGXYxhFKF0JjzhFjoodO6TPOtOreYPGM6S+20QB0QlEAgzkYVXBO0ut/p50mt
Soy1FdD+oWDUvuSo0ldL8nqzLHHF8ZWo51wy5fPFh/gCbikqdhNqEOz+q0zjRqujbTUVoo2zgpBu
fZdR/eNYvw5ZLSUermVZY4myZxExq6hJh1rTTD+v8qT3vGXvwSiBgHbzEodsJNmfbptg1iMHSMf4
5AVJsOVrAlzpV9ZzmB4d64+JXONVZSg+Mc6jkSQRreA9NE9fraY29GpEvB9vIJoMXt7M5kPdkYIC
g3kMJA8Qd4vk9h98brUi3YS8mKx5ppPHxBCp6MatCsGORfc6tNYCHs7pOHq/ONSWkXEuDf6pLBd2
jgo//BwPE2WNOA7lrRQSKDJzOe2Iz7bfi5I4t4sOAluvG3zf7NRKvATgEFJGds4W1xJux7RQV+j5
kiLdcaKvSv1euLeJU7kpYaXDgMXVOLLRb9G8pHU/W6W2tnxMq8liGloYiHoHT18Fuy4AVM/nPh7g
+Z7dKIzBlU/w5SF+nzonQdFoQ6PFPuCm05sp9gxWNBQe4voN3YJPkSiAwKGxgJ8F2dWQWx6Io+b+
G8Q8hw7TIqDDwQYDFfYMTrbMuIc4V+zZFgmhRz9Wr+U+K536IDEcgd3dIQekZqxaG93XZdlK7Ubm
wlYMFlaLtk4YZ26f3Uw9Sn/o8tNQCOz1DC1fIA1ei7WgdjluHUTNUdKAXF3VXLQlZBcESr8EIeXq
7MzmtRoC8bqlAcXD5/px7KHtk+F+aU0DlM7yJUxKMKMXJBu7gooEIiLUx9tvU5NEP8dDPV9y13qA
Uz4LhTBFu6psVylxPp6B0ZdYEl8XJiBjInjIN+NGRl5rdkSGss7daIp2gybxPtRJorNvsGcMrtWx
Y2+T4Wymb9qlOAJR4DcWIIP0XqJCyAr+rNxxo+gZSfDlf/d7SfggUEAPA9ErxIRdnm4tRBBOdokr
3YyY5dGZeI3BPKflcu2PQ7BmfUOAY1tvB+2EDGCtnFsYi08Jm/2ZDlkjPlNxVml7MCtzPgn4qs7W
3mAuklTGH0AFQV+sD0f7pSAzX64xLlNk0tJRAwesIN4qzdK7SZIuPcSDBc3JUrPQ0myuXeGwoUC0
jjK2Sw2TR9bz/LaJMuvzeOtePSaLA69mw0bYI8UmqKe5ccbAiHt6dHhHog44yNv+BdP8HLpA98VA
BYzlDdYSL0LUlKXIij46M3uVTRdjCjXQZbOE+FFsIMl3Y5lLOvJdY1yBrQvKH3vlggMRtV0kor1A
nxZM9JzIYYp1y356Y6dFQMTnxbd643HeiIbbryF2DV61BQCimLAvxm8gDPSpInBy9um/CvCAONwe
fJetvjoTXBqedbkhw8g7PvmeZTttuQtFGI0CSmRZOcEkCNJcrtFSblgv7DG3zSUE9BO9vglORrcK
vNa6Zh86ssFR+tpT6p3J4C1t3uT/m9/CzGSdk8sZLcWH23KFRx/FHzmM0ZhHrWy4xPu3IOn0bbvG
b5uIPFMidWrto3kmtc4QvJsCvL9NYDRE/Pe2ss2W66H7VLSKqH8EtUWt9pUDNC09MPHkLxwdSODF
zjgwJpeaT1sZ6VTY1Tcb9YXq4xCl8MINYYyLgfJbhQln3z1Np12cAsFKvB+9mremDgzhbB2EkFxE
okW5fT/lFGwlVTY2E/es9WOw8wYrg7I5xFF8rQ1UicizFHZTrhSWYsRN6lKy8nhaw2emO2BOxnDz
olnwmFv5rb1gVHrDRRudJLO+IL0u4thKQSct2uDlupFz0JlGUsPPP3fZkiGAfMfeJy7J1G4jFpzY
BhAq0o211wlBF3cx9tM52o1XEkq8WjoMlbytpNAqjShJkfCKkAz6G3w4GVb49MPxWvIUgJM+Tar2
8yfCwXuCnin/ttlO+ydXnBrEv1EHka/Gl8ef3RPexlSFHmblncbdMirNikab+1S0Neb9fOOAqmUC
ec0U7VcwfL53PjH8UP2Eig2SgiLvUTno+i+MFg5SyjPUeuA8Qitze5k6PHJkXz5Pxu5hvStnrHwF
MjUpTpcOtkPT/0f/24H0Z1HF6sAppaykgRG6ZsbRXQ2041MAz4DFpp7axClWQe0SoCr7l6SgpOkk
t6vsHmO0lZAGTCMC8rNxo2eYwhT+9pbTRckdv9n/wsWtd5wSK4XrL/1McYSIZiWhLESACchVMmz4
dt1CBaYxkY6ISscLfGJUyJ6YFJee43nikI3MkEjhfDSiSiCtsvvp5t2Jyk22KVcP6bIGOXORtbYr
3NSLeHSZhZIogfUoaHEF4IfaWwLNFIUxzwUWyeQzZjSyCY921ssOKv5507Lod9CgiRVX5QCvwnOI
+Dg9GBzcQAWwRaWncBtAWtiztVWj2QjTADDrWhxUf+4kcpDfXWgTii0NKu+bX9TD9gPAwRH8W939
YS/McWr8rrpm5aJxx6J1tONIQ4NUAeOpGWZCi+lyvT7Pt9iV97Bs79mDEfn646KURgMukaADTxz3
nxpvpYt9WtFrXRgff6jL/sNEDSCgTBJzcqcuJCK152kdSZk86PozDboTZGheOfxR7jr3znxGVPNp
YzE4uubi1ENOYQOLVCx+TJjtUh3hA+T8iDJSvlmE8Nlqn7H7IrGnidyyriwVETRRTJKwtcGBZ8zu
3ywaDVk/EroSbExUk3JJyNcyO9ZQdw6GJUlycn8ynIjfN5TiOCrGMjpUPhlXlaBBUHU4MHwHFjlk
0AYsVc9VXDl0nkGnIDdD741rs/0w0Slbngey4F4coj44NvQay3qydaipA+SW8vL/b0AmItcjGGge
m42N3OUldtvQAXEy7KVKKbmN0QoJSK6S3qDd7U2YZtINxL/GHuWDQ9z8+f3evgaNU85iUb2FYVLq
1YA8XhEUepC8k8UKQVhbqandv2aMUloTbhsc+L9mZjStK4VQtaQ+ALdy3uHaSmlXyd4lh07mC8L8
I2SWPicAaUARfq6d4xSj4HE8HjyI5Kya/H+dUjkmzpHqzYHBjZXuKOnXtV6lSIuGk6vtwFvrCZF/
IjZkhwIcjUlgLzmyKxsvoqcRMctkBvcWNs6zm1hmSUPFytGo86Re1g483QwGCwfaCC8rHUgjKCfS
FCs/IkDqHXRBu8SVrbyvOUp/ye3NIKRjcFsV6B+gm/Tq2OtSsfGoXxJmJisMjwqNniIeEe6uss7S
nG3ulwK1n20FeoTqhs15wcElIlF1oIk/3eVJcL5aWJaZpQeh0Ld1BVr3a9FXz1sNmba0FWdDiyth
RRtqwSz3kMPgv1OAuRmkmpZpmIgHbbt5POI4+7L1kCNkTcBFdxwWny8KBLssZA7nuwD+XGIa4Vxc
AlawJS0kE/K5jIBoT551iF/HP5TQdXO28ErEWVTWFAUOfo9BfROl1CZ2SDW0G4aGqodrkh8te5fo
zNKjJNlCgR7OUwccQfaj1AbjxmLgtLQyok48nXQY6cPkiuZB9OvnW38bG6NSayVzJEeQhQO36pe9
kJm+Mwjz3fBjpudbffbJPdeBeh60WixOW6uawcfwSOm8tbP5gbgRmr6m/J8EuGyps+SxArdLBGuV
2BiMpwYRlrBBbwICM+i3GmCvxynj2usU1EQjA0uwfxEdeALtFsEkct4xkCxBBP1fX25UephbI3LZ
cP1IUGWEIbjWcEvFcJEBp59ddTuHWQbhbjJ4bth9fYuLrH81HN1RUjTZzoscBH6Y3hqbOsNG956b
r098iY0+vkftkKxeY/Cwg60ORC7uYupCy5meUMM1XKvbEOZB8gjgQmKCHndXF2HU/Xrom3dNeKaY
v/cpCRQi9AKegqscxwxsPKNg9OBugwmbjD90XVB61V9o+H96J3Cao7+AVG82egOh5i3TmRuxP/QK
UjDaF5LyP0Hjv6+wp1qAKSghUa0pvIxZc+J7/i1QnMaWq5bYYjdUP/ZT//VHYqOHJW/1gH4AdaxL
hd0ojcGxGqx1e89UX3/VgAy0g9Bo0b8FdVlofjJT0r41C39eOAecL528AgakP87lQWTnUAbg9T8b
SGEAeI/npZgdP9q7ZpvFlAzdvA6UsnzmBTZ++GDE1Msm8MEyAORgpuJYrv1dhPdtufqGVKp492sY
arcmeC5Mx4TzN3WcuQINL/VNLjlxUlv8JiMBuafJSb7Vp5L8k6YNa37BFC8y7UVXNade4b7zbHAS
5aTGiercV3gRBV83suee8RZ3tyu1Zdtvdw/j4M3byfpKExWSPbPnidwmn7ms0hagOUZ8+AFMbJsc
LVxaqFz1PHHyRm2kcUK+wTL/ySWfiSmmI80IeMRK7Cku5F1MJrl/ZfL6uw3TBeh8HPLkrfdYx5m/
YHForQFzn8ulI4NDhDJJ34z5Wjiy7storWYQcRopPp0D2TrXvRww6+sC4X2IkkVLa2Qw5fIOLFvf
hCHd85S5yks0qwCyZODBahxq4mlzKX6le9W67nKzQQbBeXWD6wiItSpgdyMiGDJCiVvbhAlk0phU
yJb9sj40zc1GgLidG5lpQMgjGXUVBDEmPseSLhr7JhokPB0kTgYSjOP6W28oyaVaGqarYOAElb/T
E2QGUQRxYDNgbFAiOvcUYTzKFnTTyUaEZLvmzVoQObvA7OUsbvVaMCMH8XdU0IEd/8V1tBAmg8zS
TEmKQbEz7DBwa06mGfZ/s+mVIxTfcWhM6Ggnxo5GiYNHmDcqeBmYLWDVM/U+7m9GYZJjpYZ1jyRy
rBK0D8jC2ytwCGBHU/dgR9MTpUuDxZudw24HuZnSQNQiVW/wWN0FpX4RPCAxuO97gB6D4m63eHlr
CTVMeb8wWzMsReF0O9m+JWT13nVsNjsPCnuJVb2Ojdkv5plRyvAZLxcXczax2xF5Kh/Eanjr7bSF
COt2wz70XDfVDRf7M1s3vPdmA24hKbZUkMH/D6vAXnXZhpAVrGHoDxbpR/WV6MYgWjT6z0z8PeOh
tMhR7m3o7g82bzzHYjqvYUxiuCJOfs8xjvKzbs3sQghr3pnk+mhCQUrbDoUhMIRy5qRbdi49Rnbx
yhIQYs8qAINT7MGmbiQxGPxPp23gSwCcm+fk4ReKEtaNv6claWYyt/rr2D3gYiV3mVqI+LSPm93q
m/yNP85ndmKy405Tbr6aYQHYLUYn5c+W52gnL2XUMj8kH9F69yY7XCtlv6Csd3BBPq3Uy+1ut+Wc
apdmkNP6VkHkWVBE8kVejWiWtweItwNVpcu+jIqeFF2smirBbA4VSmDckSlQ17mcuhDgFunKkvFN
6NKHRpbKWPglRfJGc4ft1v979QykG2q4cQRZxeBcvzDYR4QM4LsxE08ZRMTp6EmHhVYFKoHUQtWW
cmur57hYu4WquBy468dIBxAwvw/Ookdtc4V/E94OKb7tJmiYRLGgsBIXNJ2r1DhAEogjEeAQLM2R
tCOVJfnJ1i9rIiiVUVRpfUnAvs8opKDGo38YavMMA702FmITfilH4vByLJ4Zox6ob2bMQJynVGI2
/GGRejRNU0XNPY+bXCfn7ij2K4NjjYEjAe42BPkYoWyiKOwWoUi9cAbxjr8idJVjZ95agRS+76pI
+ZyiEfcUjV3h3yRkDrn1veTt8AzyUIyl3Gqb7QK8XHao8CS90HH6hL0T98g7fKmlH/InNUybiJpw
BEpWjoEPBQ4WoYQiPFDqDbnERrdaiwiu01ojRMeY3UaEsEodQZAGk9ppHFoAJnGQbyIX3/wsFnU5
PpO/M1omFbdB/DWR+SjV1R93QAkZGgvlco95o26gSteWQ4BzSOqr0RxSCxSrEIfH55Jw2o3OPw7O
uIDu4mbOTUviIutktHlBAHjk3FKafaQjkQ+3/r3oQAvkLsY4EDxigOFlbr/5gvBOc7EqFCVhkltI
ZMlFi2v5ikhDoUFRXZfMHdm/3fFg6xFZFyKOSTo/yFJ6y/1KP8/MLjPzajejHSyqMIbNZdJpSh2O
uZBGxi3dXNDVvjJ/hyC/DWOgsovokCZPhM+V4mEG1x6XpiqnfsldlMkFX75VAwW7+Em40U1eku1c
UREDwXzWo7JHE5dQDXVEJNHNVNMD9dgrsZypRDwCLhqcKFzCsyt0pFh4Di5uqALeimOEKITogdQA
C3G34UsPUKsDPIkxGQHoasN+3W3GRad9xcr738E3wy+FTf8rb0XVM1iLK2YsB4estsWsmykk9cNn
oILQG3Z1+3xhrdc9OZF85s65uykbsLzf6epeadBAQqhqT5DJ4JPd/LbXEvHNUlbi9+w+xJhlB5R7
fxDXXL6wD/jaSAI1YavGMPVEjCD13GDp9TPT8y8RI12icLvkuGSeNAVNj+3ehDkEARQ4rp03evJj
9FBBPx/W2WwE8NZiv6jxaG7xUO6dvFzFrV3jlm1H2ZxCSB43h2C9rDwNUzatSsRatdiYSrLpy3Xb
UK5ybaXaBsQploGFA3i2i09i4BxZZcvm70ATizIHsAWzFTn1h3Jd6CuTX02GWHcpMMlRqapRKU8j
60nXEcHIP4Tt73w/pDxCSEpsKwRRq0MQwueo+1dstQg03J1RAMk3BTZeBO96QE2ZFWRkKXMif+CR
JYIDbDKFr3t5zrRVsqI1ZsgEwhO0YszjmsjPyL69QOClFySMuhl0XoqYt7IuwsJ5iFhW9Tl6kv6e
3f94l3/G1icTjX/AviqV53WcTy9Ve7zCIoF39i+P626vmHEehZ0hGrD6RFSdZFDhcJd3Mu5onRwJ
AL+P/UoijCquDz1w3n0YvtG7wX2uRjuRI4bYrrBja/ZzORXXEFObILPT4rrXd1usE1Ekpd234mfE
Cc4leTzfltcxZyy62IPrFXi1ebo0CCC9kuCrlkEMivgborHSC6gTGo+mFRybIMJ6dWgSy82JBmvy
pJ7SNBbrX4cM7Cr0NMxMFVbO1D4hAUwgKwkmZmdQhP/lJX9oc8Y+ctsEiT3hROeOItT8a0oPg8Jw
mmBIMtWddqNWXusIA5FCTZ0tldBgw17vovcel5F6wY8PrtC+AD/rAF5KKAQgrET6eL88n3WneLzf
BOBAcjEKGK79RwBzBvZubKIt/ft8pvApjY2SnG87yvd9mkvbJslyqE81eE3s6xzSorzFflxUtSL7
5bK9ctPUJoKBJ8SFmSrjNRwSKrDkxDkrYoBaNs3b+BLP/0j6MgRblIWo3aYcIdJu3pZJpi0s0OBC
a96rQgzlFiXt31SlCzMEDgWsJMrWO4P6/hnZr1XGxkMgvxGdToDkMhGiehaWFM6sOaHEGYYCiSw8
nwl01zlDGeTyaEvILVARww+dNqPcAqJBj/yaiUHy9Oey1PNrXGlp0SzSIxw/c7AiBtxQca3cLhQK
3pT2DfN0sVvI23BO2hd00ycYyOxBscqZK+Vv+pNR81nj26Xpf5aqYSkBJEqDjszngz24plP8aFsC
9EgW3Y2uSiA4T8X66chzhrLwYelAJxvpyQBLNGTby1msJBKZLW+Qq4jUivyvsBRgOz50iMMQ1ssx
Gu8/opJIxkyKXkvCjHWoFQof5fbVzXEazqZkH/YUm8uNMVP3NYiRB+fE+TjVaQOnuOpTNxmDuTOg
KJCMeFUFgawZ10U48uAysQbA1uqhPLiiJYfPk5VJa7wgdc0dq/p6SLXKb5pze57J/inldqErmHi3
jwHa8ZDSL0cus8eGvc164On3EPs5c2c9RwDChHKwUAlfHqhOdUvY2bmROaHd5Ye9vGCuXwHaKvJ8
WnnYfXVzbto/Fapx1jNz7VtClKDX4xOo3yUXr8ZjGxogEBMn+Dr3XXNjCVEoRET0VUReyLatf7Ig
N9oVFCAtAyMIyeebX8vePps8WN2dNFlUUOQAa2GPdf65+nD2q56oTtzDpnqea7m+/bCFjOnYjyWI
OJi3s/aWNjYYx8YwNxuL6i9UMRqBkyLYs9iLlp+fnUgHsMiOxvsznTiM9fMj1qB6EmN9kuZEjxsh
3ZxhJsmtSEx957uzYjvTJRL4LHbjWNAGBMfcvdlZn2jP1R5285kFRba8cyxjeu2ahFMZ52He1ZS1
Bhf8riyIO+qUXiHZzcsFpRbHTqyGgjP17VsLlS4lWiSY4Ebmv73s3Q1ofXsnrr3UkRVdHQDn0fEE
cgFdtIJBn5iHecAkGoi53IMj/2PXxQtCUnfd4Bsy5MMtkIr0M9ylWyqpqfvfoZCUdaLrntJIQDLI
0e5fiFn2zncS5kct49/EXCH7K88JMKH/JYgOsY8NRpDjpbiC+wLERBUqRJgmlG8gav4QxILqMjF2
GUMjshEveLrx91Q4WWLIu+takLTWxVfX0R9d9KJZjSt0cAcAqyEVBgeXNDdnMriIfd60wObGnjk4
F2XtwkU5TS6afCB/wK2iYUcVdq3v16jgBuS4PyBDP51I/clvD/Z2I7uNBagt3IdkNAYum+kxiaw8
EMSz0k5PF3qBxp/x+kgE/BhYlF+1af25FIjVe1Kvw8FEdDFX7gEj9JuGO1RKaD0FlTNGv/I8BAJn
Ctu/zvwEow3x/odqv6t12NNnOlhctQfvaRvnBJ71os+jK9DBXXU7QhZqx5tBPh694TsQPh8k0w+q
HhcHq+3gtU7wcSUg8gNQOe3KddLLeygu2+dvuzP/DSKjxOTxR07CetqYONUg4CQjjpJOBd7xiFDD
yeZ1atvXsaJDTC0RmRGEjf22r07VNpveCyOezrFLOpmsbSMy5QrdWlC+5bq+9sOi8TZSSinFBHXE
ed5vZZodPK+v+S1BNS4BHEBnaBJSUiDqjYrAmf/XlNHN79QFOOVy4ZOZfqr6WHu32pN/WxKwpVq8
aXoxvy1O+Y5NSdSlwztjD5VB+89uCXZL4X4ZsgdG2PFhZ/9FHIQoXzyzQBcKH/acMjlHYunptigb
nHWVS+gLeVuJ7/EfWjOtLGcQA4qzWnUAlDOXLfcNDlvs0Falr1zRLOW16vBGwLEk/35CAZ9bA8XK
3Rkk05n8RfxMUq2GU45cMN4pyC0kR5GDfWutQxnY/xPZyNphaRAroLcQ0UrSxrnPmeaTAqSn4Ohb
bXHjtY9+ClDKIw3Gj99NIzGqC6dHjz7wT856sQuaK7s6mdKyNJfb9ZConypalDlh4hciYKtRQaU7
tHs2HJE5vbobgv10kv7Sk63NWPOCGNx9D2IOccFtAk9xsWpjbI00XUNTndqTRVwhZPEviXVHoVb6
iexxWF6yUlMoFNvMueYYpog5WPY7OpT9ay7aJa+DDeQo/DgiTlhIy/0oiHEkhMc7SP3pj97w6RYs
4+Pw0ayoPkWLmv66LnkFGxIBDsodcGrVcslDrsxmB1rzrdXZ2cy7duoalHRAm+lRslb0+losbIWq
Rq/MYamn7Qn3/b8sZL7u/pxLCh1kJ2Sfax2WLsYE1m+YIb960EWPQPDb9lNQRVumTdaN9vrWLacd
Wg18JR3vdBUQkd59XjcNRu68UUgEHTQ76H7TRiE48NwT8Fz8JnR/SAlxy6+Xfk39Pj2qKxW1ZNOF
dDZb8WWa/t0+UH5+Zofc3433q7fL0lOFnAMAQQ7uk6M5AgtQYOavZlrWU7QDLyPfpjHoKDjl+X+n
JYFJk/D+vRnUxL4wNLRAn8o7lhjEXXbgtVTkdPca9zJ/yL6aRMDDBe2b5Jf8qXPGmNcQgBCeC6Tl
Nje4qvRD/lhdIP/OPYVuZmJ+z9zoFUobqkps0nJtBF7XccmMrEMpfDX4Hx/TxnKWTM9dJ10y7Kyg
DptFyhQT1Xy6feO+ddr2bgjpeZQlB5n0+XrR4xCszWlIPbCQh7F+FbzTyKcW2xhbV3+UsvEKJjX8
7b6NHhcoWdai5i9VlQUuUFhRfX6a1deFWAUgBxarTKSrqG2mGGcXMGDNLfIW8ftsp+OqqM4W6I61
VqtHNpy6qsXgrBXaNdZHsvHXtBOonicSnKjroDFW+bpRo4mCwXPksJN1uJ781aVHXZkkgunQ5TNC
OnoGoLOVcfoIof9ymmMHokCkODsxlUf7fvVCAIRu0LOv1oHrvNezS8qtJJZ8335/SRjCb8IKRunY
modrNMoKUpODTLQ7zBVmoL7L/2Bdom8O1VpJaplIy+5kmjtJykIdMsxSyJZ1n5lP243qbGX+Jpri
fmXzOkt9/M1GpJlm3rpU940q0HadLmUBv/TLWuewriCq3D+W3i0oZOx2CtX3/5N6+PkpSPfeB1/e
o784uZGwlGB+YdbiJAAW27Vwa+ZgbAfMPHHR/90BumsczPEow2J37h4mcCh9omMVVYKb4kUurTF7
gf3Pe1lzu+vI/BWGL9bEY1KKzBnl2Z+FlFVv7qZIl84xkTM3dSSYuh2uAzVhwOoFk3EAozG8F49X
NsrabMa1U0mMSzKbk44NT8QDrziv1rhhq7sRVknHztKmWkRLTlT9RVw1eFcQzVyIhF7A+rhU6k2j
NRGg/3dZcZc0MUdItOq1ycsJP6whNt8birvCBGSRKLymH4EyT/kWyXjCSgGuYlXBeWVZ/72nIU94
PfK4H3EBIFu4MrPbyByJUQ+LF5erBNG8Hw43854fzKzYk20lIKXyDf7BaEjLILjVU4d1yrqeaURm
p3A2e+Q9pNaLR0oSgDyP1gSSTpVYkWXiKXkZfkWr40hbyt/e6osbxNxou1B7LQ0PNWPhAkdPVcff
vZaT13XGKjdcUgTqWp55i87L409v7lLw+gADaiT9RRyu+XGlPNbQQN0hKPycVbrjxvR28wUqmLZ5
jRnmL6jJBuFU85PEDrZE6ANXw6ZChHabhprHbFK4YxU4mIU8fxqwcpiJrvjvmyriOt8alefdHE/9
v7QiDe81jpleuFCwyuXTHedLZRwCmHzzkeUWBeRbVm78BzSWawAJSuylznTUeQMKFAkgAMyLBhFQ
yP+MiVhi+b04a3rBCedJyTg5cbM6tWiOcZB8Mp1TJ6eKiCLiBvAX8Sahl0+Qvo1TQmGBJqMgGDMC
cLXUeI32U0fL/ON4AwAlLYPCwgEv+bQiMgOlcJs8+MOBJYkdIh7pBi9ZCLgFhtGUIJDyfAr0PzlW
pJIi3wSpxY9E22IsSoe4Pueq+mFNObaPuRlEUSFRD001f4AZicltW1yHIfc0TA6oiBKbjALtoP0v
+H5S+YLrifz43yH4/q3jb3u/jaVSl8piCGnwtkkA/lftj51btfG/OrWfW5aO2n7mmaswyoe8KIR0
T71sCe6lZt/vu77N0COoEpJXs4pIH/kgi5Do50eBWfO4i5aLFcddlmzBxjyO76yUDVvCAdJwPpEN
zHy94P6F0xnOaM55eNhM31WznG/CbTXfzaMDWTb4PZg6AxvB5/MlDro2FggmoV3bEEfHOlm0AZcf
pwiIDc/FhMZUq8VQyha8F7YN4Z7+qrcnpr5I3zWb90q6cAntlVXgflUxZMAnzmTC0oW4o0GDMqzB
FDk6toKSFUDJsvCC4PouBbHugJEnn0E23kxBP46854KX35y7VVXtrXD7N4omwrSCcxSufZV+W2F6
pl4geX04978B1L37S7lfNKet3Q3ed+9QmqST6b4JvERxiJk6dPOasfvfUVV8sM31nuyGfNBzbPi5
D3PID7yPhUNCnrPPwRaKpV6e6CDmkZEiXqCTojVQcC/7jx1pa8Awvmt3NVVsdfa7eNHd5lj1lL9V
r0GfHsDiiw68aYt54uWpK/mUFpHiAtd3eLkjSpycKxmaVYLkLN3ba8HVVu0qpeWd4DxS7w/+46pf
URZaOsDDXI4ZNCoq4U6Kf9zA+wDpHZOzQwbx5kEk+AubcSDr0Ii7OcZHWh8dRztNZhoPwxByl77z
CT7CeYjzPfCBMO4RLQvjC9fxNaoQn/KnrpxeQ+BJvfImcAr6cVYlkSWgsu8Q/aSfXTGcNQGsZ1bD
UIn22+nsXk9j8ZGm12Z5G3YYCVpTovppWCZ848K1jRHaUtyYnqL5efwHwqTt3RP7jFdTKLW0vnVm
Jq4WmpPWc9jVPqjIPi4PZyce7kFoJKO+SrckG5w6VumbiLd+XE+TJpRcDS7p+SSbNbGTaIfjvmQo
DXRt8/4+JH22kHmvT69e4buhe0986K7dlGiVOpIb+9pqXqlOzhVbJCwUhiQVu208opLy5+EGh3nc
sx77LY3bbK7zuX4eo6X4S3+yijRAjIxH1EuFIBOwP4xhppCF2ZJvwkJ4Oi9/+HxsvjsaczgP936/
cBuQ7qB9SBzAGHGga77lFIHX0BGXpulfI4kL3SmDw0EWB+D4jSGiXukEDspzsnYHPY6vrz7jTb2s
SFBq9306t5JFuB6i7aNpfhLPJjBtFNk8K6/5hdfBkDwMMXy/js6WUtP06Nk8zmrT+bKXwbK9R1V4
umbNnWqQd4GMNUc08R+WOYLwYgoimGnjj08yP3kijFvX7/mUBgEgIToNwjFQsgCWzs0NDw+Tm20G
cn9RG9ZxSRiNYmYhn638hLgsP+uh25oPpgNE+E/76jMOmtYQBC4pdb3N12/9vzzfKoED5Cs8SLs9
OSq154Cb0MZP9pxA4VuCzd66a3oiZwTebJZzgHx3pCV4NohrG+avJPtqzUjTeci48cuRUBjeR3xT
wbCrUgG4rjtgPvJwBGBPrGYisfXczivMwi/3PU9oYVPShjxclyq0OiOFuicmv/LvfgIM2dLeD4d3
2pij+N8fUto7rq6SWZ2H/poM5DIuchBxwqE3aV/2bwE1fx4ndiXxy2SlWsnNIQPKw8TeRJnNxJ8V
D4mbLNYE1CH+Jm24fUnzrM3+7sOV+pND2E4O9AQg7p/UDz5nTudaXovyGNYasUJsz9+TrrNP1Fdx
paH5Vh4hoJotVqYYUNPHRLS2JEyMHvgx2RwKjcIGWdWIq0otSwQQ5rbOVR1twkBhxceSzzybKgUr
p9YWhWXjGrc/umqIEMkIyTuTdiYWt/F0WnTlI5Dcfd0WwE8DTksQMrdI/j4PAUn1TVfgVz0KdQA8
TMR22XQZ5q64nQORriqjNh2vA+y2db2wD3E5klN4o4Qk6HrP6l6nq7e7twraCVEYr6v4VWOOJwwI
tF15D9Se8Hk1cTwmodLOgZb89S2juD5keDXnzG2V6/T5Og7oXsZioxwwA9u7Ex982IB1Qe41ijyN
GlzYv/V+qBfdo6rUlnLBPFDGrTq4lQwsXPJEstjD83gfZG97toLqs3X5xuH4093KKJu97DVGm3TM
vX5S5uKeb0h0Zp934dElllYVUs5CvF7ZXzWktb4ZSY+RMNSHXPOkUuoSbPgj508J6Sc5d0JSGxmx
UEGP791Esyt+L/RqpOnwWmg31fEn2zWJ7NNtZHjYQCqXoqx8JNrsN1XknRfFOCeC5IoIhP4tbuBy
RFbULvHaJWZzFvLVJFFRuyzjhCWhByVakFz9uOI8A1LyMTQvNPtaRg3nmxljanyAcXoiKDFssVBT
xwfsw8Z3ZPYo0YkV4WplAYwhE0rgaAbizoDVqWFFF3lT8rfV0iMAUBK65Ry7+DMQMCqA9hUssvjA
AlPwaFEnJ6ot3KWKyYvyiWi+dkfJqIumAnPdF6UUAUtISEdX6OSHdfmSU+32k4DV3BDn5HP6AIhy
jxLFis9KOBqlBJVRiowHxaeoaZ6ugzsRtevisu4uFsU43ayo8IGqFI4QsZ+IIZoikGvm1B/qgLW9
kC3eA07Mw2JJIlZayJduy7JMPMfPecZSFUqbYaYJ2IOMGhUD/OnwxcbPeaewtO8i9uLqWZsC4Z+Z
aOW37wbEMAGZFKMN8kKXrqTg+lFMd3yCMqKENXZ1agXsO93PZcAdP1M6MOwgmmhpexGBn6wSOwir
4HBFaGO/17+XJmtdTbC0xqeBPTnaep633ZpDDyNc0EkWJSIrm/uZk61jOWjeRGAp2lMCuCG+gH/c
s1qxWvdv7BCa9xyk522f5nPYjWb6QuRtJlWrG9vJKB/lfbz1n9N2gU24XrieIa3KeEYaOcimJQky
unmkSX7wimk15QJysLEukRYV5PwQbh/kxLqCBvom/CT56OEcluiGyv7A7blT/kttq/apRsnjrkZX
rWoBRtyuIrGo6t+X7X3oY9sGoxPaGZj4k59fdIwgCgxUI9mhp++brNNswG1uaPjXsplN0yDoDQhu
tUkV4+1iQeBQhPwG4e59iRF4ViOoXh3kOw6fs0dSktM2Vr+M9uMh4ZTSV7/mN1Au1drCU/5jpOXK
dxDGLNFI0YjHRqIXTsT0nbmAsn9xzvPVfs64SGsmKW/SCqefO9q9NyQMawm94fvjtueYNr7NCFHl
d37QzfA7HcIpK/SBI9BtwQuKTxgjbCbT0/bt0uBhRK9AMUb/OxR2ovM1UOPaYWrdqVPzzW+LD0BT
sTxaqK/UfkN2O/DgGXitnHqwVArXjIEWpMsjTbFFyEonzqmrrDdXBnxGVc83GL2vJSEM40GvqcxK
hN5NO2aFbu7Tiv5DwEbQQxpMBcGI56/UrAQQh6I2RMWeEBoofWMP4+51ojuo+vmDQZHTvXM0rQCG
igNrDIRJD7+oJtqP3JZjZ/yIDVY2EFPlZ8S2MJXwl3jKW4uyKG0pgy11J9JiOWKX6XikNpEO302A
f90DyhEW5EcLlP8D6L5CRMyvDj6HGDFEQxsr5QCJXpSMCZOYUn338KPVENhaLux3mzybxeEtpvCZ
s/7LQKogXd8jaZIz7+Pg77L9K9sDUw5QAu79/zIR5IQV1V31Gh26RMcfZ0xbXDRSwi/80EbBK1jW
rX5QzqYHR0zlqL24RCMaH6E/fXllmgo4lB1235tOyNg/akQdRyTYb7P0AslJGYb2YX1imFNKEzLp
Ek9ehcZskpBduXyXOb7IJ62osZGZDZimoDRj54+Xbc9SupEOFq/LZriEsKZ9aU4PQIglkOYhg+08
jiXXyiicCzFzZgAfxFmJVW5LirsdPFIBzMZyrwL7N3oqM4OC0bASchbO6vmflIUIR6zOeOztC7Tq
RHafvPuplT5TUQPmfgxWbm8q1sNf7JGtiXDrytyU+wBth/YdFEFHL79ie7NhXUySWcYiyU9/Vo58
97zAINZtU0lCyZGvVar0a2uiAkmuZda/jfpWTGEHopdEC1LrH1AI5Ydo46RWH+Zz16OZVTdx6QT/
r/GsnacD+89dyUAW/AnmXaQBmnrR4dP8GPfjB9+7ZMyCMeP/9ANQLLi412P3gogQ10OUYbxZLsiJ
HgjNNQryXNNKOoS2ePzWYuvmtxgp1bt/AjS57Ksufqm1kHmI78T1XeVLhKRBauFQjxrThMDnVeeX
k80rXNSzQBAiEoiyE20elyTB/uxj0p4OMHj38YVsRautM+Eld+MmWA3Jg1l7laIJFsdauL+/4uej
vjC7cOyc57VfFChf9wSz9oXPY6YleUwdLwsezouD5WDLeJ8LatQTy6kT0FxPYinjcd4t1MeVdhmg
mKgZWPSywIpwsumrjtY/lp4um83jZA54zJlE5j1Su1LIP1LJmRza/Ba2kLqx+IAjX6qtIcAYxw1Z
FcTmjIEoQ4tSNXgVdAuPX1QqJB4cHGwf8TqwjzYWqZB0zNNqrV2P+Ku03viyaGdEJxbemwQ+2lbf
9atGbCA7I4kVz22gkPqee3G4+7wX6jL7AMHOvXT4hi8rkbGPMjd6c9PWLK9rNdsvF5NsSBfp73Sk
n+zPF6O5cub5+ev+mqGuGQ+tt1h81yrmiIq3maR8AhdGO3SEK+oyVfqkWNgOhc9GOuTbU6DDBEk6
wxJDxVZOqO2rbWc+1JVGy8Q9NDhRhLX0Gpjm4GtKtIE14zxGaF4cW8e4pLohtqP6NevXFyoPU9ex
2OKKdfVMBUG0U6i5RFup1PHd+g6VuhOePWAt84yfacO1NcH/NpM+LPw+VUrQGdewHdJqud7oLseP
y5KgCam4MAI65dTYG8r9kfte7KqhImVtDY8XgytMZIf1Huu49y9LvqS3M3O6is/dhLbF7nF6J8yU
IC+kDWX7kE+PUyjTTGyR+ZwLRx4/MDNRKAuU/4ZqtuWwQuopNitIdSQIyzna4iiLsNnVkkH3J8A/
PGtIyhjYeB7ps221SK2+ZzxcATu80ovUbrACLn5bJCZddP6HxVkhCoOeQt0bvES56GFzHJ8FM9LV
pZSnc8XEAdtzb0MyFk4shXzMbTGDyuoXfj3KrcIPcUbiR7GhSSpPTT09Imiu5l/BMyMCBvgPwLi1
giWV5RSMQFEkkBtFxOeneFSnV9760DVV1V2d45+AyJCyzFf1HnkKghuZzTgkg3fRwYzoaX5R3JkC
h0ASCMCgWAIVni2hfMf2ikyMmbYOm/ra85J8R7JPy8PCv9rH9xfoOYpK9I6ERwUzts58cDe3JXtK
qTcD7aWi92c/KYcabzsBgZf3wRi2VdxcQk41F4mrVjYbV+TpeglyPUD9FR6iudyezHf0x8zo+fX8
XsQuWnvcMeRw3GS21eMZ+RNEQ9aTBY3uzfJokrnrMtYdpzHOHcve9oUSAsepBIC+UYQdWUH0CPmP
ML7lyJD4fNWbGpvPBV7SNeypiuHwpUQiwYSe6Re2pHw9NDfbzEeS5fFfc5hu+cvq/Snd3abFJSsw
FQqbUUN1FbGa2YoL8w7iB4JQpBVSdJL8RGJxJIV2qcM6AJ45WwjR5VwRMU7V0phchLXd0K0O0jGT
nA8M81FSuxT5rLd3vbNHAR26G5GuIiZmY1eod7iIwegMPYjYAcLkubU/vsP5mrMrslI+e2MAtpGw
5eXmboDq5ffj85kIcQVvtZ9zNYeJ9vaGBoygXStkw7PgVgYg31DJ28F/0lzQ3b2uRlXIzDwg22Cx
b7MEZDDvRqAWFc7TQ1Uu+vVaLeUin3UcJNFJdTQ8J1Xy1xCu71A4Mu64o62MJjPgf9kbduWOt82H
3vgLtPk75TBmSDbnKKU/GdmytWfxA8hIq1uU/PTV6OU4yvseH/jnVGdYEuE/hfSr/dbq2Wy37+Ak
yK2wDIscD7uCBD8CUsLEIR0kgBjCNUEJRaGkbCWhzsBwSlb/dY5sWMz3CEvlyH8wJ82CT9v5bhmL
0+mFvjDEIzVlWsXSwt0Qch99AOo9tPa8dH+jvwuHv3feczXi0Zp71u2omH/NOd0CUy0gJAxk9eff
4WqVBmhoVDeywdhT4YmvN6f5JWVR7H2zonWSmr1rxM2x8dDd5oqCMeDURiJb8wB6PIo2oAJx9SIs
dn7rL5vnd0qynzLZVLhyn1J9221EJvHRdasuwwwajo634ffnt646JHn2x7vmqX4/gyj3uoKmYq7T
XMhUJUyFtHl9ydp+nx2ITOJCtK2Zcx7ZVKiwxfAtomZs2IEJRYjcMdA2f/RO1DT+eWddOaCB6d5p
9uAyJEHely8LIniTqUVVWszSMeGkrOz4ZgPjQrbG9vviH42xfINb16z0E2xJ8T9yIbM7iEpV4okL
yiys210vx39GDAu4UtYWEp/h7Rydwyk7R/3GYhWs39uuMFuC9yI+rCBw5okPelWXiHM3/EZWaE/1
1HG2OpCTrHJh/QBRIlJMHItcV4Lo/CzpeDHG4KnVthdWyayKb67pZ1lIqASHBffqdRw9LfsxOPXn
iICW21iK/SkDnmBgQCmvyda6rEekFkLidT2i34kH8MVGS1P9QIYY1M0wS1ig54z752VTuEr4Bxcb
LmseG5Be/Dv/EtDOKngVxmLfHqflGzKwazBEroIqgPFefdTHDg5EuPznCPzn9BTqnb+7i6WLJD2t
c2J2MHgfzPxglwx9B00EcrcsmW2Zm27LTJhfkVwqK0eUqqfGifKWuKX6vC0fsSD1V/vuurifEA86
p7vIYR7TqQruufeHQjsoCxd9FdkE95fkx6IRzuDD18ULkHQugEPLWl0Rkw+oVHsePx57LWFQOrbP
oTBCt4T3QMUUx/QPP9AE8q0gWmYzJgDzaLeRXfdh0rFrAWi/K+60cXhGTc6JbHJ4saTncQ4PbU23
J3AM6kZZ3d2DYeouYHUgTwyGr4gYi3cQhhiCp6r8oHB5ZgvXExWRqOGR2gGH4YV6EiY+I8314X99
hXpPaWNzQNoGnUBVGeIsCX6VFujG28etGTDhvZwfLW4t6FgRIlUomyMqJBGzri1eYFH4tRMIqBX3
pDSINvfJRRerJW5pgn3wNY2uilosggothsq/oTl0CH9ZaHdJCRvHbq9EUqNfK0nwhFDtWV3fAIHV
r5AVRuCrEJlLE7TrKK2XaEwLxQ5Qd+T9yvGPWkGjVfRaPsg55BhH0iez9+lL6oQlW3kq5+6+ha5o
RWqDWs6+m7EMbAOtenJ6GgTXktJiRNt8RTwrocP1RsqxeoSOGc4pjB2KXen0btG85ZGI0rEL0d5t
f/7JLCVPmBT3p6C2GRPDGzRDklW664CcvWzmgXP8alAT5/yCRHshjRXCRxelhiAVgYzqq/CY5rHa
AsdiqJSVI1EGwr79NxX44NstalS0bb8LsCoYBxDRh8v5QbbgUKSqXXrR2Fx/ltTwR6+kBBopGmZC
gjKplt/xEKdhtOBYrm1yWh03rM3y9uAO/CvRnP+cSc9Uh3wbK2JbLnygzkwwZU04e+zd/lMO4Cuq
FUx67ye2t5800VVpBtHU6DYx3mXrb5N0aXGEt8jtQdW1/9ylbvGKewfUNttTRqZz09eR/ZM7TS50
ESOLKXg+msNF51GY4wCZnUW783WFNktnv38clpfEZPeMp2EIuNu1RuhaAvCfJy/z4zKPDt8QENWl
Zkddk/4Ll7bm7ExPuviRRWrcssiqh5CQaAywotQDk1qhJjzKxUfaXZd8IiKpgVuTDtU/QoNlgkDQ
wOCDhRNulMZ4sAJF92GIqe7Kt6tC+yMkoCUbwv4JHZJ4nUKPXaFrmQYb89ApJS1OoVz3sTh9XEKW
JNIkPEz1qzeLBlSacs4zYtgML4ABUB3dIlz130dWGxFGaAllqcDpf8ub3L0Lj4LoL0u9TqRP214n
IvmFGdsClhZ8QlOF55q8E+PvZ7NaeWcHBLaGVqBt8KgRrHAg4Wh7eBq63V0PvCw2idasFs/eHmQO
+tFc/ia+psGjhMr1NL9/dRwK0dp2anuHW7D+gX+w1K6mJYGpVamvw7iF2nBE0kZ7N4a+7xu+/Wav
jENN9xBMMZzhdfP2ab7wUmA7aLAvgVdBZ8LD8sW/dPQv/Y7SxO0ygGZd/A1MYIG9nqa9ICGH6YVz
me13caG5yGLS4aOeFZsLK5jsJ8v4GUfrZ3kiI9ArbgdmJLN7eA36vt6gcyA02ykY61pHcePFz0t6
RHh4HHVUbhuDEjfEKHnU1IdF6rumS80xmgQktxayVotbm6eHceyHP0KXTLSPKkJYCmOsjYoep45R
QQrZUHXKMwKCp1lPffJ7Ue0O4bM6JhZGbFwNx31W886b4KpqBlor6gV0nPgjvie87NpBtWjIih47
49+rSYykNipEX6evtILL8sFwQjykDa5H+64VM8ZemxN8R/LfNNd/mTH1U85D2Fs4Q8KCG5qP33ls
BdB3hg6gwlb9B61SDzygJGD264iYCXCjHiJqliGIHc7VYO9vTAIPBdfrm1CXwnGcfRm+EXj288ik
Z4L3pak9g1VwGpOOnZRd28p0TWdp5DqHKBZKj+1/wcWl1gfhCe8KkmoLKqJwjSWtH3qdsyvXkBHV
HlYKYSi+hTu/fgioclNnZtOBUdUzf0IhmGJgPvq+GvxppygIcsjXWiFafto63kVME92z78sZf7CD
SOXy31RRsTlZnO+ECIBqv3YS7jGjd92AJkW+v3NZq5vXN1IBP5jhqRWd0M2zSE4GISrqn9+NEI+R
0KJ376MFQUghfDk8XgqXfFvDdl9gHDjfchwAzIcNOAbT2DgFJ1hHxiUrU0lR+yC158U2wMO8ywPF
nUXeyt2kZlQnesCMgM8t3fI1ONT/Gt8J3k/QFDL3PaqWeMluWxx2HOnui5P/MTaSmMzBiAdDdZrb
CNNVFAPHoAimjfONkgC8MfuQyV+WmAqhraM+tgVH9H2kbnl7UW7cTNC21x7fyG+PEypDQZRCkNnb
AGl9vgm+lUgpm/I6m3cs/q6gcqsEd9W/Ba8A2xcU3HH1H7uTejM2q7qEoxHzbdhGGRiVYpKcIOJd
MPQtm1/3nyl4CIewdaRa423NkDJDD9tuUDhprUzOf2JBh+ZTodT3qMgouPx/9sdBNC4qpuhoCxAN
RSJ20uyhp3YbalSDA8agO7pBVjwuQkqYBcTTHpNQps2ZD270R+D6gV8nIETKnXFoJevbpe6rEUwM
JJAs0g8l0PeVODRn/x6l9d1ZZivW9uQ5SHExD/kwCAI1kusNpktdXcrkN5NdpNQiaLHam8cWXZEz
Lk/ilJNQYQoIBzTjlZEmcukyiCdUoayk5BxGYJsxoA1JdFihVtCQylgGgJghwXWfZGA0V5G4XWzU
WuGKLty6Yn+BbQPuD6Q5Q/elIB9LUIXacz9sNMrEksI1saDjmYYHxi42uPEByh9ICalj8J1QqSS9
p2sLiPU58cspetdzR0resNMymdqgm5q2+KSbb52hKEYVcI3YAjLk3FUDJOvE8G6m3yn6TrdwOYR7
/MyraRbX3R9MTOP6rwxVEXi9DQFkWKNzeCLvQmJsvdi8AIeAHXPHrQxDvfqEuMPW7Oh2m+5FNxyD
/aiPgK/4ncieMO+x35hEcqZqglFT4dS9eT2B6HN1Dw9KARhhffhMyEusYaZn/zwruwfWmQVRX0Nf
IytBB0cEWF1UUwyMbYuMcsKvyf+Ri9O7mIUClJnOxZFEXfvHwkZ64fjy2KZwlG2wpVkBpkFugR8+
kB+WRwmuPeKcPJABQdynWLYsvualDDzk/AykdLesHxe5Q7XpECtv7JScYnLYM7oHGjTgnhCiUge8
RYwAzrn4yQCF5yx9gT03ir57lS7h+J3qt+aSllTEhp48UoTafQ1yyJOPUnlMls3dxUnjBSTozG09
l8hgcOZ39+xS/wc2GvFKx+nzJkcCPcxHwn3OQpH3GKFKhQ4CAuZPxNQUSiRUENov0FUh5gphwTfM
SB7r6JCXLnHIbjZ7rh6zy3CEMiVj3H6Wv7QaVAQfQVUacbma+4kD+Yj4p4J9ccwi9pul6CN1Tkz+
mya0KqJzZ46MViQTeqpvQCpd3E0hfg6awSVkFw2s0mFjsRAw0A7asIK8+7mUVns9oRlBqhcHo0sZ
BSyIHxRhDw7IxLE40n5qxiL/9KW1P40Z+Glu2794peo7O0Vvit59Rwd0kaS1CDBD/YabNYcIaZnu
GL95BLaWBdghhZz/cLSJnjLz4n7Y2ZJPgy/+/qXDIavaD+F6MckPJZhrO92Vz74Q04N5HQeDUfRh
hMSsS6sIw4vClGZgDSTdkVGGfh5Hk7eWpqTFj2P0beSi047su3U21/02jyY7q1Bo+PGBX16Lefmh
XTHb7xz9ygUUxvllxJn0tRGf9cqBFXCFkbkGrnAVuU0aeqzYyTBKk1Sg+aNTfTYG/rAR4wWh3cgF
kIQ/HxZneQPzdneNBlpv2MylFHvYY9S9FGu5JVHRxs848kV0Gb1HZv7Ofq8C/miwM3j3CeP9S35N
/TViOA2AR9Dn+5JALGQoKyZQDtpDFSfkOnottm+gIJpgUIltUid0/L8Xd+B9LSucCP4adaRwbOvp
E+SnhlnPXwoZcJSAIw5hmXwR8TrLwltyhMpXPboDLjr9mHkaTJVLtssNt+YDOHJCNgFdTWtNWD5X
UvXiJ17rNHYpSYGfICaCKnhDbJSsq7qhzOeoseueFhkh/h9PorhRQZqZiaxvOuQFalYRQ8Nl2kGN
k5exXrJESeTjhsWoENqHQgCYnZgBE9iOxDNWpLyoVr7WB+y7kBGOS95bAU6PoaMpXfVhOyjDR4pM
6Qv9bK+QUxV6+mDPmqn4H0jD7oV4imrkbZ8A0aj+dINWvmX2JJhNV5TMV3rnGrRorUcRkP7jV4Oe
RBLNV+BdwaC6WV1chqYu92dgOJmn0TSzy+0Jeg22xwdtWKH+XIkjin5w3uiXioNrbgzCWNCAkCRO
KoUJdKK+ETZt9sc0X8QO0U0wyt57N2KDE7Oh/mBjSzwRt4x3/pYDNPIZXHE7uDjZWUDzJWKunnFT
5t7R3hJC8malgBGj183S52NJbK/poacZwZREnxKOXBigEegi+yzr+b14ScaFkojWyVISpnt972Fr
ac6Me1sZH7Tt7mfK32FVwCaLrc3mJ+oyNDAUUfMkkSgSDj8kNbJRbL9G1tGbYg0cVRPoonWJAdFz
g7A8rUrywqAIVMykJW6J45IcCS0HW0PJzRenOvCPbwMowOS9HmgO0PCTOQokat5AZL0DBX1eCvLb
tjjDU0mWHELSEO2NO9r0nIu3wH2slXdWEmZC+rBcSqy7i5OKZNUyYi+oPYBbAEK5hl2azA52nyVP
hv6XAvC7W6Tlpge8tYxG6jlB1+WpFyJaw6svQcf68sa7gzT8eG7pgVbC6D+7Ev6fXdo5vVWiBhDO
JyGCNrF7VlM5PFY/L8RwvngCOdk/nElkN9XoFc3RqQgIf456ycTik2stfGexK30q3GYhD6Wol4Fj
4RsFVDNsU15ZKXXhzwGcF3z6dKMFuuIaOB/hTpzCA+Errlfcg9tDjEzmalXvQxJEpvth3KpSj24c
oZU5f5coGnh+IXgC2fYc5El5RFi5ZTAeGPjIUGZyVVCAAPDw+vyR3Y4Skfian+EAXifrtrYwDVTj
qnwQyUihOjr2RIGQ5Evwchq7y2I9ZFdBr4dxtOMobJZLisra5o13IGNUIo9sL9tNqq3UpVVPOTR1
rQHZnQBVrD+0/8yFrEXiAiFV6ZamMUknR9wseO7tLMHVaBpBPXhoCnAyzkyzeVwtB+dliG1FjUUn
pZhRVlre7vbTDOfQ2bhOaSXQjnuLItCtbrcgwi7J1286bKVxAeYX1zC/QQDf0UdjNj/CNCUtQg9q
VjDi2G+7MEfkKLOWAKq/L8IOUl8ebWOH5tsd8g4+Gsc8x20iw2NpTltkg0gmWftOXY9cPDOjMGhe
CW7NNKawl1W8ppmn/ojvhtVaVDapOCOjYBG3c8YC2LhGU//uSV5iuOUxRXwcdv3QDjrFQ2u4P8v6
rrpXfiLw+HZfLg7qHyxZfZusHpZqnK62Byy7ra92Zd8MHcLz6WU/5Um8S3gkcHkMn5v75sUNSD8m
JuEgUSmEldkVRjlLAcqbol0chCjivzgnYgxqnZXZdPxLqqq5YEHoWvftbbdlHPgEFr167Igi0FYN
8z3rFco4RAXYoZia6tsqBCBckE+DYGcPZ70t65jgEFKTyJK/M4UnKKRGo9UQxwoWsbHYhvf6EdrX
i/Pn808mshtXecVy9YI/AqqEnMGCqzUH3IjMleX4U6s9znI3cpscYszGmaWDLWJUQ3vQ/qXOb1g0
dlwt29gwt//VL0ZbpD6pqki1egdwMcW8y3ZO97vHXI1rqP2+SASNCkITuHQ3Cc4M3VPWtg3Z/Wiz
Cn8ccqLMMFbIO1IO5dVT4N8BxTAkgJyLX3UWowPO3Qbg3EDbIsrN6Acwd5bCQHZvEfVzsh/P6CU2
EG0tbYiET9nOi0hWudV4Jt3FWHie8eInucJLbnAIG5RESG+fdwq0gSlLievs8O2FlapZEV4tppVT
vf2dW5Q3zsh8eP8V3qArMp2UbxY2C1DRSHeiix6hr/zwChzi6bpr7gxBXVPxBmeeqdo6Yfq+f7vO
n63enKPHxsX5rZakACexRvr8s3XFgJ22k3n5fIAN58t7LONASjXoS9zMxz8xMVoZ70BeGl6qsNLD
7b5s+enq0UJuymXG3EVJ76rxDiISbY7WSxdz/lC5EoGsWHGXigOp9nofiesP58YZX8QTpB6n4XtJ
KyZ71drqH/xnCFnbZKEyh7BLZroNV9Xd43o0oiFIfJCk+YZPpwyqNd6RuuZD3hKkBQPu252y97Zd
P1qzVp3GcH0gsqD61kNziI5ULVnd9L8EBDGIJvgTXrEasoXDULEmNy2AYt0M2KIYTnGF5WxD1Df4
0cNG/HaSskEWowbsZkE/Ok/5vjMuY2rnWo8qi6P0yHWZsItXfZHOmftIpkhFKeMq5Fo9Kdbf6SS7
wI/j5m1/n3kgiikfDltQFA+722IsWYli22O0W7PFydVjSJv1h2VsyWjhPL/awuhdzVEeM/bstKSU
ex91bpgU+g2ncOiEWDsEWwJ6nAQrlUMJqv2FYa5KXYI6MGgJ5mr/SmH/TfjAdpeSrN7vJI/YvbJ3
GaiKLRSDooB/Hv/4IIOP11M+pfy+Pii5ijucrDWh6f2iX6pUbWpZMuJeRSbXX8RMP7ugwswk93Gf
4sHorfyfTsxkjX0LzLmlTsVaB4/tlKibobLulPjsMURzAzN1lZ3tnY9oirJuT+ObwYq1tds3pv3C
0xju7PHFURI3goLEghXyyPCNOGWXHH740dlkTexTtgujmgTQ0QEIsXhkALvU+rH7k2a2CkQUodJM
oKlK6fhF75ZVK6LssNG2nd4o6pBLMxZg/hjyOTjnvp6KWsRSXAnuDmGO1VmCepMA1lTfuq95QkSo
CYQqEM+EMbPw674LHGvF9PZLWnhdZ2E1daiV+vqzvg3mF3H47gnduFR0K5l5GgBKJPMVNTRj/p0S
kQo33Y9JeI62Yze9kOblnBG6h6k5Koqau5xdHVMsdIeWmtyX2Rd+OxpszRw3S6YTccukmVdbUEyW
qyzvDTGPvmxnAxhXmT+R7Zpa60THNLkVlgHXxBxdIPIYa6Z5wWEAbEMzYxixHFCCcc5XfgkRBTC0
pX9+rSpShUNPIn5retkee314Xudl36WWUOstZqZWfjkMIkpCxRzF38PyP08A9d3lZrFOfLvBSIrr
+O3v2Wt77+U8LtUGDuI40QLoQAgJEDLNA5Srxp8N85pIrDPzZwYf5tMOgV58wXi4cVABSFZbbaif
YcCW9K+mJalkcCYrPJog/vKvQEtQdOSHNeiptiturnAY13RatZmx13np9+jKh110zT13+dBD8uFG
WprObW4DtudlYm3W9skuINaOujRHIqf5+fti8u/g4sbKIoRRcvASCkZiNitd6r0VtSxvlHp+jC4f
0HM1m1DaDMwHuph5opQe06qUJUc4o9POYw4bmtfh3iDy1Vb15nDz3megEWXExx/3OgSeRPFF4fEP
YN/CEneYjZc+ait/yNzx518RR9q2nZai5hU11smL6IF9NzcikgOVki7F95n/zsFEJ+zXpLwx9Rj2
rgE4zdxe4NDeEsD3C2IMOBw6bK6hmIpBOi7u52kNuNkw/U1hlyRv+F3XinytJ2OjTzgP4wOp7nqi
8fOamv4FOo27tpLomTLw4AMJ7Pg/fMJp2LR8odjNwfDW3zpj+HnGp2Eo+MyII0Z5sYOZPib6AQ6s
I7bNTZp9Sp4EZfFbLI/66cVqPkl68Ko3fNq2HTcHbdDQhzVaNvPK2ynbMPUlAkRuMacGcQq6LQlk
WI2HuGTY2ykpJj0qo08yVMI03OkZRvpTo0EOYxthwGQKa2CfkWGEwJBTUsVUXRuN0X8UpVcGJJyc
1L6E1Jj7GPqqfa2lwOiQPTSNebdE1cdlISGVKyZ25nKkNP02x0zX5FpjUuTCn1M1dUEZt4QjwTAB
4k9ZwkdkhZ2oHCxVlGmPgKIDhbIVMOEYivwk4eb+JPsevpjXD+50ZQ5MxwUCooyb+qI2mhouPrxG
AAEW9aYzaNe6G1ArUs3YU21Q3+bVPTJhl/YUeie0/BayedE99p/yS+Uxso1Z4BWVVxzQ1/lt4v+D
Xs6Y87gVvphf3Usl6r1fol4HJ7yFqtHsKJmfh3pvjDGCZg6+d0uUNroj095jQVL4kA5TAcTN81jU
bcGNMrNfik0wTPXYIX/b3pM/sXxZvWyqJ61qKUs6cF0oqtbD0lG4l/AZIfEoMNl+2Zuw2TSp+Q4C
xuKvJArN+tmX7ZeRC6F8azM7O8VaJrlVL6wPkjGwqWnQkyQFzONT1GvCpmFsnjHK4h1uYOAsCqKR
69hhNDlipHc5RxvcuxVeyPPkCMLOCOv0ogRP0cX+ZLLvCJTJu1gh32tiz2smvdAKB/4TCfQFvlzc
28MCCoCbORCznu3XMrgwlJORiqBzCkoQuNFy9iT3WMciONCfUHiNF4JYYK34JhYxEbA7Wqb9Vzsg
HQiPwadczMD7sfVFp+GGaEjScA9ys5uxlxMBQcRmbQJ544Ap40ADk51UBWcZfqLoQT6W3RBxfRtH
yU6YPvZk69nRWL8YtuCnLl7V38qmFVUVYlWAtekiXkDKW9ksGnN1n3FLWMatSK9HAxRGNAaK3+0h
kLCY1PW/gFxG7X3OXJBKyypo324OFn5WWt9BVz4aczNocpWtGHSEVcM5221kclAujZiEVNAZG/YU
Vs0N+DrzeNLwRVqEc5p5d5wk8MPHD4Wx8KyZ6WfuQAfvMjjVTAXpSDYr6N3LP9QM6WwbeWFK4Z/q
R2/bXzzMjjbcULpEo0ITXI0Y0GMFpRm4uWWaakzusiRyDK4+pkEUMsLL3THbZ4qccODRCdViRyox
h8f82KQjdEIY+LKUlirQXQuZ/BYte6AXozZV8UKct9ApEztHCRKR8jlW8Kw8dgJq5vVMbL05vifT
r6HIOVxI01adczELDmGfr7Qf5hamxMmi/c0Te5UWwAt5fCqMqsxUsrsn3ig7bXmnoeguf37OtCw1
GTv83sf9Xv9xEFOqmMzbY2C02xIMrc45aD06APG3Lj5xPF8cM2wHeM/r7dv1BWPiMWjwFX92Jme6
BzDz/irLxm5VzJ6kz5o38dFyRsn+21wfQ1BdI8+12uNQ+cyRwU2Vu+qw0/+x7bgdLKzHcyrLjAOk
/GWA6x+j8ANdnKUW4JsdT1xFQ2i/uJ6u1xlv12cexfwmfUiLkq+Ua7jmrXjIaMmY5tRXassSEeJA
WjJhIuZLo4z22GxToIU9C3NWZlP+ZMQ5tu7mH6o5/upqpLaWxcDqojsf6/JlAkr3dtg4VPHQ4Adv
6xUzalz0DPNmPkuv8HCXDMJFtV5RUTjDh75dBB5sa+4Q8eme6YyEgAo1FW1fARLfnckQFV86rAy0
UFxp1UjEIKd0dQ5gPAA6byZ1HJER3Q6z65SYJITft7+V0Fw2QwVEOBu6nzz04DAjCRMUPIrLmKj/
efAX9N02D/M+pGT5h+/Q+XULT4SweMwcToak/pq48g7jv/6A3eLpZ67FvD5zmgpmj5bZXY2IrXRM
yiuIzQ7PtPD+Hm5Jw/fejV3Yydx0CW4INPttz5Dv0RsONCmSb1weD0JNb/8KfkaAByR/abcy/LjI
B8Bn/h9lRJjRivrxxGmUBC+G1EeSkERydlPjG/GzVjDzrKKWQQIVxgvPZ2k04DJSvh1ZEdpHJZSO
FQaQJRZeotGdDxyd9Dm/8nrFugCYuEhIAv0yA2fnYTbepxWYRjFERXWAGPvZLQ+oNuJmOLrIC2kp
QMcvjrMZOaPQBR9THKQey37Lm801Chlz2Q/2MK9AKYVaq3IVIz8BAVU/jEZXXSpIXLWocHn8mAYt
sCz8QPMEDf0/q/19a+PoYL5TvprM6QZ8oOgercAWubb4cmqwCPsx7ZnvP4o8jBssJaQadDzR7KbI
KaNX+MznU6G0gklu1n+QzxNSxJdcOAx7NiR74blfegBEukVjrEt8guoWY1WjJU/UfUvYnqMHsZB2
Cdqy522FG71EFHF969GU0iH5SndLmzZwipoXNWf7AN9k2chLUrKB6+biByon47gW9KBAP6ZbwkgT
v4tjhtxUmbrk53nmBOMrlr+nnAI3WTffKdlS6uB3gsF5HzIzpgi14FZ97QDcaLYC7S2CrSTWX57q
1bYjkL45AAFoouqzyvA4aLcaxKxzWuQe6a+wsSWxsh+L9GXK7/FyPXyf1YAUYB1+iBSJcM8rRasX
RXt38rzFREu011pDXN/fiwalAFXDx1b7mjeGIaRnzubmMQzvbLjURXViGVd89LyNy9jtUND0yT/Q
TFAqggFacCvZmD8goNBxiLfSzlnDEoJYgvo94u8OdmeB++PBJqsfGGM7e47BcrmPnQ5qii2U7g6Q
tZcZGZ3H6IEbxcPnTXfuvanPvcxSg1eGini5rfpvYLAD6Je80RSzVRrOaAZYAcVes/GLuPxQ28DH
jgJg0q487KWnuOrYkzQg1TOEs3zTPXBDJr93tmjAC5Y1xMptokpi16lbX8cWnQ5g2egcgXiIeeW5
RLzyEAp68Rq05b3c3Fqi05+JHpGC7z85ztC+qJnU6AlQ3GAFDsiAz3XPykjl5v5TnKXUTiadzBzE
fSI2iRCa3Hdjfhmw2DpNskBaCXEN0B+In7JnOs2RC7wVcqhXrpVjcwlVvl7uzIUV9cTokD7y8YWS
UqVN7NGXau5qMK8lQBakcMEcTk8MdaVNnJ2KK8pZmRx29rcv7+PZrN1QS2rB9YFrsG9kHYRaKxGV
FENB2rpv9ZINkJagtQ5J13R7pd/5CV3KlITeWA4UdepXIHKM3CtY7r9tOL5w91CxbLPrZLMXk7xP
cBBphj0bBJuleoh623DPscO7GkM4W8chCD6gPQdsVNurEBxwVJ3tJmgWQdAWe0J8PDPPuKkkAJ2C
2SAgAXYnI0YO4LD7wRRZGsCcBv4c09Mkxgxv03rpH8tV+ilA2qZUAw1ZoC4XjpepfDan8m8yWXcz
kO/XC5fCrJsY2shVaOrQquN8f6UTh9wGCDh72X3mzL7EFEqxzjgbzxoymdpCr0LQpxrY4vvAVtWW
fJ1G2fdRiiXgopUH67UVlmJsFR82idpycLyMfJ7dDDFeTETfsVuMEEm2mO3EF3cUc7cWXEFgmexv
8xZLGdFbpFiYYwqePusMTGsjxxFjehHN34P2Ahnf1VYXoU3ED9zTlwxJkXQxw4MVwwIkDCk9Qsw2
TJraiUjz08RJNL4SFXCcSA3gBPjkTRYGxdwYei9fcuhxiX/F0M5KJ7kWVrLXsEqTY7FKsE2yGE9l
SvXU74zmPRfZzhIdrHQs0q4TWTqVfUzmsWXVI9r6eqmpBPAdzD6HCrpA8hcJE8vZ51j4I44fFPTt
zpaGYdnMUE3mBm56iDTXUF1716S2klX2+NemiWtYXR6/sTAEocWkF65VbjeeBXlmZP76955UKgHu
7EJEIi8vGMogVUaJMtcakj45LJn4Jp73wxYDGIHqV2lpsgJdawZZ6OzX1TyUoeruE8d6xwNIBQ5n
tRpLOdarv2aYUvmPb7nEOHMHP5wF1c35hB1w05ObAa+vGJaqJWDyQylejGrAgD/OdvLQ8m0W7tXa
KmErp9jo1O2e/7fdT7g/o049woYDL3Sh97Qs1s6V97mTXhMxF87qBwlddI4LHyEl2/cWmYnvxDnD
tI6r3ho31/bLY7+sT5jCQuCjYpsHeXPUHQmKw4gUFLosS2i19AD8q/YKUBp9czV+D7uthEVcDAGS
0Cqoa2TCH3saqNHBKx2sxdDfSAH5/xNk5d67LTstUP+YnO/hW/paS7+qsSoKFWiKqsgFvPRJCD02
ZmdefEuWbdTCLV9GSU99iMBQl9ZARqhrKznYkCkU+NBSKCnxAfyQGnFpcC6Yq1JIVDwu5kt1oysC
Yat0gfXSftf3Fc09sctrd85pSDrPiyBVwqis7vKvlM1Ej25HkWP3Kdu1Kh3V1n4tcNmrSs0MuJ6f
Hznlrk0VntSg8951n+vPr89vpDTqJh2EoMvRZAifwtPtQhx7gqguJ8oHN/0D8BqJbv+byJtSveXW
r9XvcuKcR5Yu5tGJ4g+irmHpxS5OebdicB0ih3eHOQNBtbGkJ/kq1q+BObLrgAp7OM3/RET38xdR
17mJ6/6mQD/CNLxQUXL1L32K0zwq7WtR811I5eW2myaqMex16TWnSNkoBQy2fpQiEcoSjE6uO45m
/pVqVSFl/QyxBUcYpzO86EBXkph1LRstZL0FuBhyVKmnSImx5cmpuNETm16Zg98Sv1ULsbkM0eIA
Xds8eqffuElnWNr4/smjSpE/1Q0JkxUVLpBPFYSwKwi45VK9jnAABXzwkOn7DJnSU8ZAX327OwPp
7ZuTgqA3iljAYD2RfMISOL1moomzfl6cfvszL+lLehVNLxD2/Mvc/2fBCV2fVHxVr+TEeK6KheWK
ZvfiF7af+aX8F/PiTIW+WqD8PS8f9Nx9HNsVmOJrVvpUy6tH7C6Os3YdcX0EWxzsroxfH0QyQS0D
9NGkNpMNtQGxoAFrsSd83mOXHLYOqGE4oa8dI2ba07Yt3zZAZfGv7IguAEVP3VWameXAFj3MCS9m
V/7SqacYD902cNZFsRIuMIr4yPTGE+0zPT6yfWFPaeiYge3fqmxZJYg5C7TERFixV2UJjObnvtyZ
JxLFFgiKIMeamNptE4hiP3ZrQZtDWxbPbcywS0Jo9D5y9ZsUcCaoXk8QXQF1jDlywbNyGxNjoAam
v8FKbjFVXlQovYHiaNxKo/r7XDgIQlrx6b3TiCmEFOaZjynClXwzbNXKZtmcLg50LghLAHl0B7sh
CfUDxH7qwEQeICfPso8uneAD9M9fcYuKfzpwpXwgTGmD69wWli1QuTAeUYMr+ISe2E5NVzhx0Px/
XxC/PufBotPqCL4JN6Mg8QpUvnIfrL9rMKkEhx9MGzofglhzVVykChVkC4/aUgkFM8+CV8L8m4dp
+e4zn1SgsxTSykcrpP1bm4KgDN7FsbvNCDdgQOuqYvDcv2bP/uDk5Zwid5U1jkCcAIAEgHXyNsqc
7YXmx4uanNPs7NxilT8yuffks6Z90hgyzH3IjEZWrtMC/cLsybEzZzgUgvzbR9UyBxgXWN5LPlhu
nRLVn8EzdklN3WHQovo+7ay3PZRRazdVx2LiFdHMNdFPCQqZuFPz1isykQ/rY6WjclPhf6k7+9Xq
0kgOPyRTEDKW9kSkW2yvKw93m9+kDwFSQPTYIel5E0kyx56wKV8CncGwAXt8AFoGQA37FAW/1Sra
WUhSQUi8oauqtQxcWCXIEdJz++iebqfXB+HWk8c9t1C8ces5XUxJbP02SmmcxxzLcDiDUZ+FRQwb
eKWAQIHeEC/1Ga1SSKg6BX5YJSjPcH7+UQdlohsz4tt8L7a55x6BjbehcS45jFWReoQjQYFR8tf6
0otoV7FpQLQsLJvbk0bJgdgmoEbeb4oplzi2OGindZsmaWwbI96iBKakguK9gwJ5c21G6Gar2d11
5spoEAWH6WHITs/a2gpy2unP2xH+8HkMahwJV/VBG4OaKU6vJq6kE7Q6Izrp76fPqyrmAg0flc/H
W72QfOeCi7kZFCY33XWxbn58sxtiYpgExR84pg78or7DVU3HtUyEWoRVkg0HpCSluDpQCB1PoBSr
HDloQfX6WlZfgoun5R7kOY8eZKopRFl/oSG+UFcfuLvyTjxeq9SZEOnVV0E3jlDPc6mICxn77DEr
YhhtSqMehHIy2zNYDH443g46YHDqk5IuUgSouGI7hKAYQ2O1UdczdZAQ1OL79FJuJmm6TwMX8rXE
KpTrij5NhoW0e1bYDUrndKWMX2iZ4Cg1MoSs8r30CPC+fqt4aEXGM/tNYTLoHoK5xwGKXhlCZB95
xD7FAU6URPcF+Y0NpMM46t5a7JupS6eFEtFfOdB/dsE0kxmdGFGKzYInExwX0/tO/I3w6OapWzCV
HEQodZbhDzLRSgOo43Sr70NmVD5FFzjxPL8NSImvsPIvMcBA4huuMtTRRDWM2fqLQE73pO0defYk
q7mRsKTpEZTI9xhICAbv3xivYaFLDqHR21SsI0JEEzm0S9ksgCjlf4o37jhHHbR6h/9cE1XdanD+
eOYS/Vq/GbUhVJUstWtUjGJTsCEYlhvVBnVdISOvMY6ouwDyDkSQxLnfEBfdrJ/mJp/eUA14fXy5
ZY7G/FkYIx9oqPPnx0xUfbZoh5QpvrIox1kXMSg1rmIZJ6gVyotO3JhTH6g02xPCpat6EhWGw2WL
YzwvkTf4vIkwdlXTwusan7dulZaNkpwtw3tvZ4YNqzwTmNwGbo38brCZwEGvCR0uP/lxZ9meI8/k
rnki4Z0LdAfhT3E6b+G7x8+gxFkybzGaTzSYyQ0vW/WH97SvyNQxH9vvvhob9Z0f7THqIWp4TOL0
082T/6f/Js7IpA0Akv7qtokEbOtH2NI4A4fNyB9LRr8HJy2yCMxRdG9c2h3GBnWtiviaKc9oJSqG
4RcQtjbwJAc+oykbCyV+nZl/vGqmqNrLaqP7r2ldCPhaedA6f6OjGCrhPGZEhR2s9Ko7aiLP5M3P
MRhhdW8j16/U+3JXtHIOiNwt+bkz2ssTqN8ijT7w3vsVtlIw50hjtyOTQkp8WRPJ6oK0gW0AWr+e
F3pf7gXbbC4BpCO7nJABSqPqoy6Cp9nkUY0JSMnI7Zv8Kln1638XjVpd0h/rKn+Iivu7ZZjsLqAX
QB9urba3EpU6AODe0WV27+kQ1rosLTcBR9fO5pz9gcIhvUWZ/QD6i5l91Qi9r2D9nn0DzHmyi1jp
jNwIVwHBKhoMIVakkar+VZOsJPGs8aL7Wbiq2hiTpwIgC8uDULwlUDs+cxhCRCyKQgNSUqxZBlgl
XCEvHVAwJSB9bjd139gYdyUKXH1QZ404ojXbhiIsDm0X1t7DClA7XN/+rS3WLpF1I7UhmsFrTLIl
Mw3XpSCsm+wFBQV0mkfacOGA+wFZ1lITw2aOe4dWMyt2K7PF7cuUPLtvYHYR8+oLo2VgLZZ8pDD4
Ybwj8GQIsgr9JMJ4bpnR5mEwtF+jruam10c7ZZsagp8D8auAruj3+pTThlXDNy310zIJE2gU8Cz1
exVxo541npmav56cHLX0gjG+6TkqZXoEoyaiDc4W1vhMkPFcZHIoVl0HFfojLo5aQhRTbP9xiv44
hkO1nR6/w1DAORp7jJyVRsZBIebzXysru1sikSCPDBSIvBiOMd94zEDwCjPo3lyQuoUo3L6tL348
6Y9N5IQDs+cv8vgnq6FBSRse0jonsb46YwT9WQGfp+0pzQAlvJFhsPxWsIU0wGhSD+8L8G2meAlk
hyzW9UFUw6fIp5aR/aKepiyLZgp+92YGK1sL7Ftp7ZVGdrAjZEWsDUBvO3Jgdt/PHFIA3jtrwYpt
tYk18a0XyHmfZ5bWL0eeSfT2T+lAB0wG60srtNGCvPKHykgTjegKEzHU6FLXeEFmh1D5E4Jf22b7
OzWTXy9m/Dg+Kmx3zBo2VhIjP4SEUVWWLqgi4Q9mkeYONB4nlsH+dLiL+gn6eeJvlY77R3ElEhf1
7NWKvRnP7ESo0hrg40sFU3DS4yYZcmLmRHIRGjkSF5v0QtXyB61iXQ+m0yr6OBvdWJ9w/b2FgKJp
NLtHXBSWLgAyoelLuMqUxE8jf76MsYTurHEnTIXReIwVHR23OMhjiS+VdCOTahLITgI2hdlBEipr
TD7IBfepEMWiaXdLjYzjmmlMBSZTOc/I7wIQx5llNo1lqBBsMutR59pnURTcQY118f2KVEg4UHCz
z4xids0iW50LT5jL7LTDbIi/+ZNWa8xNFCm1lpuQslxQPOolC3KzFrVrXwfF6B6W+WLGr45DQLUf
RXh8S0cTX+1XNz6rsj20EXLe4XP2ACBcm5Xu5plquLNb0GIdPKl4jRSagZzTDkNTKpsGeOp1A/6N
yYHDSofNiVd94Oklh23NFXoVzBpJgwO+CS/lbuzUiDFCW/7WOiGcq9O+4mmOesv/qyuYjUJyvLux
3h0xPz08hQ89XTVxUbKvJOX0EGCS6D7I6LZu9EhzZOYLQfqEinDuG7YfMXGP1hn0wn/ASc8H2FY5
H0SSDExd/Y1fBmox5mY8YG8m0Nn2M3aZ3/ZcKPXwk9TmmmDg768adiB/54PXxjH6oVG2gzbvct36
4u+/tl8ULNBZHz2roDwgkRD46+qy9riMlblu3EOsJqAuwEhy2wxGXjLRTcjA6zThuQoStDfswyxL
9CKL3DMxUdU9ZH+rBSDd9xHMCwFUzCqLf/RsPKrnRPNcOYeig6kDAQAy506sDmvV01tigKlZVOwS
4c0c4rEibhrHMQf9HXP7uWt6xWgyuIRvV7xCwu2RLphVPfy51YVWp40dTM0w6v16X+yur7fBr/eh
zlsT2EVlxCkQN/AokMr+kVrNNk6A3yMkFK2yTsdBVhn2WGtQnVxTRqXysOYA7M6Tgq9FMA3fiF0v
V+MDawVoUZsDS1PJ9F8Xlr4ET+KuvooOVmUK6xcftXN5bVLWrT/QmfZFvOOyiEgOGi71GUCqYAP0
mrLxNGKl6fQtkyECVbaUJY8k0gjadJ3oN+Q+qAoYatmQXUMZ2qiaQ+F9xqN8oLkiUcM32L4a+0Lu
8pFIE//nFr6+zOHAohWsL/FA06UTIAj0chiW5qNrEZ9+Lo/DKqKQg7QhQ0CdhPP7QsxFFjLMDbFv
MTcBn+N14lXdrVwiyENSieqvIZJRKrFCjTnl8IzPbgZBSfceAoWN716XZpx+2mceeZ4bYM1FHPFV
27UmqZYyCmYWP+CmvAyE4AFv5aKjtTotGZmqDh0RN4sqU07duMFtbPlXAF5KZoCmF+tTXML4JCXP
rpnqTCWFv80CJPmVzTNjyVXtq9Setzz7dDzsq3y+cNT0oVsHzeLAQPwQaVx7pjb2pcy2iigTF6MZ
wCHY6/N2HfLPe/TuursRe1dTXxW8qnUMpOA9bN8a4afQEVaYqp38woHjwRVSFSKbbDpxGHFPH1Nk
RTM1gxxsE83+MXBds3fd6xovTdzBKq75uxjr/wwn3gclSTVm5ZpgJ/JHfwlvC3hKP8Sjsck7kZxd
BLPoM12kbrQx79wZ3C10vzAA5Hrs1YsoGoVwlVilcgj3wIQC1+p74G+Fk1GVxcsLAL2kTgIj8rzy
UnKoe1TML4cTlKAbRgzBIa3cVckS02OVpDHuKbNegFtmNXbBxpM14eI4u4PczwgDT5xjZefo7hMg
othaVzU9MAAxQ87ktxhxWVaJlX4TJ24hhtlwC/VzmQfltmTXaIaIwhSz7391WWGd0Ksxs7FsuWy7
IM5hKnUEYlk+2xNuIzk72Z4dLSM9GloLRXK7vpvuvLhwo1H2NKou62OMy4yiY2YCrDTGyjZHgQiC
O0ucaCOUG/yE0LfgTrBobqFH4RBgtqZKevVtnArJhlmrRNK8qU0DGmrljzFwPF8HIjib6zLH6ZiG
Wl0ck0jfXbapfxVSJiOkfHFlNumV4Lz8uBMbJLHMV0zGbKBInV0Do/53lGgvNCKL0AAFjItqsmO0
eNC1TFOAC7er11+Z1cn1KXoB5nK6q91BL9vajUE8W5x1JvtjUq+mPPvu+24aswCOTSEFLpYTdFOA
irZxCprP5PwvCLTFnO+En1g7MECtVXhx7xBSL9PwO1fOXFsEw/S5ZhY1/KPXaIDJy447YLQHI7/a
x86iM9ZLsK8bovEwql1TJ7LGyKbXqrzH9cdPTm8TGHs7m2XW2JJIFD2dZteJLIAaOpVgs3SPT6X+
9CUip3bxJ49nj54QlWuMrmVTv6GAeBJiBoU7LG8Eb7vD182ReFN7P6GAeYw+DyqfZcgUn6GCyMUg
WF/Bv1heGPQWfMyNzn9hu/IfYPqf7Ai7lnUfEiZKN+Zdx1vQxEFDNQO47LxY/3i8OG4BHyhuJQ9Y
f5FtUVsCp1zXGSkxuUA72AAoMnh1Qw7fBV0AC0fNlMGUEUBbCST73mURCfvO8TmlQ2/sIdVCPNfl
MiBhTccGsw9LzqU48WTfm5MFucivGeTWBSTht2mkcksyoRbaCr02F6BeGkhncCJWY8i1c2XdSZVq
ELsWaOR2EmGiVOCQSgw3YLFMSXf+4M06Hj5FytV2DS6WVs8E7YtJpC0Qy/Ec/mG+eB/s7n52N2fX
XeWJ2VEiRNIHzAXBa5zNM2xLLuGgQ6/augkG5rv0DGj+HDax6XHZuAdLN+S9lLDfVKe1UDTP3i4u
bgHHn4dfCzQl1GKlLS0B9yyatHw+U5wodU6RmrkBdtX6HvZT/bR9V6D/UDGczLSRpzT7yZEFB1/H
50OjsdbZBnRGjyoyNMECd+FMj+eR9fkvEzqe7nB9QxLTWr7O/1n5yUTk44ITHZBRd+/vG1S6my0W
Y3pkoiZLPYkxFCZPp70xH6ZI33ER8I/fJ5/nZK4OxWvVphkOFMMnJPnly+qL6LdumqnyPCzjBhjN
9Nq47nFssPhhJai+IvLdM4d5x3tL8JyO7cjlHv5HUne2ZdDTKb1IWTu/k0fNxEgpLBgHF5zeUUkB
snv1hCUlvbOjaootmx8RmX6DjhPGQgCtKmDBnv4sOZSjaulAuycRK+kNiqh47NvBZjMXTW9FCLcw
x0InFKAgF644cmk302yP3C124AYDc7jkyZKRuvOMmk8BNy5g7nJ124HvDGeWVgSPYAh7MkR+RIey
vStsedjBsd3QkycqQEM9hxmOTNK3KjVDyqSuhlUghqcwxOgWQ7e878I/KTLW2IW0E6j60nwNeeZP
7AZiL9UYti7wFyTr08lyJq41DcuiQ7U5EkSmn6fHRV3JqdNp8+Y1E6+5isTYfdMgof6yg4S4vfXi
0yMGKKlfBJh97jaO4uv410sUDweEEVmsjR2Kdp7ACXnKEc5w+Du9fw/sRvPzvZACVq4yEKoqsi/2
eXjRsSJLCQICF64TpD/wAsAhc++yHNm+XHRP9bWSFP+Di2eBp6cZRParuYhoVPxuIjvLlgBuA+Mn
IPb/cZ9MdwmOBW5msyja7BScUrbBiBhOALavquFyeLHJ+HLtjwZQ1tkQn54Ag1/zhtY3BcObwBIv
8LqI6FkXwQvBvjHi6DJ/Js8TDPbW/HBoHPjTD9p5fOxhmiw1ZlHFlsUA2u9N37z/Dl7tzBmwEtRg
K9xE93FWndQRs791iFwQBJlxmFbX13oGFIvx497iQ8hjZovym0Y1XM5GcfiG8e9ltmklTieFVBdr
dB1cETELG83tmaFrhkac3i8Tm32hao4ySB1+mJKJ87a474M+a6beAyBmM0TUXntqVAfJOrMpIjwR
y44YqmFoBC15iDuHrQS1B0HTA0RZK+mszGEeS08cEd+csijMMGT4iOm4jPKuwAjcajZ2QgAwD8kN
4v323m9F8IbFyfNhqAvfHyq3ApYMtrMVPlpDumHCPbcNy0pzG8EfiIA5IivRGoAniJaxytJ7rsHz
pezsitc+OWGH4L+hE2SkE00FIx6NKUomkF4Nd+fuFkKOlcKQC4K3jAOwupeWxjLNhFC2PMazSWsb
Cm3/UifW06gMD4izfajJamfMtNLpf4E1M2dKnVDoeyX7Yruoo4T8y8vfgd/5mBUHGHJZvtS71j94
otFZumI+PiLkjuEbNPnVmoNFBLDrUOqZy386SwBh3ktfbNWT4XOstk0rujOQWkRWUUwmXItRZKEI
aeX3xn6KM96fDGytzyVpsdmrj328kVixS+j2SWfzBjSfVNkqEbZ1JSK3FuvKo0/TbEHuckOqaAfO
6H2/gd48NwBz1DXQ1ZkeGvQygEd9hE9NSHm7uUdEKv0EAWjyYvOtjoh1gyI/2uOCTLLuY8JP7NY7
JCMIT8wb5kMqUSy2ntsLo/7Pt667HUvcfBWZsQLOa2O8pHlCEdWYXDL3YrP0h7ONdkII+nwdnoSZ
Vyoza7W3v4b8ZbDZ1/oWZEgcu3jLx1qbuLhInYIcLLx8Bp4S2iMEKr4E2gue1DUNZKdLH9fri8hR
8KjuEo22OTjGc8BCyYmANLIxiHlOMFsQzMDxEAX7Je2Cz4apLVgIyUbEej31Vc6TFCfZ/o1a0b0D
9pvnkuSknH8vsqjaoDHXmaYJS39BZ2IoNg37t67FR6CT/f5fvNiIYip9anPIUawCMF3/MJNqSLPG
lAh4CE8UnVvhYCIMfqIo4twfqrp4tmH8Ki+qf65W57+t+VTjmcqYlMq4/kjZOt4S+UecCbxQoRd9
CO99lvnBCpuICugxWxNos5qso7TbYhEO0OByWOGwDesgvJlM+k4IEePak4RxVHlcu6pGKIuvC89M
iSYj8X3CtKOAxOD7cE2kHvsn+nA5BxWhIYNuHixvf/uvA7vToIEjRqRe9pu83/oG7RjbwobPuWrP
HSZkKr3FOM/ArWPTqnRXvVH+Fw0ylm5Py019y+byOeg2MzPs3Ajmto5kYyuh45Yk0dSaG7Q5Q6/C
vIXPej5TmYaJar26K2/ixKTVI2WI53ILyri8ULjsQrskRoIckENX4NT/iqH1HyHZGUp7lie4OhKr
XqFcxPx5R/dJGbyFPMtWY8kNvokUVpHxD7aJKYwCxbse1yH/xhmZ4L5SLx1eXDfYRPeDS383pw0J
+n+U25Tc6cyUETestbM6OYkGKKzp8yPMkcoJemf04vH9Zw45PgdP0JwzzpYT0vlMON9KAN+Qqsfl
DGsCc558YshsxhNUExDVgtx32JZxGeazRDPgMQnwj6F0MeeWg1c3QTwNOvJj4+GDsaXYE/a0dEvy
Axr1UBv6Uy9UtJ/DYSM005yCrSbdkNwo7Tso08HuhNJt/+hZ+nQBFrDftHSzx2QfUKNinlFNYM7s
0b8aaWQlItKU7alXnktg9Qr5Vk2QAHMMRLUo2ULcDakFquet6oL8zkX0sY6qXw/XQWmwm2attUYV
S8bxTnHU0ot2Kb32Irxvk3n+EWBWiJhUudVSdVnHxzKcgvK0JEBZhVl0e29cJR8E/7a2xv5IOkNX
yzpG2VOhL/OUBkZK1y6bnqASQdYmkp0pPcjxE23yn4f39wQVrseiGbeE8KcjvabmC5sZmhAvk5W/
QBxm2c99dtjLXCTl7b4nYuO6HbnrfqR6lPmo5qD0SavZgsgCM5aIBRCymj+CQWRFXeS9msmtNgDF
bFhQztVHUEvQVo75Ht2Un0BZTT+5EKzJVLy3KHds8p/pmNUddWovJ3tV/aqjmpGyz9KcBqVu5hTy
Mnn6rzKrvtqCLYNThLRvee9vlWSrQoNyOY0EOMhMdLTMyJCEjt9Gte0sFmhfAWHdkI4XLHLMTtcF
OlKd04GCpibis6aqyl4PVI6z2RfurxxVa9mncaikioD0NsMBsayLauVEmlZ8xTGBm0mPdhNWcMi3
hTtDpkYw5QhvjdZU8MU9ew9oNud8l83ko7gNKFNEnEHHDTllNQF/BemhngR7u9+FBEzO+7i6OosX
q26/gM3++ERs+680ZVKVYBFNvGm2xZHUJWU52h/k9UMk03MBxPupRJa4QtpWjPZYgrsPLnrQsZfH
Cf+etoCgAvE0d72uSztt9R9iZ+cbP/N/dj8B6ckyJ/R4DVGxdAyIbs9vHJjXlLCzG5aTYiOCuC9d
fOTYbXtmsIeERh/uB6X8aB8Q2pvNtP9txGMCQTiuNeVkhW6N2ZnPfS7KYe84qDl/35bOR30cr/4t
u2bw/ou58rw8PuSL49QaJ+7zjWigNv8K2FaKoiHM8c+VWxsdCDbg7r1ulygW9Z/i+uZCfT39aJtz
m5U/j4r4PZE71MVNfJds5PKMyTxJrO0x1Gn0+4SpYN8p5bRkJavaR/dRWDv+x/4tG3A96kjEU2s9
1AWBbrp3jqJQMX/FfTL8nltbtCbgztoURDKdO9SkFNKXuOI7mb6U/FgoeE5r9nok+yNMErpMEYRF
gVWTG1+SlreKca+i8P+gNZ36OktlGj9RtNzeEyanyIA+xIdONSkND4qCttpbAkom+A8804u4CB0v
21BL6Px7uW9PftITNwPg5PG34z9IJnRzuNprSL+ww11QdOHcLsNCJADeH8OIme7VTkcd4LTOOz8Z
i5HsNd1WoaKVUc+9e8QzrZcJ7lwhdSw22l8EgoGdt2Qx9SS+KvJmukj/50qxG/j0zDYWOYE/U7F3
pA2b0/IYoaPkknCb3ZK7Fa2GHynxHigKY+od23Wd3l5KaicDvOQPJncDoVnMBv8eWQHKOi6ZMc0e
9m+I884rkSF+4GP0rxM7d86DtbNIM4NnsY3987ArYVWa8dROuXGks8sudYPXSe5hOtE49Sw5GXyl
KdzzolFNjVv9p6Mt0aR/YzLIx9esOF/esH/+wlhMHnJD1klyDtBWR29dpp/ipKoeIhIWgP6AsVTB
BCTHGLRhE2jpg/57jfSqcYNW4Ua+gyw8MS3uyI8U9Fyl14m1hJxKErExABVJt+U9IUTDN09sRhoA
vqJKqlAcC0B3bXF766tQzrC8PjJFAkOwkdaMzxYsylY2Qz75h3iGecxs2HYNbOkktIT3h5WkRdli
NSyBZp7pzTb0kmrGo70lJtNek4DOkQCvDZEqI8MWNHgsnB3a9Tuggz6XLhW2QAKV0nAs6PWmqKpr
tjHvtot5W+O9f/Fo3O0/qFi+YXpLUVCciSmXlSyUlyJim9kX9I+o6CI4Tty1dff/O3PjBSYfBcBB
tsRalhdwfa0G7Id7fGpvIxrdsoHzNW/iY0W/2XYm2BUO7iPte6a0BlAgUv7dy7PfXkTYGRy+8c8t
NljhNVv3wpcV+eWspXYiT8dFt41HBkLLOTrloXWSGTZvN9Dn0qhPxrQR7fZkYKnCN900Etw3xTjg
ll7EptACwDWmGi1/qcJnO+5oKE69ApmDHWQu8OJpr7Pyy9IZTbJWhvBKttqQ9t+L8kd+1s357kBC
KqzH7gI4JICM38G5Zcmce7ovMqR/oHx/BEurOxeIGB9GuSaLstkRld/aeaDle61TpdpOK61H0xRw
DpUIMx1shpeepKD6/9rRlkVoVyTHpPLHR8pGCLRpHv0Yh4NFNaPj2mRneQGk6byvK4B27w8D0NEy
Zg08EO+sc+ZlTdXFtFwweX/opZmWdKrut1nnBQhKbdRvLBLVO6uPO3JIDJpGuh1nmj+tODQ30Z9C
Do3pone+HWGMbM8O4KDDNuAc15U2agtqDXEhSqVmhWY51wBPrr9ELO4j+7wa3+8xhurjj65NqkJ/
Ost5kQlYqOPwXG0Z5U1zBg1LCk68EZeP3Ex4aRDL+4wQdmUYG+ppJGVMKJe1nMn+b6/7Vz45H2/K
qoq7kfqR1XMjO/d8sAiI/qYLTxgxc4w3Xli9A4WXIU4Jf3C1RN2nc6lFEke/N7rLKzayV/0VWEuo
Y/DgGsD9oZrY9JuHFMeG1AUTtwNDAyTXeFB9K7OQZS3P6wkqvPDKoPPmMRkjn/b2roTxEBK+26k9
3gbswGy5WGef/0M+K76Q0gjkH8J52jgts5CHksHwQ1waXjPxI+J2igb5Z+lKyWselqnXGh962zPA
hT4GnUEZuFOUUnwJoocRSOXCm10NJJuya86H8NRKjd9Byybd9i379xwjn5VshBofPj1zRCZuOnmE
nJFHdKuAYxJQX3+Gm7L2cCC9SRLRm1N/ApY3Cqjk4Zn+Cy2JOZ4YzyKwjetzuFmx5upiqSb6KkLK
kdLMvSvfECQy/UTx02NjWbmmRI6nwBAkwCWTMWKtHol5Tv7TloiiecjwTBkQ97H7/+mvM5q7lSRr
BSxjv9zVsHG8eHM7D4zJ7rIX00nPRMOxYAzvXlO+8DECyzElHxyKMkSDnuGMLxpW3QkDngC1E6Ea
1eoRbd+ZgjShZi9NVkH7Jig6SYOIW3J9jr3OzaKczCOCQvnEpCQxEdSfpsfTSCG+An9Wal9W1rv9
aloFlBHgmXkSmc4TYGXUY4DK7iQ6Ym3MlqZ7forPhJGv+NrHFAWJoB9B0+FJ48WjANHNUI4zVuK6
B5/t2iM4C6XCPSeWB5CbXAE2dIzGjJgzwj/UfrtKKeYtF0eZctptQ8IU/SbZ9uzpgM+gpJR1SrR5
B+phjjZkbO2sjWNpzUV81eyu3dRa1nxxR/HNGmRSwp1QOd97HCo0N5hbUgBFrGeVA3WypyhORenv
8bDeeF7Gnk1eLZqE+B5eek062DNfcqJf5lBa7TTqznEWT8R/QQjkPTrbdxokT3gzx7HflD2xnSIk
QHzRD0RPd6uA7Nedfm6OPD7syfZ019yNTZT/udrQNEUvl5EuyBYlMXTmI/q0tGpXl40am42YoFiF
gVkYXIH/ZWBQfdtnbVZVfCndykHweGgr6J2lB6hY6NwuOtdg3uObXVuaKAwMF6oB8Ps/NsxKXKqf
61KheeeWH/MPyur5IG7iSBUEFWvyb63Zxhpnvx5/AR2UiEtCt2k8FSxaNtkWDjLUM7rMeqGWONSA
GCNV9eWkdpqTeXlRa/pMw2qAHe+w6K/7tVjsOp7K6sKj8k8jbLrSDBRVULSlggHxJhhObLWq2JZi
wGfQMo7scGh8O4lFlmZIXxDXGcnmya32I56zGMoCAGu2sNKOyxYlIqbYYmq0gsL1Mc+A1nOMAQYO
J5sbuExJST3kY1uSRV1Hh+A/2RPHG3N2LtVTRKG2SgUsoZdMnE2EygZoHWdZAm6fIhyJcGXV8S51
I3LMn95FeXiqdHP9I4AV+s4pngavlKlijXh+sHxuL3sm7qWnRz0zZs5ogBhGvfNjsiJy6OC4UAAv
bgdJ98zfeqW8N2L74lGwa6hWrjeW0JhnpjWuwxUK799y4Ftc7VWAFjrpQB65yzt6NLpZj3kZmXAJ
p0icA9pzTJ3axGZ0juBJNBCyZCxlkVXnV11HHzhWl7WVn22Xn/6mZ6FyqDqCWggPxfIygqkK3SjH
hIBV/H4eqYJ/iLTYvHr3r+EKNBL1nR8QMMSXxnkaJUtK8iFzGYv7lfik6AYtqbHxwowgweLkiwkC
Ff3+Q3hE2ru0v8+cbIi1ON0o3WzqNYArRppjDGUVQXjDvD+9xVstA6pX7EPVHCmhBMQK+veYkma0
Y9UBD04gvXo1ylLTT1hkffzVOSIKCIhzGfGp5kf7sqx+uYicgo0vc+KIPK9loYQgwj9QbUjWA2BK
rIqQiZ0th+ua8/ip1osVUv+QVa8Liftaj+e2vjpOxJwSORv1QtjW5TBLlE+wpdmdL/WhLCUG6ZPm
QocbmweHUbwOg/rINmubQFBOOgRP/fKgqy9OejjpYEbCtW7ZiH2EtuGEPUF4Ds9xMPm5xe8pBW/F
Jeoasfdb3yIMCfhDrdZTIZORT6dvqQT3qTsnZS+9h8yVx5iwZEwEEw2GBOPiZQR2dJJTpYDazod2
gqmwPjQC1z4JBTpHeRXGj+Lq4BPJ+s4a8ZIN1l6HDyBwTSqKQmNMVQrjipr4UmcotvU2qIOwG1Oq
4bzFcTzxOXBOSRA9U74j7m+VQbAOy0UIAVUYjgQXLSKBCtduLJX1WLzbYxy9MMOICJflpqnThbBv
CtolTYULNoK71LVm5gFdyKJUGfZKPV2Fn+CzANK/unXxBfM2hWQERK39ybvQxakIxR0Bdso3xHOs
AXmgewXZQHrAeVkpPYdjauHuiCr9hIZafnbCCkp+SxMhTdOHmdKbbT6H/YUzLXpBC6rEfqYa8snl
QxZcXrjcH7bjxQylXPTo6Of3VOk3VN+xqqcKU8sheZt6vw/xXUPzj2OuaA7kggDX+2vttFm/AZ2X
jbs5NmgIWf9aO2hJVPhJlvN9nvzE3CY5VnYPSxUT7ove66ER7zzhUfXki2OKFZZESxioH0SWx+s2
Y66T8PMDdCIbCcjvQUKS+X5I3JS3fEnTXP3DhkGETOCWLmaR0CTMjpe6R5oVk5MX7lSFnhmH0ENp
31On1e8cDqCcjZ184mRzBD58LgPh+KyXPlgrinKOZgfWVI4YehOlxkdi96ploMZslIP962qMtJKV
6aOkplvWsBWgtPa8xTAziKWoJ+fMq/C9HUoXmJIbcShIyCXZx/JahZgETjtDKsoeRFs5ymT+LabE
IrxORaX6f3HrKtDXlS3tMO3DBEpnpZ5KJw8ElgEaNGtL891mhqn/zfBaenOl4fEKSi4nJXW3ZA8g
+OtfofR8yMNBH84EK81SnaCetX3ZsqDjRV7FYRuvwZaFrp5+1kOkIQiomnZOxAFPHMXZcyUh490Y
Wkt47T8uFXuJm1SDLI4WyRtATOFU6M9B9EQxUAbNHChsEwn/hvT3ZsrupKMjCYYbvlIKIVxbfDvd
lRyVym7ZQvDuZ3IdnsywZ/iY2mHlQEtTnf945FvG1O5m/ffErtRW+dFisy90dptaV0siIzRBKWSU
e+2Xw4kIQZgzzO7RIEXml4Rwb4HEF4gIhnEr+Dws598lP//m/LcEiYNTy6K/22fB6wR+pJ25EMFQ
NADZ8VkVZ5NInpLn8UdoctKPv48EUEojuJfyZOBr785NdRtgn6vXVONo/CLuuqMDmvS55UE32OMm
1GMzm9ZXdbHPWPGah9dx6BwrKuixTlTBpfNQaXsgnwCKjnjn6uX9ayysqRzlaJgWUKWQarg9Zzlm
sir29SxXI+IFj2ona6UeJHo2UiXULz04BtGFvJphByGxGcL7nRtPDLt+wqoAb4QI/IZDdaqnrqPg
yWf7ugnBRLOk6tn82diclFNCAHFk9uYciChLFTu5Rwq7FGCkiRT3RQyHzJJJLvsBE6uGHt0w73qE
fTBRfUfftxnH4DJx/9xbzhmBrwPJlTwrLPIYZ/wXHpkKnDY6Ok8yFTD+yN8foNeBnKK4p7+q/hwc
vEWGmpWOdEAuMQ/IqZ5laeDVLKOBkB2IGnrZY64BDABiOJSjFcf19B7OlpRxbyMwopnsIm78zgkX
FR6Tq5MMgc/5NjAv4VrFx0oRNtMDO7OmQjqx6sApyldLj/gmDJTTIT4o7APue14da79BbYl9VJbf
d2yWViTrAfgim+AJ7F9wT1Co9E7cRK76jztxQGccEHcQfhrzvt1hDMcF3iyeN7xDAfjOIpXTvffq
gMLo5xq2m1oEMVHDsD6dNwNW7y18ANKXnuc3uZDm40DfRICaAIlXf0Ru6HEkJvT7BUczmEL9CGvG
JcFDunBK/khmpTkN20BbniCTZYTAxRPOl3UyvBOi5ryrbOJ7Z1c8dO+mxjYAIQhzcT0TL/3/cvz5
o6CGNUPOlzDouhV8YuXCkBgoKkRIkd64vHY3ICSEfT7MLz2jdpUNsk776Fz2eBfS/S82kMfQhJV9
1k48pJeIRwi1wcgMZDbUx0noivl3TiI+yC0ea5C3yP7Jkkpw+71TnFcQZT9RUbAe5LL6Prgo6Yqr
Gv+v/vFVbpvCXAtAjk9LPKnzrojZPzVnUSLPUdlhRQ1oj7Q+DJu4qS5aKtHNnOPLoKsgeks7x9/h
xujyPyAGeYl7XTMzxCfDYtX7TXWBtaGc35H0Ba+Jnqplhlv5g+jrMjJHwuuAHvC5TvrSOsooW4Xs
A7AlEE3fBke/QmLKJUAx0D4rFG202SsC1Bp9faYR1ncSd6PJNal17+jGGBLMEv1VPx66vS08seJg
GChaz9K82gZxhvetoV8t8X1FGi8amK+xs4oEYSByaKz28RE3+9Jx0cjctkQ8UVgR2L8qEvUGu7Hu
7p44V5qnRb1kBs7ha+elPU04yK2aFpPVRSqIgAkCaId4MWxvBD9U9krALlLcNhvnk8MzhnMHedsQ
ywlUoyAYibB34JzzGPaclEzxtWxVfHVpuw9h7bT3d9rz7AbOzi0Hc3VWJf2mGIVvNDRWmIxfJhlp
6LKg/bAcArG3SLJen6VaIxFUwL7DXV6M6mS6LEiFfoQmoX1FpAFL9OszjEV1X29v2oTRds0PbXmN
S+NbdAABZnrjTn4+Pbn900zQNJJpQUyQKjcJoE0ydjvAEYPZ/ynQuiU1IHaMlzRoNLF29Qv70ORc
PZ9BsRFHAsLOJ56fAKQM8Xkj/XJmPkFPC/rCu/01RYavO//rgdwc61XihMTXzXgqjM7BZKzBcAgA
Htk1vNzXmh2lmTz5ZXdCiP8EiLdvG0QasRoU+Ijhx0ZIgxsIbsGFGyPVDHaocC/oX2oQjRyhznJt
SHg9bo52Jhx1UCl6dyc2fl/2KqJTTnohVKhJ5Byx5F2mszCfErIbbP9SKS4lOKCG0c6y/E+wcAke
6O+gsnfm6SnD/wyDEep0T2iZLh50hNV20bs4U8J+PCQKiXMIj52DrvVCA/4rHDgxzoVH+TqMTjPz
Wsv3/JzNLokh2+DE+5clAAyuOYhm7kkxgqyayv+xfycJL49wu3iugDBgUyD7ghsvrTFcBRgxiBPH
37kWzg1gpJvZqCA1wamtZeFMn6BCF3mWNOA9rCzsUoFyLaP29GLbGKx493aEKQk3S7FNB8t3ZWHm
vH6iF/wFFg7p53TbQfIM0C1oDC60PMa8RlBkwh5V5Jhkj1VDn0vNCTTsAb7V5cD44RJG0OFUZnBg
Gz2CvLkqxo08jfi9fHxqFrG4DogAXl7zyHXrUVS+mUsFJQTlPdoTQnUv/xjXLEswIpQ3tz975+R+
0y5Mv1t4188uXs62h5lOJ2Y6dsNvXRWxdUNpGcYbx3nP4Xhj3M4aSnsiyWkRwiQZGkQGet0GglTG
kxdAdp+1GJa597PpDuoYfyAKKXJorAHxAZLwZ8e1Jsv/d1x7OeUWFZGpLjVaHlw7WXZKAtQI6A4p
QP/AykyhKE6XFlajOiKmhJ4SaO9Pue6syIB42aeshDroPCSpM2c7Q5t/3oIg1pNxDWRkDPcmu/Sv
urnirkd/XLIk/8o3xevVu7fNSwwbQ6P/+0OvOvcURjZoknC5s6ZhPbG39xPB4f00O8sxPgvxesLV
KQWcKb/0keeUrdokQGP829ux00clWE62FH8d2HsenjvDGQIQIPkngin2O74upLQUk9BSyObpKPUM
hp1jntItx7L4gji2Mi+fIfxe7dKeJNg8lh/DoSH+hqPig+kFNgVc3ZvmxmChmLFn2LfnyowN0CMH
MFIA7c6iiXM39rTg0zFLNuQeX1Jfa82usdJZ04qKkPVCBstWVUDyGjcqh+VRb0zAx4xj5+bNQUSm
LEx9Hp3T3a5N3WzNhF5QQkfYb/ggH9DfyyGHy2hw/yuo39jW6ZdccMyhuHZ7OkrcbXYFBY1cZfh/
i9My+/UwJg2au+EPf7Cj3ntN2mN/81LXwOHaN5MJUBQhw+CPxZq58CWwZJs+GmuH4BIke7v+74r5
5p+axnHi2TMje9QPPow4d1G0ZxYbEoFQr8Az+lJ5BdjCYAMpe4dzlPp/jOIXk7tKa8UFo6I2ZceS
Fe+0J7KpgFBclnKBsn4TJ2UjCqtVrJ5jYp1ijWOlY4qRzlzXaab+3J/420hoDWROxoydxpYu5BO1
+JEpbXm98rwqEJzrKXTNwlEVUbrRXkrbrWGTS42biBMmTCnFzlcnL3b9iR8r8PSDmnUSSmpY0vM4
+mTYFBGH8BkjYVE96NTGhOg2CfX8rrOt/AySC8h54oLhAr9M/fIrvWkluNCQ+CPvEMDUg9Esnvis
vF2Iz7o0zptaj07yGY5eZcbhuFmCtbMgzj83oe3jTLK7t+hnRxfY46LmbtLYPsuUTFOTVhXlFeF8
Qr/rPH2WkBzrPB2zYpvIIAlq617ca7wMDwc1ZeebVl2FESoKqDw6/cBFSMIO8w4gxrK9ROkMVWaV
k+XkG+Ne8Blzx75BtS/GKV0o3LGwvKTogiobGOsMOdY8mjUzZ/XkHSTP3RSh0Cel1jpF9YnlG0hj
/C2/q5MDQJpNsUSWlBEL0pv+LPPnHurTbjmEdRLwZdjasUv0E+fwNtNnMJvibStq3i5qpmjqUIRG
w4UiKgShh1uhSdcHtkZiC+q3/hYxJJMF1GiiDHG/gOrdBLIuJyvjAoy1Q5ZbtbzIydc2VLiy4Zo3
q0KMfHjm4WPt9wSvdPNxDGEj6yl4N8CEkaYemC2QFQ2ZkaS5+RyiUNYvUHKvwik9R/DAng6GcvcY
wP7pHZXZiLaug9UHuGOra5lAYT1MR9Lu70lUMV/YB5MNtZkpkbHA9s5+e4VYJ5yGZUxWDILXLWKS
0QqEvQBR+Jv+52UlQXy1bXU/D+/RBVzxoVwI+ZNPTZ2ooJ/C8shKldk8uGJ78x5B8JpXeyUkFI81
jBzsW2ey8QmOEaqKTpBKw7nuS6plzgtUHpCTLqRhwWreDYb5Y9sOSyy0muyuuGkmg21v5lFPZzrM
Jmxm5wgX3GDmEa868wH2aLi2+h91p8j138necfy+vc5GMqQ+A3ajODr6y8X3hniovAWK5ivepUnO
lfNRYahURUGAIe+j/kZ67O7EUDuofLDO7XfmNcZunuurjtBIiKGo2RsbbuODUJsDo9rHnv0scQfb
m9+o/Gfl2rpdEe/9uS7/rb0NS8zrj02dM4NlZ1yQsJWpv5DP0mwYCxO16ma6eDDdEHOLhGJsP3g7
IuH6/8HY69qhDYTSR5dU4WnlXtCMDy3hUZk+EpCCuUTh8utwtptOKnObv/gPcDTUyEcX5x4oTQe6
4SfglVPlUk9lWhJ3j6P7M3q8rVqvvl5bKSF2u9ZqFT23+tyLkGwRiGjPizRjyenRBLWDK+ZFPv//
OJF8NIP3pUEvNmLWGtr65pUFxbnWdoP44n/4c22PhJ+u7tHbIS2wfuLTzAixZYd5oKrlFUFKkFZO
mdLzYQPEGwJitn1kGNfJpAx1Xs9hCnK2ZsZG+6wgE02gobG31O4wf43tHEQAkmnDhyu6mFqPhJNp
vCJ3iYWwTjqeH+NnGd1vI1KZ1uVhnb3EVR2/THzDDuQcYufCSimHh+WowVNwRJlWmzkleJzt++mj
5wpTKbsYYgHZGIwOemEoc2/+auCck79L0JydiYF4vE7lcbJMdxXceuIWjJ3BTPra1sUXkJEMqB5E
46Ox1BYYh02eFc/l4DXL4/swBqMdkimDAMb1jSg1/ErP1FNpRZrP7ky82lixEFS1Z0YsBVVzhq+N
Y95YMzYwNxwF3pkqbzdcdkpspUEwKSSedhcvv0ev8uCVbHIvDSyuRAAMMWYFIHeSFSRaRdMS6Fex
8fZLhNaoavWece0QoKJzXWK0E4fVlq3jOSRkr/bJYb296Fuehz89jXowtvFYV8loU/+zBPe3m7HO
XY+zlRcdQpDOVzUdtvTqhQZsrjCfPk7om9olqh9PbHGlNpGpGm50nx6L8d0EJciz6JBImHxbWj6T
OtXolWs1GZWDSHwIAXvUd5QcmQ0Z23x4iJAY8rV2JJilGtxHNitZZtNq+A3ltJEYwHk/dasscKrw
eP3a/ObYmzDzN9zV85AsGCgBVKt2Yka6ayRstMvRIDh6vM1hOq+1/yRIM3gQrXtAom4Yc5hcHPf2
Q6IhMu46a5z6R+ZyoE9VzYLjsSIG1Ef+j6GP0zu9aCGbV4igFPtF/YmEMofKXmYtEUtdFXvT5XrE
0QOH91j5jssPDb5TBmqh8cxX9Fr3kd9xYLk5yOPupYaAeEeOXyXT0q66bRjOS326UyIHA13iYbus
IeBLyCUorZTN9TzlRq7iEAQOq4zaNoaTmzscHjK32ClIKXF8l6TTb/uD7nTULzZfPZqFAXwxFrVk
5c+Q9iWtSqkF3ZXuYXVeSIX/KK/13JGh2uc59t3TtJRgZfSucYJ/SEC9NELmjp52eG3ZzE1mxyyC
XMXmSjLIpItY61fNGpVna45BPdqSYaQyTQCl6/4MRL3eKl6PkAk4l4sMx3giU7hgiYNTTIoTpoPu
hg8ldNtzgdKoR+52rvtD4al2+GLb1qlJnQVQamiXQll2GIFmfvnw5dAy5bSLe79dqj7xD9bTTvQi
gySztxfH6d+EybBz9pDqBQsVdiw7L9VeFixUyDHo4HxZ/G//6xgemYDm61ds9dE5IyTiKb5jDlgz
cUTv/6bFy4vqWjfTdXlLl9uHPcClLbndmW9X8ATROT896VcysBeRzhhFM6peq/uCp/X23mA5bIqG
2GWRKYFCQuJ+ln9koY5JORxgzgqaJDz44arV+vUDQOXT1mKejfmLfTusR93vCaevIr74XUzEuNRp
RCyUMngPspiIxhDi55x8PPbzUIsXDuUJZYA1tdsHCqMtW3ySsnxWsO8Z3tT/PKa+hmJN36eJf/7P
cV3KQyx/JOwpH1J2HtSVHU0pK6ytqSrJIUjXYuqqWAx+FVoE7e2ffODmyNzEyAgQTmtIXch60cIZ
y55R4JcJtRRwEUQDZTdcwBuJIEQAhX8uo7lok+LA4GVA4p2V7qPNHXXy9xNzwP5Ey8U2nzKlBAoY
8yKWgcgZcS/jdflrFqVSPdLQvLAH7Q/fgzWneZzvASmsRzjx0vfzKYT6Cr02QiQPuMpJuhX4vH5E
eFr2uAJLd0U7SZP5YMTrxKhtXW/NIAX8Vezr7GNwJQ8x5CJ4kjLd0EIZ368sm1vPyS5+WFAF0Tzm
PvxplZRU8ZD4vXdQUuiAk0+aCz6dnlIwFYgwHexnAfkkp56LXZG8fp0pKIDaPLTjDHt5oCqChl3P
BKSJiMKbUpbpXsStY7dnyBWwzMBHJAjovB2hXFi/1zykK+RWcrOqdKSPHiltGey+BaaI8v+co47Y
5yLUQtg1KUguWJx2MGR5Cuvg/SMl1dawXji6hNWnyASu/hA+JC1GSu3LnFi0xOsOMvqAqxgq3hOJ
H/4LWc96WEpqYVX90ZY4j1f7vbnt8kRLh0jffcMAltde4dFuL0at/qT5IrMzZV3IDf3Xw1WLNgG7
p1w+EEXUrVsba99FK2cmcjHQS7FW85uN2WMOror4IFDi1jfNf+dzIvj4wwhjeBhj+n3BIWZNnndn
itJ4SWY3rcfMKNayCKt1YnNwcbyjVQR6Wol2EarG6/HFNrRPoP1P4nOp0rbKx5lcVuxenWpw5Zw3
sD5vAPSdyYxjUit5Wc1FZhE0Im9Tifr4MUU3t4Eo1Zd6A9UDkh/93l5go1rgGHBChNEGnqC7uJWf
e8sNjJONDOzpUggIi9G5PYHY4a4rDlynp4g1CWRnsXyJn/Bv+FSbdD6ld4lJjrEnWyehDGupYCu0
iXQGMoIvjRECj9+oJoh5iVDlbz0HSsLyA+KDLOsWbL+MzspTyyjMA9kM+IsYGo6JU5EM9kA7ihCn
IewWuipVF0MAeOPnznWpUKdXREMP+WC8yL6D3dvJQRuPdrxVFumaE244haHyBOk7DtmKIPAR6d6M
aACg5WY51/09OQocQotPe6sjNMSRjlXJ3WS7bkiNAzBo9n8YW7+znJheXLYZXjGPeYru3AZzzPN4
MQr2gs4PFli5/PIw8dUKi5WHOTyIzpJ6c9hS6MASEv/7YDZHZ/MXf8yTWtgUG88RYdiRj2+wYqPx
1KmDO0lRRrPhuHVJq3lbuAr7IWrg8wZKoM0mDJhKdRSNpWSXovYmCFq15fN2sNUlD1TKXqi7L8bW
RXs6Yhc/FGNS2nhVWN+9s6QAtlkNLKBayYNq8pKBLcqy/xTPUgAW/y9j81u2rrskbmDNSve7obSX
v24/dZIR14CtaqMq0Awk7bKgD0xIAbw0VGIMKU8GoPxtfFCt+WNKgIQzCM2WGkUx9Y1jGQZvojWB
ZmdZb5XtSx7QtNfL80AfSWDB3tNjwdMlk1yLjPjufyFPKahVNzurwr1KS21kyKHX5dNdu2G8+u+e
XyS4B9Z9QfIc42AigQ6Ss+Q4+caeXBewqgF4qNdkajcqGIX4xPgMEh3oSl7cwTM65wVxlmauQXa4
kfzntxUICPOluTOWAD/5SlISUJMRFiBvvrYEUwoXtSM7iWAJza5n8cyHACGsFcQwhCHIUW9U7W6/
sY4hL1I7rlJk1aw5VnX6ZXXPTXd3VdJpHitN1nx+Br/YzIMNqgaoVmVMdd7rHw57Fy2ahJ3WKqPH
zWkrUCHK9+yJMa0c/aZeUF+AlWckFub2M7SIXOQPbPGgQ1CDEiJScyKBLUtnEi7F1YTg/Xf81iCa
znkU9zybyutUf8g70Tj5metgB6Ew0wHRRP4IiqoNy8LSMqu2FblJXCrh5R4pREmEYynXT4VWvlnF
sRsKrzqXTlviTJhS37AGh9vSyZ6Rhc8X++cFplNhOGpnoT2P7Ene4jri5Y7JPzV6e740y+diEvrA
Xq24XpHWcZP+P495oSn/wWv8VcN5wPhVnxra91On0+zkm+fgFk1hytegGhUbZbYiGIkiKc80EwUq
odsptxQ04+KPkr4TC4VgRUpZhpPWcdqmrBC0+d95vKNxkDksjPMhQJHwDkPeTkz6SUPKCbRxCowi
+KB7NywlcDsZzrILL3QtY5su4wGgbzEZwYy2d+uhMrelHlIlJ8QgxknR8m+HF7sKLBCRkMdJ5iBp
sIPlYsNxnukU4J7gL+JAFVhaUoL5VH07v1J1bXJeYBSUr/k1QDjil7i25bYjya6dNSUYXv4lmbJo
hWa8k4tEuNJrUEEwFfm9Z0lRYWIBjKVCE8104eGL8QfRUEDEgskJO7gUM8O9b8qxSm/buLKMCB3t
HFSqL9qyH95Fe+XJrQ/A+e22ZSry2wVurvIk8PURLujyL5dlqVc3Yz3XEXbA+Lswb7GYJmG6kyRX
t6y7wqbwgT5udPJVclff8dJAWenT7b6lhsOhP1H2Vn9E+e7WZJOS4nVMLbSpdQC+tDeA3YldYZO+
PYZB6Kup9Fi/ZqPvIzvMIE9fOa1S8MrezvCBpHTIJ132sp7eIpMPV2ZmrbR2E/LyCCqqN/q6Qw/7
aY7iHS6/0BMUPiG1cgUNdFW3/1yYt4AglY82p23NQAnp/fK0445mgscdoGrlP9uhCl+ySac3abxO
4t9FP5VsNgxDKRl3nrP+xJix/TRYoBKbZn7QlzGciontz/KpLxOOA1f1Q0PNDorJs3qNULTJZur+
yRYP/eJgZ+6dSmn3hLEbteEyqtz/J1APXulb6dPnZkrXFgWWNO6YS7Ymgt7i7ZgeH9X2hkJ4oJRm
Vi9ufWbv6URBSL2AU/yxgF1TEX6Xg18SHfJ6sgL8IESTxPeHdpOullu3VR9hD0GU+Z8JC+/VzF+m
zrAKksP4+sOVuQ1IwEP7D1Ea7SS7X/npKbi18jQxf8oI7IaIVZoTSnpnvpr4ob/WtopMEw5LqSuh
JRmoiJN43haR0NTKmbWJ+6Jd9n0WuLD/9+oEdv1CsTG8uNWbXySqMFTHZajVsvtSF6eHj2IVNaeL
/sF5g3KqHuouZUUoWPdz+uauoAMsnGVS+h0HhcydSyVMA4qGIPIzq+uWiCGMenJICPn6hhNcYPB+
Q89ocDpFWv9XGzDaY0FEUZpAfGEsw3SetnB0QHUeS2DcNNhUOqvJ8n6FpQB6cKFl6H4x7SLMr+gN
LNmkQJq2PlqJqUzT7mOvGz9xgCTUXFCZebSYQYPL4zhUN1hDC9udwRJ7yx60fU+Bir9he6SJELt4
IjXvqDT6NOCQ8uxuXGKrNh6OwLj/WgqcBrbk2J3hshWjnTKSX3x72k78wtO+34wEgKMvbl7aZYLR
Dubc57phc0eR+MpDSzdZ/txH9Yd6isSkFpA5+ySBCHqW6WgPsFYb8OuJM2f3cpRl0ldOAwwlEP+w
YHs5IFAAbczkXvdhATWpgL4wbEETPGMuqwTck33Eluc0Rv7rhPU9oWnjRfCXO75PqOtx0rnmRcpw
4vYKWhWqnV2jyd6wtlfla7bFRPceuoYOS1VasOQcxFI/Tf+IVZW3Aqi1wdAV3BqZjNAwvfqkyOe8
fFLCNWcoxcKS29bwPROruFnIRNbDpgNTlfyzEkPdgrA4hhODCZf2nQcWioe+sdwDliwY+q0H6nZF
lQdZQKEANBzRUMqFgHFh7sa4cofa6gh5gFq4qqcXAxTpS1oMfBKvETkf+RaTqCwaJcznSmgHcMad
atz23sQOpgYPtFRT3m/az/7B8gUcke8jEXLW4qNjeYYVxL2ycbxPmxFxRHC3WTwClxCVxObrVMx6
OciZCz+ioDLPZz0M7Whf9AwUyy2Hn6hpiADHwLjarWLiGDDzDGMl8XNJuTW/V/onTKiL5XPbzmx/
rwgefNK4f0ddEWI89vXKV8PhU5YqKD+ILJFeJvmI1OydUwFAfB75EzqknTep0GU5+uBAzbcZxiFM
kAiNCXqhbO8KdM2pHMBjqJAlsFcAcm0v2wXxNhbUOWjV2Iz25E2u5ctXM0S3EISjuPNlyMzjPNXJ
eqKzfJ/V7GGECxBvWOUj1xYNuxPLdLftyFh3kHeEzvyxqF1lvWBAOpJIMY/lFD6D9xoDUDaDxk04
89/7AfqtdPrEP8v7uEplSGUXqtZ9BKPM1u42QxtbQmIa97OInze9S2M23HWX+BT0XWp4x6qdhOaz
aEzwjSIZhnQCn8LFRe3STZ2pM3FquXdBzOZtJq5TsuKXnjbcUDtIL7ramDORt0LMkjXvpdIidmsV
1HMB1Tyr5wmMRJmJRedDmCg6S9r4i+8URBIFjRm+5EJmMP4KaJZxndZDbkPaFu6NgvOnv8EMMpU5
nwA48AIq+TJTYnmJYCBS1PmqjksEXlLo3hKZKUp5SKwAiKCFHNJaYVGda9CUYBjXe4Yzl6ZaSTuN
Y68MluUr2OCX9SYmKL5M3ZzKwxwm6tl30mQpGBYDdtMQNVQACJPxbmXdzh4lJuGhAPR5UkHizLlh
YhxWrjh3o/+7DsllUx6R4FCXX1p8APbil2AMeCUQUF6FJyLubwwY78ArL9INSEG6BmYlHDrR9+qG
p/aeBWBOC3dfQCyKtBbtPYueKlZlgUZwPPvVwL3w7cT58PvFKKGbyrhkkZF7+59mcskU/N7bAEzP
EuKKJwmWTkm6vfMqQtEOlnCSZ0HdyVhTJ9IENDkegvJTn0YE/S+NDZPnvnYOlpRUoJfpgYS6/Hjz
k/v3F2d7BH42+2XFC+VPKuGV4jdIgFR1gxju/N9LUYRGB7NdDTCDlxmzfdwrALuSRgiqRgr/CGUe
OWqJZzNdQ2a+jOxtmdH7IKHT99x7Qllg/zBf//CfV3g1lJfPgyfNbwKqbKO3xvgyTumuZjnWwsM8
7ZxJuK6WEw1Z2Pul50qB7kM220caYaY75zh37jPrLDcdm/WnYKl9oTLaGIypgpNJp+gxODKFOZXz
GjxJ6vVtDTvI4hCT9ecR+ChaUIMiv+MzHfR0DYLcsL/QnU/T0a5fV2kvTyhX5UpAEB1Xs7sU9prY
bSh+eQEutxEnLXLwNJoW2jcusL3576h/5rZO4L2LRlUE7r40t9qpCEz9S7ABHV5wzFahEAUyVw0f
GO4LTbDzMG8tmkYY0/3kGQbxPCWeQgG5DtyRBZzn3CARxWDuHmp08Ms5UUd9G1xoTSSmlMIr529v
Ap7aihy2ZiowVaPD/eJSHmq+fP6QnMYXil0uW7frqcVLIw4vkuUbjyaurmlpz80tpITq7DnXm79p
JN3uN/Bdg/SDWSLNk07nf9/oRaE6Ainbd4ynRn17LTsJsf8vQfI5sjO32uLxsgLCaFu94WfA0Tsw
2bndsGbZlOssQaFUvRmjaO5D2Q3s3P3Xtc0qQMlIr76+SL5j/dac67NE7f5Fto8qR2MUc3hvFYNv
+qfffHWL2PolILkx6JcXPw327LnOq/W4xFI+Tg2gy6JL3ZiARQ2gblEqr+vTMZdNAYI0mKmrsTOW
+XWph+Yjs3vLvf9GDttIJeB3iFo+ro63PLT6wTSxeO5Nfq3FcUxCdkYj34Ckd4C3jDxvw/Q/yhr9
881WiMgZRSRr7GhCdPixFVNRe54sNQz5zVNixPLA6ywj+iBuZSFwiYcR+D/lJ7RtHbVxqBHOrInV
1cvFTCWwur42ReWvBIn7JqlNG4uN3Zz1pPGxVOBQTaAwDlcXWq9QiB9MwO0SA1xBu5YxheFVzkCr
Pc/1J092Aw8DWTyx1814WOqVoGCOAvwm46GDvOtRgr7HCgt8qm/fE7W8lAcyJ+PeTmw2aq+CYo45
oeok3LDwnA5uH/kyRlFs1C4KjPHKss2fFnEvnOYsc8pi61B68Fk5ba2VZAcJBjXmjcFPaMHrl56X
s7d3Vf9HywFYTtk5Opprw5TH0tNJkpn5rAC33uWwCrFoWfgME5eiE0yVn4TMnuRjZOdLd6uk9sLM
YlXshiYiSKeZluM5e17BB4By1IAVdsiRRgEIjHPkGUBGugkB9De/kowffupUyCBK+wsL7YtN+Nb2
9hVaHeYnf7K2D7tp+z/TY2lMkcMJpP0jZr17x7/Pde1/5Rij0OFla8n6/vIr0PhXoip4JRZGuJT3
jzp7HhpTr3Ci4+TeR25sZsutOpPRtH/hNuUtIEHd027/3/olN+TbmCarOvG/fP4MDdE0uxXIXtMG
7ZcAW5wDEk8or/5zMEVyCJH+hOr0+LvoexFz/QSc8fbtPoqnv/wokyG4D1BXN+5gQi/CeWOh/HnJ
1AVcgAazv5LnUPesTJ42InxiYGU5xoWBebsTl1CMhUjTEikQfmt+MOGyWmQotLBGlXtPjHGiehD5
rQqvAhrnaRbsQesHeeLzAzwLdFgkkDLvuWAAa7AGHlvbtHUfgXCefydLlgtM7YPiRU6zKocicu+V
dbtiGHNm/fCHusjXWgLskMn6zIYCK48qo714YUVESNp6ono8mIt1GlCTrWGTQQj1e8q8SW/LVhEA
3rt5d/Fhws9WWZi5ej9mguxj3GzkZZOLTqN4UGRLwv/DzjSMwgbSOMOhZ6KkOQsvNrgZtNa/dpp3
+VjH8K0cME5+SXU8dR2xmj6WVwvWR/yxIGXbEmFLObrzM8tUtD8swQpD40rjcQXHkvagrrif8Pa9
6d8ARVUkGVWQWJrmhvc4WJHCZX79IG9vtVpHQ0UE8mLuo0QbNsLn0gcT6UE9Vl/VB6tRPk7cv4p4
ql/F09JGZ74sUM2Gp1xAV1XPotDEmFcbqrZIZxbFRRjtC10tW4YlxWDuM2XZ96dTacRFJLzcPqho
lf1ZlMdyHMe6Y09LOLJC9EGxoWCqZyq2Vd3gZRUSskh2r2/YU2UOBHThxcAajXzoFXB+iTi9zWjy
Bo61TXzd/o/R3bkel6jYNlUmKEsgNwnZu80LN8/GYaGEKbMDlpZ0IlaJVVHWsZHzI9kwhoAKd88T
Vw0R19Jw1LHdVaKs/OPLJ2UPmroWKiwcCTFoYXLeAiJ4tDvRCqfrZXkNdMRJ8iwOKbv8EwVyB7RQ
g0YsZ07uq7smtVxjL0OO4xvLQdig2WZWFKqJ3tjTCaMBGIjeEzzTQHj8Mp6DuHNBTlsHHBoy9/Q9
sxWDVcX7cfWAHEhMPJwUiihTkeBpY423PhVyQU09kvlyWjOJhrE52QdQ7JBu1PWEVNAJZmE0IuFy
dCI+EJcR3WT7MoCtKv7rPModFTOo38pybx7xgx9QoreYEOfhFCR7bfef/UxDLcKELHsvfNhScysh
hZogtBA1i4jNGyCwezM6Y/MURZb8rMRokeCzalGfCBeBluw1ox4VGfleRgmrtAKh4PzJ2+z5eq59
9dDCzWl6G1bljg8x17aYvJfZ8rOMHo5irQOyA8ZeouyTKw5yiYXv7VQNOGumEijwc7dNPaXVx1uM
zT7iXinqzBm5Fua7Sy+kpmqhxLNImdaiakuWi0y9i/3YlfQkPy71MZuMoxW77bQrYeWaLNZU+w5w
ot2/MlHo5rOP5rn8EXbNh54qFgROs1L37AsAmZ+nrp2BaJHfvx/PExwzcIIiYbiNo4OwaXYjYFaZ
0kFHA67zB+jro0pegW0ecSXky2e9ahKa5nPXjIQxWzSWibcuIKPaRl0ccdOI6opR9TBDPf7YaVSi
o2ubAS3yxHcjDsud85jQQTKj4fugNzzvDnaZ0GziJlVRZkmb37Q8PtAbnQEmA6ei402H3sQzdtdQ
w2GyFvfHIh9A8GPJ1L/4woXfcxVopNLFldYYLHggnVccy4AKfwF8xD2RfjCS8IyOFeIANWJxiiHI
H3xqsuMpXE4fkSjKSDPb7/jvbnR4CjxgC5IQDBnOqZ44Cc0nQuhDYrU7orMK2RlrtqlZv1+QuAln
JH6aI2IJKSpv0i6BvfcyTwsuCeW30pGn4inGeWiqKMJ6wUJaSkFNGPHljGXsquQMLOeeowRgOSxH
Qo3lGNDUzK3inY0eOTELTg4O3qTUphvjpUpRipwXcb18oOjN5a3ZSvuFaFtM3TIqPmYfbbNNXOVG
dqqwuaimCR6jeL/Ih9nxNuM3Cw+T18r+VcsXSGNOHW/xdor1CoWeOmXsjvtAt/XVQlgoFmlE6VWt
SUWa5quiavCkWPjQiv9guShqq1IB0Wla325++o8RZMjCkhmVUnDbn/WZ1WSD3I0+3VUPKTEWYMSd
2VJD4lbETc4Kpifga4h/dhJfrk9OCxX8jqImbFfXycK+1OwqSMqvbGR6LRqsCydCX4iVCUblhr7b
NG9Omww9Dtpf9FPeAu/Q7VriI1j35uzkTZ+wTT+T1ea/S6+TU6C97WxE75iii283qHhzuObPlgA9
b42QNTP4qr5D1lZxGN7/UrSiTioHyyD+UfU3TzhS2Li1xRlyN6D8/3eMCefWPMP/CdBue9lQi2o5
a2mI+uiNwVKXRf5T2I2Qm88YHCL1EFB68btpTVSCT8h1mSfMJvtp3UENrTZQbb+qaHaN6wjuDR4+
4cAXj1ZntjI2Wcx1xwx/PYbe/JzD3rg7mUI47BYD+G45xBgPVqI9B0qipGNVjQRSjHgnMhfGhz62
YP5kLXjwXHRNOITeQAfvLXwO/ZESfbgJvlAPwFWR3e+1Vrd5LIQQFXX6hU08a/9BxHf4qPPO0yxr
VH/Rp6BeLcJ00TJa7XcTbdB6qLXzGGPAjMRmzZfYkXRgeeLoUxdK33kWD7oFeNIuprgUT0j1pRfV
j//zDZOxJ4kcQ96KE6O0GCGPfTtDYuZ9amSvPbALsgLss55h8/WqOvJ0biYQeSg6Ea45fkTbTGWI
SzWX2jMJNCaDc3RoaTb4LzqCA7KsqraeeWQWtqoKvgp0uLiKXWVngjyK/jplX7hpjy8h2g2pT7pY
2zLexf2qtU6WOJZ/MTBwMqTYGj6YszH0O9zV9gtXjXochwHADhzHfMHWJEkNj/8tUhjYiZOtALoi
4dkaMlLB3iidxY0tPZML6rr4Py2b95EhyweGlY0Qp9S91TvdJLbCJ64PHyh0LYcCcjTLpZzcH42x
oAA2f2k2FM0YQcLFva7m0+RS9MsmeKzSJ/XF+HKOX2Zdhq5Yu6ToKIS2zlTVM0y3W64QllLBlU8m
BLcNj3e13SmTuRO14MRYV532gLXfainTDIv5jUFiS/ayUDk1DHXU26fO7B1PqT+fdjKEfnQK3VJe
vkRQHUldPiZ495djzmWXAnWtJXJ87uiAIt4GOMilwpGMFifh80gBDJzBUy4NzV9g1NRuR8JXgAj0
yWmDKzj5KGBTNFxfhTmEt+3rDlY+Tz9sA4cgH5CEESLeVyEkYvbspl4B4i0H8kG7MtlJWj5ubVQs
nE/lYu1oZnK5DmSk1AkEEIrEZN+7KDM6VcO/qM1Xis4h5Dp5OBtWiZ23fcfqr7VKIVWPqMyATPx6
0RgkxyHBzBLyHdtCruGuqcvS3iKLAWtEvHnADVWOYrtCUwNqcI3qR8JMhxTfRKwY/VYEd3MDMNO+
VNRyrjyaoL7NKIrT4zdica+oWMR9+2+m0Tz7uZAyZFwzQPve0j7jxzMfxRKrq1C5jAD8tSAL7ntm
sCBjtgLczoBsHzIJPjQocC2xK1FRo9d5wKJkwC/Z5qLlYE8QngTDcyuTJNFstisqTsIjfWQ3ytb8
Ne3BPm0R26syKP7/sdIlovrzo2h7D2ZNjPFEF6bXJCCld0UaTSo0lvb9vogOEPS1f9317sSkyCya
lfmkTmy9bPvGyFz9MmZTJAZg81DmGN97tNm7djM5f/+jmbvJRUwlRuWL5cQJq5BQ0JG1R7CrazuD
jvjXsZMLQLdjsytrh9U+tdVufB7M6PxXZTeoBse9eYCqThLTmGdUBrf+XAQf5BqcnVp849UWejYL
LcN8+ymzBwOXBVPRzmX+mE2Rf/bEpaZUr7PvM2M3xp9bcTTnEin3eBYpHFGSZs65aYOVMbMYa47d
J134N7AA9BDlgW+6AMmAGo4CmjjC3TGfME10R5BR1bP/CSNQCIyZZ0znjBqC8+6e5gMffqChBpA/
vzQWE0PpDlACcedOV2TOtLmiASUpuS9+ozgBDBIsu1UV9MiVtj/FV9xGbbqTm2Gc/saPEoIDpLab
td0iI+41PtHRRJWxUs1UrHsu8DLRgh0Ar/xDf9CT9Qe5T6asARTSVlXjg5rF8FiZhbvuBxzF17ES
RVA3oE5Ut3SSL8mTu5/hQGNgM3Y8i1OxxSvjB8ndQScyeXqU1s6RnJshcZSoMig15DA5tHuR9NsM
rFqY82KnGuf1OWVAtHVLlSuuG3edm5/CVb2b1G5fYbFTBjVUqvXnEqjjipu58u7U/g+g3bjyl0s1
4fGS1X5IbjbR1UvG75OtMC6vWCSxEEK3SPFSGu8Kexl/DS1Rk47J3+jeiT6jxVNcalU0BN75ycAX
xRqBp+xrtREgYXMwuEY5r1reHCo5BkZxjDAoCJ1wfQf9nQGZfT6dXK7ERf8X4nWBwbcwhGJ9A2WG
+FFf8RWy3/uvqSTBqrKU9Xqu+GG3GmFkOT52IxrTu/tsFk1d7ZFHXJgCpEVOhkDRuFLfMHaJ8TiK
QKWZVOgd9Q3YBWjuduCXB80+ENhpNpV4z5fJzL08BARLegJAOXTjPu6aDTVmuEWA9uWfYudK6Ktc
0GN2qoa5+rg48gWpRhpjWEkMwjAjzR801nTwFn0WLlV+pi0dLds54keaOKT/Bt7TM2c7UsHHZlhX
Wz5duOQ+XoPeU2knKcnvfVHDb8itDjb2cBD3FrRnJoKAKm+jvM5BtaOH3g9ijly4WyQSkfxYltST
ACDd7AQ/K4ZvCwtdqT+ahW7dCHtt+s8kgjbZE+oxQxr+RIDNwAJMyYY1ezwG7uiUM/SIXbGG/u37
ACOoJgYcQELMuhiJyEJ/TL45u58Oe2L2iXSUkmre2SLR5fwE7I92Rhxaip3x1SK4CBwQIxofCrFy
mE+ZEJvFSJBMp2mln0KngrjmC5RckBd8bqvXYm09zzJcfj/y7S0WxqX1VQv/elftxU/YN35KZFsN
3ZMYZLIN8KTFAXBcXio9lGt/2eo1EcFgJljiV2rb03yqC0p0dyWyCHZiSnGOUQdXhF4ESNDYIkDJ
eAAgo0NvYyxEK5UOoSZ5kU0Y+ALe9c6Q+dYLwMWksir/jc2EiiZ/5+LyzfHJ8UOSSsxZ25haMBGJ
HOCCTGKspn/8SiWrUHiTZf01vYMunObNULln1Hh7UEqDLsnRFOM6/aNaWyHZRfe4Y4i7iJwQjmso
nk8a+V93Ndi1zvINU8IV5zgXCnGap93HOdSpTjdinASTAasFqxtJ06EfVA1OsIagXDijxnDUQwQ6
uwbK/+RbwS9H/gT5gRq9I+csMdhIzNIj5Nr364x626+BUyH7fin6RzRB9X/sxtFbUHk2EmJwKb/f
85eESdV0HQ7p4g5ErE9JuX0XIeVXNI9RNkdhkHd99W7z9paXDdJGnzTK7t1Bk1iC8wrG6AVvnLUQ
vMerqgQ/SpCnbUzbC4G29zSf3L2gmwtRFc//+De1r6jYmbfMVotaoLgzGTI4x2QHv2s+Xnx5/hFB
tCGb30CW+hOxdZxwUDVSs2REZ1tg0VhYCMJkNHPuXVoZZUUnpWurV5DpWpoUWBJHG44jOatYR6d7
r99GtAB9dZq/GLUY/B7lM+7ctdOKJtA5JEJwtSGhvq9xvnkZMm1T8bhAiXbBglpJIZOr7cc8zrQ7
DrjpgJeEfoCyV0Pent5Yca+Hs++PfbkiDDObhE9HBY2V7sJ6mIRwooNh2Xlg+SRA3wyPkH1aoK9A
MIxA+86IOhv5Xw0YCNufwRn5f12MBk2NkFeRVj7C9Vrx/MkBDmmIi7p/R6QIVPLs61678eTGT+EW
grlK7CS2ugSEmPDtxoagFFBZWogDPAJYcfmM8Syrs+BcTC5BcT1LQ7yeNdhNNOOT+oQ7hSHYYc0E
80VQxDP5pl07J7C8k+fBL6SF4CHJVaIOMYq6L8OzOhAqptZ58t+zeP1XnC5NDx5Mds79HoThcaeR
oDREHk19TcKIF9VZHHuD3YQ6Mi73HjpEhErDtxUgx7qZhmeEhCCmHYUWiqiyShjCpDEFndeIgbHI
p6esl2dPSkiTlQRoAgkLR+CEllnrtpmw//SfSUUqezbJWHNrjatyqnT41OgudDqMocO0tjObe+EP
3JbP1p462c1+28Efm8cbkyb+tsV/LuZwztQSQnYJt6MuCRpG//hKFpvEQEtx3X6QgqIB708XlTmH
S6CWb/hcpdK1d+FZRwKrgelIOW5TJei/pfvgoVwG2VH1lQGwLMNPCxNKfHmYqpcZ/FjeHOl1HFbM
FVBosgMdq3be2ePUvajyphtPCy1a99Ic5LLR7lSptwkyogJLiaLjuGjNMJB5XGCv1ZAOz9eecA+C
b9kOH/50tO0G1H6YGJEuEb4Y5oTbodcLhPG2znwUq9f1c1L0nYu2o7mqWA/GH2QsLBNxmuNpxhTr
pQAariPCtLyXZh/o4+mYcKuRPyieRVYbEAyuhqzpbokulng9dwveXY0Y5SlhfpG4aMho4DSBTGZt
WeLNrwawcfYCgrJ8THBiStXbO1lAOKV72Ae2v190pKxb9fRJugTAO83TYOGbqodsctGGEoj74551
j8DN0YCr2o1YP4+gvm2iMmx7vYLyYfXzAE+01V4mg65mXaFlJ8pIU7zFNYIcFm6KpzsNxJRZlOlT
hyH5PMI/pboWF5taJP0OYPWqPPHimbcdBlanxHBsSS/a8kmZzh2TxD3QeEJt7ZgN/LIx3kqOjInP
EFU+Xt8nz7eZl5Lcnzg1zqgR/5UMEmeHws0g8oGa4Yu0J0+Hie9nH44RJ2H5HWbF5Q42G184o6oP
mrLWBjoUK4mB4jT27ckGLX6lrKuZPZUB9VdouVan9AK/0HA3no0ZiDgVrig804zC6K+gwZFA7RC+
RD7OVLmCyvCdCriMkSEYFmIfQbERApxGM2cvTVOjjW/CRAbtRwbwctLmiY83OYs8QiFqfwbz18b/
5xbeosl1DQd/W+S1krDAKTUxEfObj2UyzRFacn8ORHyNoy03CtJ/P5DlmrmMemLeXr69iCnZmQqu
wW+veIeA4C5W/3I3pYDxjOA9rFuLlxpXFY6C+dYjdY1uNfQaSKlGwBP+U9jwVNAHv4SZ37zg1iZt
v6DqhXSxKNcJRMFgr7tIBgfwaX157QGmyndr/c2VomWTMy0wSQLMy8u5E/lpKXd1JyjX8XAHBP3V
dPbi+v4Sc3WYc7UOgK2c4+8D6R6pLYFrKUWKyOR8pqOpHlSGPGBVRloPaoTiDa0ZGnXgl5b3dP1r
/vjutew96TsfWxo+5O72lYuMY8DTeAtXMBKyKAS2O1oclBJ9MOBS1ZQU5UUtyzPocr8e3dXOe2pl
EYEDDYSU3Z5hpo7M+kfZCWTypXhc6oNKO3ZqqZ2g8WoH1VF55g8VhpaYhd6tYXB+wZO3UMuY2WaK
xNhViDBaI9D1N5CAtMy2zxLQili2/VCDwd8lIr6UIAkhMia/XNCGS9iV75MK4SK+4w3I/huFp+HG
ZkHz3sLI62LvVPaX0YWggLoGCesgKXfCwegkFij2oUy36fRyF8hVPO84uLrKv+9KLb30Rj3p6oi8
oQY68BN9MG34YiHWmPHCGq2vkd7Z4TCUdRzEgTKL6RTzHfiMZ1tl2qvTWIbRSf8cR+k4FHAezr0s
wrkxQMzWLE80boIOOzDlvujI1eYtDHrqcAhA8tylmQJdyYm2QaHtaaYc2oPajErBxxGA2SF9zMmF
GnRqlreZMAYn01R7dI9EZt9uNK2TI6zvhNwF83J6KykLg9FM6qotRrXP1p3G/9yBJ/SHFBzLEJLN
NvNezDBbOmNcRUWLwE6Jp/esnyi2HFwiins8K7gZN/X9cNcDXkivYX4doUpgpQJMaFt/ZTkks2GI
h5yjHtOXv9XSUZ+OKAmpcR7NsymYW/LMOVhCEsxN0XjO3rr2rpvU6UrXABP2gGkOV2rmT24RUlnC
vEUyj9QyOVg4jFAXgxVLQP/ofJ+6Xc/6EVKCnGjW9ANJr5EUcGL8pDg5RQeYsoPOFmFfLYdjuVxb
cNIsurvHqLw2rKyYDNz5NGIcvGI/txtgEURG8XZLYZtaLitD99q5MsyAeY7P5MbKB6kYEtcQph1X
3GhsNOTicAtLqPf0DdqJ+6+mHPI8ge2m/Cw/rbdgaW1wFuquyXIAb/5Q7tWCREzF+2SIF6ayOqka
LmMsp8y3n4lshUyZoG1S5OzkoAUWpk8O7Bk8D6G04r8ByAY9gnTizRllUwdBNcfP625gCrfvS3bS
YQ/Zy7xVAv5t2ZZReLDgc+KfyNCErFFRYl3mw3yI0oOO7Hgn6UYC52b1zWEovB2f/3atrCmPgNAN
W0eQEziQFDX1J/rGJqvV8AJXwwB97EbwBaNCYha54B1PJFg9h9LeV1F29+JqEbtNQL1Dp7p0bDHT
e3iVhXmKXF0BA89Gx5kG/vwx5YqOobNqNY08GtkBhvwXpasgPPARlf7YjWLqCnj8wjGChP20LKuE
zqP8kbBMEs8Qeppb6j2nLQx17d4zgG+OZLPfEvpfi/+0HGThrxELv9SHQ1wm5A9tbd05K2bBU4cM
Pjs+ncIJKnhpsbLAazst890ANuAWNEIVXVCQlFDb3j+8iiPc4E0EeQ8rjLWFkDsjfSRLhiszBFsP
qjZLTWrntQ6A76rQmqYVMtbKhiguSjpTbTWnJoe/AY7KZIXcIz2+fHdnYIkb0jLmw/0Pkxzw19Yw
Q5XoNfxyxq38BMDYXqq0me0ASAPjlIA/XeLGBEobqotxCVh0tCcGPzHdFS1r2yFcR+Dpj1taC6oS
PykfTzYdAyuKq8PALJL1nKT1VpDMr0vTlnmu8ySNzEblOqbCYOQj+iewAn2lykrI72UbTklhDg4P
OEC8Wi5CBN8MYXg/y3yr478NeD67uDB06MQW8/sTHeV8l+vvt8giDcrULORiYxCjGwFPRir/44ia
I/4FRwzZHzrwmCzkgsuQveX9s/GECsDVe7IjOLiucxJprxquaDnYKy/nOE7hY9SR4bMD+RqrKjVi
1CIJ4o2B7Gp6fMJ3mAQopEImNBvfqWqIgrYyFJXILf302Lbrov4IcuxW/Lltz81zCrDZ6CHeN4Z2
BnZU59aHW3fzLHWt2f633dzYx8/0KBaNASbUhAHY4azRR9rVK4bNNOiJHCWXLF3m+Pp1toTeZ+SL
mNMaWVqQIecK3hMdZ6EXT+MMd+ec7ThHgfFiu/MwtJHUqPxqdU5N32ZfUq5xyqGHeTf9GoKmHOHp
V0cgrgCGsRlaAizFSD+XFvwYErvT3bXI4gqg17f/rgVAwJzXKxLkOSOrXGt9kAmMAFhUdwiI5w/9
p3FPEMr+C95eX+xeN6Ac1fvJ4kMPoSeCNTqSOQmOxGsS9cYTNFYAohrXoz+QqZtjHGE5AIjbp2qB
RoBjhJO+Hiyl3xl44HoK4M8suLVV8LinqCI1m9T5/8qCMJIO0R7Qq0tcMuLFb8QKUCXMAZNVpj3P
W9o83TZUtNaCnwcnS8TdrSOsSlNfQ3UI6anGufSnn/8wj+5ZhUfwMe/0bOvHG3M14U+8/X2G9Nhb
mkPAd36FhAvBxNq2+dSmbUfR1fhrY/VCQ1+TdI/51SM0LHkL/eo8NncBeZfZyCXBzwLXeyequJ0i
QYmI2xihm2A6yvcHKUGyoAhB9oRBGehSwMu3LEIcmJpNoz+J7tWfWG//VbKn0wDdFhL5t7OS0EOx
gNbU52LLRYJLdE6/GNS28DYStySWz/MrY4r5u4PPmW7nBBEujKItO+/vtdH1g0IP+Mfs38YIBS/1
6Vcd1LIUyLdh+kdtiK15hN6hXj1tX97OmgolUbrwyzFrZGTrzkeo6DCYY8zHsx/Svq1THhXgQmN3
rlF2XHDY4mezean1K4jwgrwHZiLbA7ihOCTJ3f6y6ZYSCreRilPHUL4SSD4SC8NMDMrFpAW/DEAk
gcKNIXC3T6kv6KE9eBghzhGsHWGOSWjPS7YzscO+3RD69zFgOBxmryh18HeHN0n2vprFMLV3MLVz
1LitCDhC2O7P92ei9R0g15R0jA9c/xV2RQe9kqT9mZmqyzOvOgeAwnsc+JA4EJsE9r5LRVHBSGj0
Gf8iOop8g31aXCWxP9sGo/+rAeQfSV3hjLBnvtemRUtdYT+R41AXUY+1D1MVttviWIh8U4TMaY49
YfPALtvhJWqk2Lb/1kC5WxrpvuQc3krKYwUUBKPrmXzrJxLDDwr4ADpeL53hqMKMui27QWivLvxq
oznJ4fzsFPvwFU682lTh5yO9508HBJmt0baAgaIv6X1RfH8KO2kPzSt5ncnM7Ucplk4SiSLepnRm
KQ4v7+VZfex1Aiz0xSv3SfFc5YTC3PCxqm4wEuzyOf++9wq2nAnKxno7l7nFlHZKJXtDNqI2tP9W
PF1vdUn9JeR1bOxEl2GLJaV4eZ74Y2WGjGAIgo+lHOFMVTyCZ/DcCI8Jk/PTTOTfc8qLxnRCqAPQ
5WQIukZGNZWMDMg6ICq3LOih/qIZ0FqCYrpp44LJ+O/1ybX7KbIM3benlk9zYyUebnizaX6aMbQM
glXW+8RPcAPSRs4a60GH+oJT+2Nrxf9aGCS5jqT+WTDfP8cKUSOZQKYC4QsBRZ8JnGORLhWQz5NJ
AJ4lq7Ui27PHUBDU0kJQ1NYn1Jmnblr+n13pFhj+LkX2803OFFs5/AQASNliv6i6VKZfTVVvCOGN
CacaN7N8QclYgjw0QgOusgdWNFU79GiPYWNU53qiUf0Q4bG1JtdF7GslA2C0DKGVyHfUBAU6E1Qb
9gcH+T4+4q2askiPidPauFEXrAE1LUc77d7HD5zeXjOa7976uwVJWobIq/HKCV3YbY3BoTovGx/Z
N+trKaQNdc6sWhUkvK244R+3FbgbA8onXKaPO9UHylQdD3qJ74x+14pUXIc9Eslb61tLoKOmxJ95
eNOOtpCv5RaK46UNT7rSUsP3ELBqBxWPVzndxe2adgJrdAkHpInQk1YRhE+y5LikIo+JftbpTSK3
+G/pBIGD/bwhYwPCyAPhkjcL8+DyJvrdQtXkadFuMLI87D+RLucoDwQyxNx20+M0OZsbhb1iHOOF
Jct9uYU9ecnu9Fodpgs+vzLu7svWc+j1Dp64SRmFBQfBt4QTKZMAgfPdl4Pa7Ikzxyslb4mMX8iK
hIxNexP6YJCkF1Jgz6edMmG7ZTATQu+5V6X6QHTbL0N4c2fyrf7TCthIXVlTFYSMnge7GHa2+DBS
gcq1w/ylg9KPHopRh7JFey9e4dpRv+eYTlpn+NItT0VGkRfrDRz8A2oSuUPgsI57/fkcGNVGCU4e
NOPycjYJpzRLLIBTPiX0QsiydNx8auuBp2BeMMjEuvxx++KjJpdTyvV4BMG8ml0Uq7I1CWHdr0OZ
yvOxJhYhpwchlOwZ8W2TFMPkqMtgLvYKGtznkAHIFedhd3NXeLSTTcfQ5eboXK0P5DKvMHdpXp71
JkGisinuDCM0AFvKTEaFjJs/Ya3grXGhAVu7myZiKU1IitGIqdWMw4r3pKFyvaDrMlpI4HzSCNwn
0l6EvA1i92cvLm/MawRvZNEN92gl/4dqotGeJefKOZzXWkaJbo9d/59yKckIbiJYD062y31Mkga0
M9lTL97Wq0uG0+ap7P1Dz+zmtL0KeqhiGS12qqKOeseK+DwI8KsrONZ9cUgS3LHPqJ/K05p+cVBO
TKSnnWDISkmX3RxJIX+tRNXuq+ifFtrCeBp5PVWgbtVbaKG53fXYqsdALZunV/kM5hb5tTdB2nzv
AT9HZ1w1zwkHbv/lgCW2mKuAfyyIbDue2jGQXO17KLVZHR2mu6ecbK3fiFPT2GVAcXzsw6D0kYcO
Uc5isYxfY73qsOL7Fx373TDPJNuhH4B+lNwzaxnJr2cPVbHiCCQ7pDqvuAUot7nh38Ke2JdySbE0
dLpfahHNaByNooe7kOgviYoj3K4bya658MAdma9rM88j7O41m1dG4/9iyMz9shCVZcmO5bLb3o3l
6YccsbTwGzZ9TpyhWu8Q4UvIDGWGr3KNSq2bz6sru31XQ/6TSYLccoD7Je99LKwaSs9p2p8A2Go8
pjqDk0f5uUnWBWTX4/W59zmxDNxjuztK1uhDRfIEAWoK+CRpkZkO3ldowSFS+quJ5UDmYONyohZe
PFlJymiUweLYYWe/W3iNmb2fNcxkqEfKgQoUEUwmO6wwHqRfO4hz5UsFxFDBZqc5YwbEtruU3zmp
OsRD5fzQo7MbmCxqPHaaIBln4P/HfE2u2rW5a+See5OrflF62WmEnXPfiF022Wo8YufsZPP2vkRA
VXVpT0ioQhvFpGYVbWSbaCoN70rWJ6rNF1PYk4FEUW0tP/SsaO8Ei/x3CGTepKXfT8o036PMzWWD
9amp9/KhywKu9Vil9ZmiYIQWG6/W6/9ILekvv3XZjsFRQui428kr3074zd2q+q+gBs5frcAgm2O+
xrh6MUY1+c5jqnbm1du7r87g4CtFCqGbZY0f3OPB6vOKnzXkuvPEQquy1q0rgGc9RTWsKbwoSLcz
9IvH+IOSs9SeMTAxgnxiLzXMthkjnvdVJtH8rrS3tbhmxwdkiDP+O/nc6na7MvzUizJZcHxQRe9A
dWDuq5MYTZ0L0rpdnJfXsJNCdGpQmKBJ7S8XBKsFYs7qPDCXDBDNebBD1K0SNS0nHZyPN9+Djlil
64Ql0yJDxWAqsMuFF3/S7gZhzrNzjj7wuSjkya4HDuc7MEYIXUjodS/So8A7GPMtpUA6Oh2V1Lto
jqGtg2LF4yqEyInp4NPHWmWMVpudIVuhi9GDyv3yQ586SYBODMM9r+HjkxZRw+Vw87k0+tOxIRJj
dLhVhw3+grsz+t1abwJaKXH9mF69oqFynvO8Cxml9WnwPDWokOvnuuUQpAvNEQgsdl5xbMw58EIU
PZjRKKlhrfaf599Vnuu7j0OCpcLdg5r5+UbxtDYhtOuo8sZLAg3h8HsiL0Y7O5bAOfIt8FTgUIpG
Jl2Zom091IlujDBQgHYykaa/UqxIPIATd9DfwyLglDSa5ZbfP2xcvrEXe8BejvWpEVmCWXmW4rvI
HiYhifZkPp8TYpPr8fpXjJu+VmkYsRsss3ldOWy7gPlwm8jXMAEqlwhcWWUQgRGTMHpDB59dVhCL
zC+/UXqv2iD4CWJH7SMv0S1NDZz8zyMBD6Y2bDSI9RM2FchWP+YIs+aan9IOTlhAbPYR6JKjoMYj
HqGaTDtbF6RVI2/8gfgdEo776euzF2NpVNOly8LAWJnAhhG9Qkex4x0byv+xkicfSBpSA946Msdn
PVdd5mfHxw7EZVP4QfFQVQ9SS5wf51LVtaQalv1scKTWmOZ7QnEIcFz+tUZ9dcOAwu2dzSPpQUVu
PVzIXoXL6FKjX3A+HtZZtaauUA+hBxOt+gblH77YITonj0dRqxnlAO96HVNXlMfnhyv/j3Wsohb6
OEf1tLV6KKkXmgNAd4Uy4qBoNqQ4PwPI7wYY9qoYFybmifclzpQRdF5r+3U8uIbQw+jFvCGB1glF
2c3i+lZm95Q3kHyGEUKhTk3YmQb4ygOu4cCtq8iedpOHB4WnjpGr8G/zhH5JZq4cV94Mu9B4TxFl
hJD1/uGm8K4uEIzXgL5N6pO54sl2Fu9iY+aencr6C2+AASTl7vF46aWp05S2WFLsG6Cu0AxU4ADa
23pDYknyxtxNnJ5vlUr4AzxGPdP653KH3LDqYlCC6ukFzj77ezEszdaI/x4ol27qBIxHt5s3m8W1
3v+DPauZJt8syjVtQt9KMZCgF3Bi+Es9YCd5FwC3z6z4gKsr5pa9fln1r1TMJBkSIKmloAx1rzWj
D5X7AeOMVY6nlU2uIOeTCwqr9yktskAS0azIJaKFW32w0AfFNOPch1cmRYeNAbyKkHzPwUQGYwXI
IuxLu7uArlBzPCbiVjvCh7JlNeBPDzja+Vi1MboVsUHbczyVCCt8zobs8GMF/4y8gGsWfx1aSKlP
BMSmO8xjG3Ue48Qv4mMUxfdLlj6m/jLIluQBB5KqAgNloDttLfA7BxtpEtK8x2vgi7WYzrZG6AvR
+maS6sCDouWcQsWpJgR6j67+9Td1xxLp52JLG96t/mQ5yi52qhYOPycyJNyJMRwTVxxkQPuy+b8F
bwWANVWanuX6tzoh47CiwqKKAOdXhwZNDrkkwGq7T+27Eq5byDg94dk4rVFM5AdkmLaTaQgtx4zW
+fHI06A2zK30pWIKndADWQvE+argCYYnCj4RwQ0Sb07UpkRw7WjGJ59h3gUdltVkiJ5ZxpamtjBH
0ykqBGCpZHV/Zre6WaK50FQExog7paYK4nVvTh3czSXfvhZDhAjvdQ+Otfz8Z7N/p+bard/ybE1K
7Pk4DKsbCLYrf2bVGCHsHumexTci27zPyJtJvk6IWy5hhMhit+b7ZEniAV6F2C47buOQKqh/KZCZ
Cplk5zRvv3y4QsKbKt+QEEAjK0FoxE4tFwLQTo9JCvKynEsCWG8mwN/fO/UzBt20gC9XkZty1yn0
lSb4VvNvJPVqrDP7qL5ad3I6lO3koC2Y+SBr3Akj26p0RFo36aECv8zXAJF84DKB2AQhON5zJFIf
6eo79CrVikPXoq9Jdpm6lYNQQm6hq8i4PlwHbptFKfTKvVu35GWWZnnLApaJhHso6jq9qzcvNUEP
QJgiTuw+sJpCA9KWWgI6t0zMLNe0gf/jvQp9r6IFlQCnekNi8Xy8kkELtj7qPel+faG/tS8cC/w2
gIwdC544bh5mwaIAuQr0lhKK8qE6cc02TYrgPBoCTeSeT5KB8HE63mdMFIPKAxKVrA2EPsTnDk66
YjiRdQpZxw0broCsgvwAtNaot/s5c790GW0reJv/Esl71lLLK70VuF8JV/622KoNOjsoKUUCbSg+
DrrUF8amuUw0g1tGE82sjGihmSqu6OZOu5Pjcpjc5VJCVWyZ/JGlLxy/8SEvoD7F1U0i/IiSzJwS
W6XaQ4O2IUzxoKZmEypQnCg8FhDqGlJIf3JEuDxLiT0+cVVoozeeoK5BPEEJZxNjk4f6jkYy1qAr
AqBoHBxcL68e7X+AzqggjO+CYkMpP6jTYzUWBs2D5dKFBYwGhaO63MsWj4KVEl3mCRgD6d7ViiyR
BQ6ziqeESb8pnkfJvxgRSkBLMmX410FqevPyxUDrF6HCTGZJocT+IBRWbniZk6O+Z6cJM5zsOwU8
lQ7w2l9Xd5vcOLxJ9WQtv2pgoJI2ZwbmPYf314W32QmuApexFCxMG5bXALSuM/H1tvX7vucGiEhW
zHR113P0BlibiK23RMR0dHcqnOL2OtXXOga8G1S27UtDzh4uQ5nC5sd1+Roexfg4jW/1W7SJ4yuc
RXbkyMOjFUkxjRm6pSHF1XdrnnY89SkHLWSskhWduD73Cvy+8lGumqYPr20DttKY4ypPQyRiwyNY
xJGXivdIoUlWtSS9rJFo5+gSyzwCkATLBk/a68ih+Xv1XU9nx/BfCc9mupQa2m2oTquWB8G+1hEN
KB0wqYG3XIyTfu691fq5tMqgyiaTLr8Pqpf82oaSNOJrrZqAi3o7zf1XStxiz1M4SZyKIix2uKHP
8QZohJ5jN+nf8DFN6uxIQK03AK+7UzgFnuke4Md/eoBjTfv+O5pQ/RwG0uiRjtaXd0eROt8hSyZr
0Fox2D7NJwWNIYudp2th6XmL1w60EBZ/NxUKWjymtQLb6kPYkUNCHDc1vHIzJey7rd4CuGP3jUem
mX0aJvgBaoGB2Xa989EJ6kq2JrHBSqKllyRl+IaXKIlOx5a2X3Zn94LHhx0jdGCygxS3K5PRnIJP
+zfDMpWZNz1MVGR3suNuJnxJ8tZQi6Kke9DPjwJp/n8iKr95UD2g3+o2yggx3hlxFdZ6aP16Dy3K
3D38IqH6Qitzn4VfTdj2MtiJcbKLI6OdrmRC87gvo+S4B1X28KmC5QXi8rdwO4tK+pwwp/Wnv2nJ
HS1o+xseGr1jL+vPpQWoUMZ6IFXnzez26ADp9w/kBWhuFIfPt2EXEvvH+ABzBuQkpqyQgwRqlTsq
vXSppbQMYq1vRqpjN1BqFaIVr3FFhU8Gmcu85R0lLyYoiAZOI+qqTgb8mTlu+Ick6U09IkJFpwJo
JiLpHyYZepZmNd0n+15T5XbsRHkEe1RFL9MXZ5FPHjiS/Ye6Pyei+/aQVm4eT5A0HfMbK71TzS8f
J4CXtW7P7b+rh2DCwdypXVLyvCGp9g7moHF0C49fCY0ge4vs1DgIH6JiACybS1d4YgDyEczp7n9s
JmXVMZ4GbqgkaWU6VKdCYMtn7p5BqLYIifgGEu5wALqhJv3owPTgFn9/urM+vIdgvxIEO+gUuWBu
ejquM9yAZy0hQ+yWhKSp3yauA/tJ7WyxVODawbBigjXf17Ifl+c5vVLOonjwDJzmoR5nLvNSHdmj
j490bWinKNThD/Qu3GZjkwJEWrqBNul+fw48UURY9sH33tSA29khOusesP1bjOjbxNMh4K9u9Agy
hEfoePn3Goi60C92OvBa/vbhAytFer14jlAfSN5geF8+dPjI2vMght3yZrE/+2CGVaRYnQ/9m2Aj
/Yu5+8v63rsfa+vtD9va7H7ZX19kh3yZbwBJVkIE3KuIFsX+yxdCXCnewLQTLY3ObmlvrQozoOhi
B1HU6pnB71Z9jBT5WrRBqELWA1fe57ZmT0G4sUsTs96PdEoVfhFmJ7D1MPk+AJHQw8ei2CG/VAzl
gLgHtk8qYMonsOeHaWQvcDwUFkJ7KAaAaaEz2FKzyQtwiZd8iJdud1VGvV2eMNwPqwjLJt8jvzmR
oNTnq9LU3xQVDHseuzlTTfFAIotLPLHmpk6Eff6KLT735Py6i9zjzxu0wQesYgNhAcj42y0FbmJL
Npd91W5XYB+4NBq3/fBssuubLlVBhv3ZzRWiq3QtjJSzvw2nFnic9SxjvYg+2H5daQ3+X+eyfbJA
pVma8Wbdva2QXqYscuh09UpUV67A5OixBZYQoCE/GlZ94AVcfybc1KQ2uP113DudANw/e3FqBMg5
HhOLGM4UvSAtD4Vqog6AdqWMrlxgv/Ebj3pCnbA9yqxYKTh0Qw0ihLtt3vpo+sn/Vlb7xrsd6a7Z
vQvojtCybVo1d4rqWqVAcuTnUb28VPxfSxs6SkT92Xix151Uj6+aYE6nk8o34NUE/sSvqaKL92B2
g516UNpNBSSGz3cDpMFVlX7LOQzFUW1YYp2l6+WHJb4sogkD61YrA3xcviBOwEjTPlgn5YjfvANz
DfPpkBLiBj8L0l/qZXBsx6rD33vrdw6jpRt3Z6iaYdN/r3UvNLmVgq2t5XtBYTgQc9cVwaF1uLli
iL01wnAkxb+jxQNNjZ2Plg6Kug3zp06H7slPn0+IFthdgLE6u/U19p4hQpDEYfubXXJb7p1zu7Uw
UyNtAoYzQWs7QdyrC+3M8xsRZb3IIj0sRopN48HCYdI4kXdYm9RUER2o+q1fPX8Zh+Z4xyuuGIuz
Mrw5zoLZUzhUnLOWo2wKHjldAN9r0kqrSoDCX4ICNSEWJkxYNpEfS1WJppy/COQqtb3m9vIzmc/i
78JDWhm1FAdDz4pAymth5WRdd8J7Gl09XEn7CyiI3fwDxTAKN/YVuPQyX7yBeVsl7sE7c/8SuQwo
tjgkVl1m9V/BoZ0wuFc/oAjFK+LVhKEtjZo58zquc44ICvz1Gy/qauZsZyNuXw7p7LLgF4MahyQT
FBJpgXLyrpHpxvV3I7oXzJUapAlzBRqXFaqHAhQ/G96P1oEivAirD6HW3jWVTvGOkrdcizgfLJf+
iAE53YhtfImoL9MfrGE456UAUomlV8dflzsP2I1Wb0BePX5DqewzmqL9aQ9Dts0zT6z/I3H/Rzq9
ILGhlOYv7EVxI64VD3+LxnWpOP2vyQk+0Md74JIBhgFf+sGce31lTbwME+RofN1Cf3WQlVMBcq6x
X4BoMvexKSlRIKSz8+1yc9yyfMiOT1MUH2UTEmz5v4y9LVMsr50MliABfFF76W8mN/X+xF0+adaI
yyG+3POD9E4v0N4HRhqDlZg5stpZqQOvfkQiJdB34SnolIFAF0pmrJzXD5XX0E3zPXjAEkewzCsZ
evy/Z85zlwkGhem8lQsbonp3HgRKIrI6qzW0QHdGVUEbxjc63quqcLAMKsDCTBjD5mUePwlym5WX
QWrDHHtl7lB9K8GeUOT48qHpTHxzb3gyHqGBagHYzJVY/HFALm05ozghXXCDrkPN4Cya3C4pQEsB
3Fz4GW+SD91CVWBVhaSJG816Qgr0dSnQaxsC6i9mBuhhpkpKbk2+fpWfL3mHfTrqgWE0VfxjJyOX
83trPTeB3+XQAW/1AmT93Pq8ESgwqopn44OvL+Pbeo2D+zCdvR8Ty1Qx08urAAGjUj/g/jKAH1u1
Nr22vOI9K3LZjIK8LqH5sZu7bxfX9W9UUfaxwagSTP44W4LzkAtOOvEK/enopTNAmXar44Q+WNge
J5Bn0OKNiSvnhb6SokW+FEXMKMrSA6Jn/pFYnP5vSg9csp6cA094lLpZIIJSx0r2HE5ioxUzL74p
Q07aUat/k9kP8wpOKBqyxiUwwTSD0f0dsbY3n5FG2G3eGrthS1kp5KDJvWgDMux6YL+n7qzMhoR/
nCluGjeVFZ3oBL1JaNQkBCCgBx/kZ/AE5LAPq7QwEp2n2BqxXtzE4A/GVbZlkTaexqthwyvJIYTj
+usc/ltIhGc/2eTLMWgkLVXwrZbWBCXEMPQ72VmelcxSACgfgP8wyI71cBxGdRvpR0snly/jzpIn
hLIZz5f8jTSV90rjlPtX/MuG6Z8GX12xVdrUHXae38s0v597dkE4Nbjfw08DvCD9sXXoPtQDWfa9
bX6dvjKl0sFDHytfrXVK2/9IDxKq9aqYr7SxehEHomi022v+4Q6utLT0a58HMrDZUXOO7HEqIJzO
8t1PGyduTvakfDZJoiHJ+G4lF4c5dQ10XvoH+chlV0lf6oyLDpyKN079zHS1b6/jOftio8CKLUd0
KBPYAWllSlv6aJH5qjkQ5wT56UaerSDGafFDYA+j7ijGR4TrQZkyKldBCx7gaQiJY/euNjTbJXCk
z+lSixdoMPYtEWANmAXXxskIERhrY4D0nhjsweG0nt57R5JWeY+ajWv3EfBrXPPCLIK7YT5/islE
pwpgLjmcfKXB+chYaSecocLzFd1GsZtinm622ENY+dSVQdJSEMON3zp9+PRVGnCheTI8c5WcmMJA
fomiRESUOyexdjxGBDCUV03crv0Tg4MnBCXcNBRxSC2mdVaM+Uw5hm/pj29/VQILWL+V1nFIkZ20
7cxMk4XfX3GdOhYqeGzOM/IJ5qQjXxkNNoAflrNcEgcZVeyAJ8zX9ArmaGrr/bZ75X15IEYwhlef
mcIL9Jfki8qVEMNYY1iYt7DZTDC7jqeJD9kOLvV6JS3w2F4sq6WfyggjzJ1ufDYTesQSC/3VDsJc
M0w+47pJx0JTHWtNRdy93OWSFxEwZDj4KKGiTdPkZsie40SKCSEyOOnBIsPGVC7fnNCBHNSA0qZM
porQiqsXLZN2JFVmwQ35CK+n7/1vdYMCtnXVKuwin32Wm2A/TX6u05LscMLfYaPCTSstB8uBQUED
ynRXpJvxDH973j1Dbgeqdncax6WCc/uaZ9W1aioFxYS+dLIMarkMweur9jT0beWkh2qrUt9/07e2
yVa1cD9ANAFXzbziGhl/i5dWthHzV86Jm9q932VuZL1pe/7nkvIC4oMmt8CfcUwJGA6PzhGEdSmg
iMKPMOYMgUJJbGLQBRQdLpDU3cnzzO/qlafL5QExxJLYwPz0ITpKbZShNHPqOZQF3yrnHJbi7ywy
SQF4VbKfpfGEcjo5TX/ef1jcrYOTAffEwZMT9EAxzQBf5NOVHQYpp6Fn1AhNQMf4EwZJtLKRyfjt
1KVv3goJsxKccQfWDExhNl2BnZfcSiSpbFyxZUJYyQrTAUgP72/Ra0DbH7Y/LRon4F4KRm4Qia4z
s5/u8NgU7ORZt0Mh4aZ36tKRF0+7gbe4FO9SWjNBFfIsfanVKFTdZ+r+uyOR+PcE6fcaN5lPezMj
HI9almeU+tRdf+yb+tCj7+1IhJloontW2TfY5Q1rN9ZMoHDLDdDMI3EUJyX9CrOAxxoyUnu3BmpM
+VIkvGByyjpCY2HNcTtnBndlvJ+0gKK3Q0Uvj5/X+deI551QlhGCw9IdqK7N0W9mJV/aYutuJPFo
G+alT6ON2vbnZB6Lh/pzisgHxd3QonzJSDm6e88HLl+nsbufV9M4h8DNFoBW4DwPVsKVCPKZ+vk/
DlbjqAVHAuYhGFcX3OoVjThQ/L4Exvf4iwThlHFAovLscdBFqzSx0de+g6ujML53ZOGaHKG0R2kn
+dYNh0sek8789XhMDI+1x/mGAyzsFH6Y+gvMoO41cXXDKQ8gRaW/jRQNCBzRT43xefjM56FwkT+r
Sq/eykl4HekEEZkG/ZNNpSb5Ichbm/+YPgHa3iwR9BgtSfIYbSw/ImE5BTIO1t/8NtaBNyiThOe4
XlhSssAqSqF822SwsRKl99RCiqfak9hXdKkn1S3WvA72nE8P1n9iv1dkto5SEyLeJCQaEY1i5Ms4
YePfsT4LZzZRgTWdrSZ78WsIgCoLH0EtruxCXTvJhS8W9GZztL2d9nwaF47hFrYb+IyNRN8whopH
LlmT0vBJk7qbqcnS2HY/ERLobsTnWKfm5GhtYGdR4bXTSZkhX07O3r7W53l+sm2YjYzvBJ30rJuR
vkeHPAGs/5FSrxUxWLWwT+Cn/w7NUKcMd3Yfx/bORkTDv4CiyzhKdWinwVg/4Jm0t6Z8BZuZ/ujD
+EJWqTcbHwY876aNVVOmVxSIxSNyULBRTe9P8lDqQvxRKbxTpBRu5AJtrCWEnXFrEki34tvUiPGF
d7zK8UAsFpC1HbIuwrwlFqnWpH2pkx9fULNJjBJPtFgsn3oyu5h64MLJKIDKgKnKVZOe09uJLaRH
WlPWAYsWm/xxQfz33j0Gu8Qmg/wpsy3+pKef5VyEAKJl7S6qxb2sDWUmqZkzaMlQwuIgY/iPDbmn
LgCIoEqHienKMj1eJXKjo9rh1RmgW8EsncBPenZxh85xfkpq2+Mwq+XoJ/Qubi/l6xpa9R6bSjrE
OYczrdr/66l9HOYj56voeZcKBItRwnOcL2wkxyYbymlkBbn4gsEMm8jVjHnudmTpe/+conzfyguk
/AvXmb28qmf9lWA+cS/bsCq8v8Q46Sy36A7QifLjp57rlvdI2cMUptHX4WQ6owQyY0BaLSirFc12
s8148t/I6RCK10CUipsyfunpMHVQM/nfAreZWnSPfnzhbUWAmT3nREqHDfpKE98ngZYWyYhuZAiX
oMN+9CxfCJ0DBmoqObJ3Q9/HdecIc1mUhs6IoY4uhE1JoNaaexkPgDNrIicvVqvc+aGDIE92pd6H
e1BcEdN5l4RQgN0s5LOUm2g3zkUArTa1wXw0b+7yCbfuQX7NvHwLqJM++tB8IGR+aN26F7abr/wR
9ZKcEwvRbrBYyoTkJsBZhPTU/tAq61xA7FrlA2hXE4DRigpuXuwKlMvhFeNntMqE7ZmWGkFSDofw
hOnrNZghZ4JvxjT5WCFM2vlfFAe0EdTaI++OJPuruHpXErmHBGvHNRxAYdbU8bjzvDm9vRE4XhLd
iqt+0hEt5u3jkYJYvsbQDFFmVYcxnm8t1oroxPE57zhKyiNv72/H9ENl+0MiJC6VZbs2bHa3sEDR
Xgd9JrOkcOuF1AjKdjpRDVU4NxChY+T1xt+1AYYg6o0bWDX7pTxZ9ISNtCDAPWb/i5a2Z7+tfyQc
/mnlv6kzfSqzPkqSmfHXnDirP6VM9F2oAPIAp3gX+qUgGvcgBOjQukzDoRYr/kdrYQV9d1n7B1Bu
6ORS9Ouz+uQAriDy0Fsbe07ptxmjwalRvStR7+l1jIAhha0LXYpxRlJSianbZYeFtucTWcGYASie
s/oK5g/kZzlWXb4te/STzrs1gXmQf0E/tmJB2bSHVqpm9IEt4MPT3PJcaU5D8X0C0zNfez6z59Di
ufc3JpLn3yVg8FPJlDuCatLpLPExp3sjT3NIgFKRkVQFh+B4d6AhR4VCWa9iOLQHdjEnY1SpDlsw
DAjMGx8GsMwy8xDOPDWAT6U4t7sBLFDSDTxBXjMAZ5DP8cYmUyBGB5X8vjNv9MpqP4iiHjAjF8Pc
leX97ujL3liWYSgorM7dyq5H+jKT1R7h3PI/kDIAfhjgzb2sRgYHs9JP6OQImzGjHKEQMvf0Q3fV
9Oo/W2BC262OLUhw3A3cC3pruc0fH+MJzy4oQlqQ23mWsTVzV8Clya6ChGtOA0HmZSor0qPkitr6
CdQjsuSOwv0DGhocIqBM8enz2sVV7zf2MJJ5X5R5iRWtTdjTwdQk37usIlQVl+412YFWmkkUZxaf
pdPxrvaQlFtWQ0fAFbxs6YHAQ47bEziXYbxPxh8gEhxWkRaaSIh+hSvl4V0pSm4lVsurs1XyZJZb
6342l/u9LVmS9VnBs18g8U56zOkK7Ol8KTHBQNhk0a5aGqqZxCTQjj/bxw9jqA1oGU+1kZ+IMjwi
2OaCmSORkQPxS6MieBNU5JeUzw5cUw0fBvXicsfjnfTiKHS3DPwQ4yIo4fzAK63/WRmXd8VkzQhv
+8xFrqTNwGxG207SHKmox+vaHPf1B47Lsoo56p2fcEDjMz/5utCBjFVuK67yXu2Fa5tpgfW83a/5
/g0OSNu3IwC38NqOEBOfsSg09x5kMHLMj5fh8gSg2l9hIVzDPYhLHL9ODFS/UQVwdlO6VhcAuA44
Vch4JfVMY/ZAiAlo4Pam3izGg5qUtfrdzHPhp9LUapPjGnKlX/8cEUetf+DWWaFAF83v/v0HXzvf
tL4vdgLXg+8DcbpsFyikN1TfenCz3MwHMJmsAhqjF3YHs+xTi8SvgewQdiYdAkZu/Rj7KjMDid4c
XTZhNUlQZCOY/vTs0YBFQLY/QZxOgG4RzsSBg2WCH1Vd/ft3Teby3DuzxxQkVYwvWiYllVd6rLo+
2h9HNnMyy2KDjs+Z/gKUexxfHvd3UNpW4kIAZ60XCxDF6emt5CLyDNr195qBHNUHiCPP1LyBr8G7
I8gypY59eu3VcbbkczfgnvLG1IsLjC3679HXr5QSuViNpzqOc+w4i6lLUtsIm5ao2M/Yr31q7BRa
kxT7XYbfmTdBBBR90ItNzIEsg3FNKD2MVyro/ArhEFBOUi8Ff7MrMgRVtu6RseXsuvpXwP9YtpqB
zCM+36eLZ+tzzpb8RNUdXdPqzVnGZeatHR8lpTkIdkiFYmNz8rj9N5P7sxdz/slPjyVeQAxPr+uW
yRWBjfAI92RiYMA0LZZtKYAIfQyUouNcH/mg5ICeXenoP+WgHVngde4FnIj9TApgmpd9XUvMPAda
TqA3UMqLNujsSFUXqJZALMe3Zu24svSJRu/18l2Pw/66RFPUSMkyzOmoG+FSqOLSJJcatKzO3fYp
/k8BZ0UWDtru66SP9VJLSzEJEa0MxpsBy/wTiC/rGR7enK8jEan7YvFKd9kcCNoDFdoCjA5TxOoh
kh3v42R7ZjItKYqP5UyGDvYgraUQf88bjJi+HKQdr3yzUo45hrePilMK1qgyF59vebyvZhrBtR3j
KoHXHLD+3fxccDZldLEe5wGa38j0ne4CkqWD31oEMP5UDuED2G0EeEyhkWQzCSXJGr9a+bwRKqVp
bBVFPJI7HnCsOmhKLk2z/AQujdoh8rQG5LUuKZPfGT/QiC3z+wxk3lRVmfS7cFTIlszYzt9hzXxm
xQD6zJcv5jXjE8qEfYIqqbVFJ/b6wHWcUj16NaIaKpPCfY+3JRSmdNdSHGY6GRYTRBWyWB/0M2nd
43uPr3YaCbPYRyToxuoYt8nL7bO3xZGNsVcrBshRqjSYGOhJMy0gDAxUfXQpnVqUVHEdBNwzlrKy
VvHkGi5IdNkCyk91HoC0m8ITkjwM8OcXsjIlrRJjX3AXguUACA+86x2HHsLnLPy4mAfC28C+fUT3
YkFifx3Rv6R08Wq18I9nYSk6UXsr51aLpPTvMsBs8GBdQlO34EDwyILcUGsaCUvTY/lj4hTSdXgU
4rZ2+Kw36Wmo5s12LazHFodQmZMq6XgB5HtQw3zzNaAmb0ExjSeUtaPLR33sXIsPGvqdopQrCaSE
qb5f5QRklCZDgkX0nZOjEtIjKKg628Ud33xdxiu58U5R2epEqeLFuDyq1gh6FTsAJo7k/2B9Rs0Q
1S1pOdM/fawxzF24OhLGX1fba84zDxUTjM45X9WZW6QSP8/dBuCi0WChe5qK2fPKoyCr8aEiY8rG
wsxs4aNeT3fl9VyZO8RnxSmCZdLnJKQj2h8cX9Xx/IGeChK2quh/66jGLRbMfVtnVjLWJ5eUgh66
xAYSgJ6Gl8W+iiCJxfMMvv7r7hjn417N7fXbaiZ+W0GhRSwbqCQq+xhgc+AxAymAiaf1MuOX2Hul
kcIau9hseb41mcME9IrmFu61woGxmYbJFh/MO+fDB3VNlXELPHx63pxEQMCmUibYDgaB5mj5obY4
NpM5+Qfnf0Z8Qj15baSnLSO7DTqYa6uI46gnzE6m6cWTQGL87jwOFbIwaTPNfHFn2zDsS6m0qH83
OyMMYpf2Hs7jqFFDm62vSfLjH8rGPaWGe82594Iz3o59Yd4FPBc4vpVo49wbj1tzmm33HLjayKfN
CUbpD/lWI3EKCl4/RdyefVwwB1Cme4pPgAfn/dG3gLDFyhZWM8YNjGuAt5m8jcJSEyHhuqDDrXs7
DmAqO5uFMgJvLnV1FA+U1colVuqlGip822l9+Y6ZKnENr4kiihljQ4QZCBA8KsEmOsD3R/5OhVFh
4Fkf6VItzapcPVqjc9uZ1q5ZgjpCEc7HhsY8t7yOAR5tHxK5tRXPm/R/cCWKSctzMJLI5uWkqt4t
e5k5z4m8zRPLcy81gV/FmQx2hSSlFmbeakUMbEbCX9pN6Z8zUci/3LWOvZ4o1Ps+x6MJa+ePmtup
ZY2j6QuilDet4st4MsgL1rs+YkbPtP+UAIhun+oNndIkQcp4O3Z20+GWVCo+RdByEhXFBS0cw8FQ
TJhEpYwEbPBE2XT0/goUj9PfsnSiBzT6BUSeJRVLMtSaa58tSyUriDfYPZ62gTsY665VfsepJ5Y+
thrsqjkFAPEpD5pEcXGDSjjiBVqfl8VUndbnluKc7+pxrdapHghNoknZZReA980DKasGXNC/+rp+
AhVRhMLjX0Sj0sX3Kkj9bEoHpEdmGJJw80wFOWaggSgyrYU+9uW7EJwiPiCkWwyFfDEpBkXLEwz8
dXUh0bDYaQ5AY2QwP/mhaOgbjdEyNoO0bz/JeELoEGDvLlKS75Xiw9E5MB5OYAUPJmjiopT2WRA9
6fC9vYBmBv0fHNsicZXC4VMfXz1+VqEGxdFiZFC/oNBRnIg6d1R9pI9vgIfbaU/NojOH/j8jvGGK
Q2asqgTVd9a3vnE2zmUN44c9YPz1PGMdIdVaaAHRJijHEVvnR4SVPbCkV8pFyW+JVkxtRhoyl4+a
AnltepuiVN+Aadu4cvqPTZipuZJkJoHq+d+e3JMkLVcTZIOfoFOGJnUojETzP9qaHJe8gPecHYW8
gEmPdCbi1vZZqbCYWbh+1Vb+m1evIjNx79tslIPHVWc9k4f51gZeJS3SrTajPw2+OiwVAtmuqoOz
mGOY3gjzh2fUxTTcgUSmSJt7qxbYT/VZ2U8ro2paqszBTmx6yBXnKFvaUV+XeM4PtmWLu4r5I8g6
b7kaJxtdln0Ym7OUataY8LBMkguTO0QWXgaRcSDM3oYYdc/r4UeGLbz1AfV+KsgJOAqELGV6aRCx
aGVKzhe9kKsAQP6gsHVfLNbkdB88T3+BHnx4KzPLF/tKeMwKLLFrFJkC2DHpHK8UXn5wSYgMgk9A
onXteNPyt6cpP+OGoUrgrhFf99pn0+xS17gxp4C3Qmpyfkn5xqiqdt1WHcwVOpg6bbJoaD1+1b9e
iKncHE8aKkucc+afAW7TQRGyRt1l9Fs68Y3gLKb4OF7kK8kaeoq9CcqVy0znnC/aUQDa/fth8x25
U+N3wAKl4CqfpXZLV0Jm+nn7xPELgbhHITyKUr79DKQ4jZ8NjTAj1B9pLoywNXgRaiJDZ0p9N6P+
XyuGCaab5kxIru5jZFNyvW79EpbTJQCXYX7kIdX062ZxZQVGt0G8ca0Lxj1TAbRvYDxrGeeIDo3F
z1YRGN3obuyCzf5Qzg/vTzjesGK2cftxdHxmCwd9mIke45ggajpiGdcvSOCcPZwBrQAVAm70yf0j
88oL5cvT4R3iv7UVLQR6fiZXV4jRWdKfc7KREe1OEeGs2nPtxqo8/E1VJgliiZ+o5oEbe1ulhvO9
wBx7DHyIlz6uXrzpbP/en1xvAZtPuGb/KjXTxBRUA4haDKppmVt7aO/MTzcqP2HxaoSN2e3Arlyb
UVJXxUPuo7m+nFV4SLajx+1BMBapeghaZfEW65k19PMW0dG9xabn05pL52ktwq4xZS1zC671VVmy
eElMAJz5PVXNvSni1QVmSn17Cate6pBUUUlDSiOMvWq5Yq3tCzhsspGmNk09fF8yulMDae5RGPy8
GkWOj0Qxua73irB+epQSnPvqx090X2898qk8xltxSwMkJgQL3uS7TzoucLV1k1Y+5oKql1CJWItm
6gNWszeIf9S4vOPep3v17eogmOYqV78ZP2Ppxg83JZbtkqFrZSXvU5yuv5bx1wX1dlzmp61w68Og
fDEuwuT1iAFzNopF7eetU8VvMAoA0vCzMNoLfWZKPeG1VVjWstbV7K0iTpwvJSilir/eCHh9Sdvk
kqyl9yrQR4zeIENmXU7WpXU/svOZQpma5f3njlu9bVpyfTtaKazY+F1wRLqL7YVv3zhgG35SMVTB
p7UF2J6ekfOYW6BaoM2n9qQEmsDaREgYv7dYDIeSML6rKDLClNne+tEmdXEAcjafSjawlx4y7nb7
Dh1SU75kerq2KKwQeX9D30OUHFf/nDDfIFZmOMUpSWfdYA7S0nTwX5ACtWjFZ3mGYT0WLM6Gsg3q
tiuaoNgWp94FfVsseWqjLpf57T0VGyaSciFlk/wveIUtht6hTCdN0JVPaQA9lBDu+H7F3KYoj+KL
9JBHIoz5dPiieVoOWicfv625xr1SaU63z0KvJdZ2zsGPa/Vl8MVO/UoC4QavXZi0hQFdE35xzi9H
Jc87y+F0ao4ypBTJY5UJ72ooHypZCKyUOF3hbZGp7bNEY7dVu8tuDrr7X21t74LDYLpPeDlGgxV3
zXh1DF1xzxu6KGsM3b0dtHyqUGTuG4q/hbE/v11UCClEAXOTsneNuPWUNgW/A5aSENtmoWMIIIu6
GqHnC0opKA4cT73zqClrh9lwf6iW75vLlY/1y85hDgSe5bD5NtDY+mCR8AUuzFb8DQvkkVxDDNAn
3N/HqjiWqsZRhFjeb/rUrQ9xH3Op0bwIZetZQzz9VRb2GgS6nN27+cXIuTUpX4SJTU5xcGQGwWhZ
Ao3WmNQQCQUcoy1JcneoXHU4rIGW8ahzrf+feTTRKh3C8Hfq6LgUkK00hE9GKLhp4+VeNBm+JTsg
7Zql5ghzR7XngxSn7DCYa8/5oqOQ9RKwpQKtDv41TUwwSwjQcUjCl7jezRLbZh5ofAtuS0Elcoyn
IZ+JvcavGLIHYJ8WTgUU2+FFr3dVcYT9+VjrN7iQCxYqC+aPERgDgAPWlpiIeBjyoZ3S3jKCXrKF
HiWAKxnQP1zSZIlN8TJLK6Kg+rTNOQkh/hlaBMYtJotHBLzkWJfzUgKrem2AVi5IFUTSoy28EAVZ
YakeY6D/2xUPUXPAveUxp4bl5qzLa+steUiKrNoQN77U4lC4eLDmYarsVODTBrysfP98JXINKjk7
wL4H7pUbvtK7y8WnF18J9oKbb8POsjTbRSO3HCw8pdVofi4HHJ01a5jJ+Gnbd0oEsWCMoXFCTc0j
o7kJYRu2AiJ8Thb74NZCLRcKKT5PopVplbiLL0XIwIS3AaKcR4xf/z+l7oefs+a7nrqkMBfLNU3/
yKwbCkgM1m5kcc6TjMqLQl2QWo2u6h7/vxukd23btY2Kn5RuCKKQH0/klA0ng7id9+pA9cYGCCsX
gNhhd1Is3FEwQGu4zSPPpQZbOOo3YrtK26JXamZk9WEL7te+tDcowQj+7Q+e75C+ViVX9HX0Ebp6
LwSsVNRxntSrOMAGp/A0SnCJFl1Q4NWvu3Uv9ASXGvbFOThDUWIjn/Cuk7drzkReRAvlRB/qZaSZ
Z5ibqkBINkajl2BpWlHEw6Nl136LNqIlf943x7812I20zYQF4PEwtJNWeu1ML+8NPaQgJcFmiFIE
g52GMdXw/71epZFa87KMDutulBSOxNRGsQTPqK6folGpRFqS/85/kx4oj/mNw2XC25zDY2fbYE2U
e6LqxPzve0rwTJapjwmjQ6HI2N65fllQPOt9TPl0WdjRFhxvrKnEOXkavB50cNF3Y74dWww3BD9S
2tapyG2pBiW7h2eAzizq6PXK9Bm2ypS+PBzhvz9qjESNnW4Xu+YuDoOlbmvzl3tvyNlUJ8TcjZUI
2vvOZgQPeAkJyCEU3rSHNR+xWOaphqp1YqcihlTzMJpAn1n46WqjyxqJASEo542TYDkJYK8EvcNT
eT8OO1z19EauZ35DNmUyq6JEeQRFMiO7pfmBEEtf7X8SuNUlsI0SgB9jbUiHy/Gh//RCd2SRJQGF
OB96QpH2OQpqmMUANj5prRHvzVy2QC65xEE9SgF2gmkPQTByJ8vgxzsFvWXD7TmY4hYH/BuFGm7W
J6uumKYZVUZqwOmJr68uD8ktzskbpkZ94s35dCo85pthy/OCq64OqC3fP9dziJUXbo+BnSMbHo46
mVC0bdBh2OD1qatVDooe/TJ51fWhUqQ4BP7TKOa6Kq9XZUa5c6BS0MF4gZFg4qkAg4rNdgbmcxXc
LQjj/MANcHVXb6Noyj21c/vdPwUMGyIPXmRqWcB8xdfFWphmJSIbS+1LpCyahCCC+81qStPtwX/e
b+4D6YW1QUNxYmR3792fLywRJ0F3A8eZByIp+WnZK+nab5hx6GsaHMM39RuVrxDAg/nFmSrjJ+i9
xCmJERgP/fE6hrrv8qMqPIIuOVXSL2Eq6Vvxbs3hrh/WVhhcdMZTLMF4pOc9dU393P60ZfFgO28e
+6FvlRUVWsUz2KCbgKMB1JeejAjjKWvzoHoWU0rzFnR05fnwwiyen2T4F+uMh9PABBdvC2rMosEi
EAbHh7pj6BLLH4Z3aXVG80PIIrVOfbK85bEWyQp6J5Oh1oHDMq75tOloYrYDG9K9u3euYio8tEQk
g0GUgjJisczQQbnuz3XKVUYBodEpCsgTr1JxGiB+LWSlk0VUs8uKsENt1Xp61FjTSGHe6aAhbHE6
0fmlIg14hx/BcW7XlN42hNs3Oi82T+wPNCWA3JDtFnplWHNM8xhQRf7ypy3Y1Np55OT5HO5b48zl
1D8FkdX+a8onsHOJpXBS6NvEuIVJdDkM2AulpcBvWJMeEd5vqq5KQNukinDmK68NRTE6K+XtUPFz
7saILWeEc6ytVw0knCfDsib7ywXgL04KN8ND5TyHyURpvxUvIAuNWvPVf1QcU/M8ShfzHB/4qSuL
Qte9V86HcmGAUnj1B1hQT9MuaqSXKV8MkWTiAXiInuOn9AWge6GW8tRTIJ5s2eosSAVmMcaYUMHA
oP+ulnwm6j7e7WSxfNXfwEjdpxgx9Mg/pJCSqLKa9Gt736GwM+CqpCMxnLTI5KNubyiJeKnq6mwC
D18kcLNoRsdw+LlRKjxB4RjzTCD8yyxYD1OmWGeyeIFypOOxeQR2zwBGH4DwznoCsYd1jO5ajDN3
MyQRfhDqYtiAnk1igwUTXmnrqKkc7VA6TI4PadTjyp3sYXpr3zzR0D8+RUfp7oPty31ULGia6IEl
lKF8hbfjSthWm849AvkOwbtWJglwwYGRSNY6mSh2+tJnUHK/pvjBH/Bd48rGIztYNiWJnsqozoUB
rI/V1ANxW4Jn3/CgnFOB4cE1i+XX0yJi75ONlHbH1TmyHl0bJyg8pl+3IFmFQob8T5lk9oQRI/R7
M+NZbRCyeC5jCFqrEeZ2Lmbee5GPLxSk5lgGSD1Nes1BihBRre0EOITS9HYj2qrL/NSYUlmVWOQ5
WgbFDEZjORKz1vK4uUlsnHYqcP8pbRptW1jpl2KvHwjrJMYCGtR95pjI2HavCXVPo8SmjF0mD++/
bxpZNDZUbLy+c4Pf6Kmj+NcHjm2BOSk0v4/AcQd8guhaj8sw86olJ0HJyMsxtBe36vUt5tnvbdn9
x3uOsfJGvM603BW2Yw1ZjXaZ4Wk+pWFYOb3tHwEO3Ft+Bo0uhMKNAUHs1WesHKGyxNes0Nvrr9WQ
QinTHiFVwHm7Jo99L8/pXNYTEqi4W2BqVt/Sji726bKZ8n4Spl660JWWVoUqk2oG+bfUbuTdVTx7
JVxOsabvYvC1SZSg+w5gpnlK8w/6icrtgZ8nkhpxtj56H1qFsVlv9sb2jrKpLPEMhMgnqrTN2TxZ
b6uS85Uj0/F+Qws05glqAbu9Ke7aFXZFOzj6chb0LiA92DYkVfkJ5dd40YIMMJ26gbG05trA2sQF
JEiIadPb7c3UiHhiPF8QgP3ISG2OJgtKm7w9Ip+q57EhJfCd/JOLrBfuONfkfTkZ6I6Fj48lxo+b
mszScTRWNM5JR2EIELa7EhnGw8W69kFoStGEKKupVT/HK8qyZF/qxn7aJJIDqFLlbcR8j5secDhF
X2KLxxvC5dV/EYuxuz3k1hN7mTHK1hCNj4EoIBGVHrRGMEAwnOu3lAPtLnlhecLnd7aVaSoSjXcL
nPkUbdkOYK3ha8KTI7W0AMi6FmqAgVfpzO1KLI+meHNOaTyieP93gQeNgEu13gILHGN1Ak4MUeNp
gQoMxWJ7nDPcQfhR78ObMSdgMw28Xk9pRyeFXjgpE/FrjJR+i5osbR0SaLImJ2Rkj5Ni5ZiNwQ3x
3PJ5wgarrm2wQdfAIEdx0ssAttvG9wE3AacWKnHIy1gXkAArpPRbwCPiIwJE4g5+E5KkS4c1irG6
41ZYNNFhNWwXw0+Qwf6xKIAkYuGCEVTuL6EI9Mykuypka0QD3P1YedtGdb7TNot8GiGOcjbJFdRx
KyQzJKJF78qgHIENCJxr02Qp34tM/qKhoDeR4jw2LXHHPzbHNpMWLISwlwqTlDOzm1D+Alrarbr8
2+vSptroF5ScYH2qkL0XQ9pzJM25NP0iuv+5UfzV8Gb0roAjqqozlA==
`protect end_protected
