`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EIJPO9OSDMvMNdOLRjwQaF6UWoBQGuoL9zzQDGu35ZPwlaCEsuX2/bXZpi1PYJWx1fIV4fCHJ2uv
SGI9TaOoYQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jR96W/xy6IU1CwVZ4OWs9uQHbt8MxEY6OnhSFsNtb0hYTN1DbC1Q7k1rAopY5R85kliEBsNMYuT4
cKz3DR/nTb0Q1MQjXvFgtNYTIJn+x3l/oYgzda29/A8PpsBi6sz8KIglPS1mIVYa6RurRv4LkYKw
EaTHjYSLD9yqzkfqJaQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l+dRl/KQgn5YC8NdqXiuF3uROWLYUXnJ8JxZFU5L4rAPmX7kzGUXJZnRPvSDiahmvJuv8ANZs5gh
xs5LoEmDF0CFompV5QwULgbR2Q6qtwhrEPfg6MLWV0rRtc667uYFE9KTsFf9JZKKO4/H6DzzAdIP
WLVbf01tBroj4IeWcXlkzK/313rQETBKihcoZIo95c6hdiOI/cthsmWnNjsjRy0+PSU4464xZnC5
TEcE7sJSPGR/fWSbLVlBZxn3OEvlbOzvjiNR8+/H97sx/ei8Vj94gc3yWS1QgQO+AcvptL0n+FEy
JyLr8oQ6zAVfPaFj40vg/JebO/peHp+yKYPY5w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KHbON44TPSwtGlB38csZ+aUEMwCA8EA+f07XdNfbRNzHCWdzgmAoOb7uBfu7KxgTm9Dt8IjH0z68
A8EQUItPb1xEcce3WQRQmtBL+94WCLdFalg3R9madXc+OvDU9lJ30/cmMgJzC7ZqYcKNxsY+MltP
9DTs2k9PQ9HK8xPytpE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wBWhADcN+GmDp1YCpVhIm6ehHfqFBS6YvXzYJFLy6Hbtd4ICJ88jM6iQIHo3AmpIauawmkob48i5
njLAuUbhiO3pjbjswXm9m5ULq7P4Zl16GePbc8+NzBZSqwO0mIMB8wKnwW++E2Rn+Nns6sn6MC2x
zonzzsSzqRzajp9fUDbbOq2tS/NGomoy1+X36PLd7Cy5AliI6CDkRHdS0IOLAwKKtEXzMUbjOg7H
Dtr1NedDgP/xgl72/c9xLklOb+LA3hVkJJO16GJEccChdA/9ulSyPIsSQmXX2bub6jXFEifZQ/8t
ihBzhm2r0HZ75QWpj/gbGRQxM/9gTCkKkqLwzg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WEJsl//nwwFukI7AawNtPva4Okhp5BPPbpvcOrHU2WhmmE+kpe4aQOMO547NxOMlZwGZ/nioOZpi
LrmS2pTou7semtJjuwLmE1hUNq1JnXEjxFJO4V4nyJ54enCYSCvNZDfgVzETNMWgvh00LJlZjybK
m78e6vo4JdsWwhR2Egwd030HGF+WhpCBmJqVrWwK5tEGZIr/dG0JtSC4lyLT4TI0WhfArNiIuILg
4hItSA/a2fFSiFfuPJXYSodzb/CpnIKOqjTcK004JEGCZJcglHRpZxK5ieOzXEV5LQE3Ouc6ACbl
rwBw6NkW9ODG4U4PpNFnPhbwmmQLP3dpSXp4+A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1658064)
`protect data_block
bMfPX2R1tFs2k3nA+qlwsBNkbgx3qwShSFbW1DEU9J0xy0SH5zI1E9Hnx/QWuf83RIOPBwA+fCGE
13QH+yuMhyH4jhttUvJhZ5L5w84xu9Af0cTYnrAtZUxLaYdahxCZ5nbxYEmyf3tC4uUiFX0GMMM4
+MIWsvmE/uomnvVSdw92MyIy77weDURQNUG4XD1citmBfHkA2BA1Frx7TicNpmxqVMf/s/cVm0vH
rRt9q6oHNlACTq0nunqJM/rKTicgEVx44gWXjfF4MbFPgPy/2dFe7JSZzPtpgHPiotPDXxMe4ENi
ra7FxRTYfjquz0uytim1UU17iGnzwNlMr6jzeptUE/2WHA5rWLpLwC707JRS8K2LrrIWsP1a8IbG
0wp309vpKW3zXvLwHMWKpRXdj/cRmJkaP4hA9GV6KrLsFdIx3sDUo1mlY5v8DVRQJ7+zlPKG6SLN
dlTCPP+A/jaO5eRW2xp1Z06Kvet1aL4VDcf6MrznfVXKGYQxg/HQuBOm1Jo9jVNXs1YIuHwWSVqJ
dng345HYrkMZPcwPSYB2EVN3eJ+NB498a3H6bPQK2KJIaXkFs0jjJSgaejoQNEfTh1wm/T+16NQa
VvewzcLLwp3L5ySMj8Xxpv5EDGJ5PwQbtZBgeoY9U1AZPmc9Muv5fI1feAuAb2NK3G2tWu81UqgR
lfG+cX+nvHPF3GDPicqdKxKPL2UVIAJiN/qsjatofqIaol9errlGmCREMT6qW4IZ2W5HzhjER5Mz
TfNBmOmXnwjC8V+pIs/KlgesVgpbhhCpKgu1DeVOhVXUrXnk2lXZWIBeP+DklSYumFiKY3VmrX1a
tTqstp9GgtcXmLFPlfbskXnC1gzjbd9gYNKhqqjDkBDNeMJJPT0ckz/fSOc9gGBv1USnuP1dDjqZ
9+qkBxhpwj2nkC1TIHLzKNz64nMu8mi59CpdO5UWhhlr+kgC1u9ba+q8o9eidEQV8iGybRlTewdj
+ep+5YPXnnMfV/8TF67JoqT3v6i86oXzpTDgBtShqr3CwJYMQXigWDwy4gwElVfo81ELTXM4Rlsf
DUm9Q6jSOuQMrZwPb8+MwqJ9shDMpRdYIMq56gO2tSLnfJe1tlIhnE79tKDlT6s8cRvaF5QjW6ZZ
Ome8Qo2iTU6uYpqeYUGG+6uvFb0unQtbrMOkbvOpZnJ9mqw7KB1xJ/HxM8pVx9CkEwlqN7KBZKjH
Aaf90utmHCKrVH/yzHAHR+jtD/zp6+m7f0fZCf9pWxhQUmpfwscPPr/T7Tk3GMc/FPMeMmCRxpZg
/E3+gnylajEL2GUkOg78Y/iUk6IWNvyJpwzavwCOU7pdypYS6Z2kmClwvQx38DZS2ud89zT/PtYz
VM7yrfiViYp3pmcPSEEoNk4QQMweDTF2hG1GTD6fvSzJ60azwbuLMLFDvK8YYC+p+OsMarEp4LEA
NxFj/GB02HfnPSz6sqtOrr/hz1rmhco/RcxS75UGZPxdGJDvy+KEd1ewkEhKT8hdlrE8auR++vWz
ML/a852/kTNTiKlSKP7HRTCijAH3ksXAIK7ZzKqsTkG6mERSBv+PXn2XvBt9/3ooZFdZWYmYGB8W
9MTpLW1u9GhzjDQZSquRaiGj9zZPuo4mZg9MGy8ZMFa9My/M68Cb9xgs+SRDpfAOcpQRGvZK+2ym
fixJmBI8ZaLL+WzFnn2/2ibhf2SAu2iPkdXEB5rqfwOJX27eX5cxqy0E3RtNeesNvWKyXTYx0NcN
OgXTedcUGZU5Mm9oYLmDcfMI5O9p120kfDiLlJEwyMBLwjiePMghf2oSSCbjx2EbJ6bNjQKjuj5D
8pH98I/i1T9tw1QC9zTqHwxtmR/UOfKrXW0YY+B8k0RRKKbZLbvTXlrnX7IPEnEkE+fQUJAYnU7T
mkgrMFeJf03ZNcm3Hi774TizWJbH2gJdhBg4FSUCMLPQ9GWzKdJYExxF18ho+fC5ucb6670/BvAr
uqlxO856ZIvW8JVk3tm2LJCVsCUXkkfpva/n7quGYBP7R9HRZ7rIQ4uLRKShr21IIc2qvCGD0uGy
vPaQvfZJg3vJhznQXeJTWCnZDMZlHXiTiqmwH9lLOKWCEYmCXVxAT3eQfG4Hv2vy+P0I7c6PD1AM
3kDT++CfzWrx64sHgKTACyedjixcMHmbFtMS0/iYHTnRk59X8u6NauyIzRxL/LiUUvRFR/Am1vg+
c1yL93IM2T/ep59beWXq4Wd+jz1/Owb0xXnfp/nMZ50lFr0LIO+8Z6Pmd4tUQ/sA1Vk7p2WYsjF4
Ca8hjXeChVQqvRuvyhChHOghbMQYt1AuzQodBd5M9vsjbHZcsMGsGOGnagVs16GAfFvIU6qTGxrJ
srqZnEBxakG+/CHmRGQcOfcF6thhB+ZxlnYKxPKJ7+ABECxVi91f28zteve6CGx3LVD/Ylwch2bM
aGL/WJMV6rRhyFJv9QWGK0oHZyUCoFbgm2atOaTNNKiLwkmlA9Ub1O2Y2ogIZFlPejv4uzqaUVEQ
59oS+guVkjoKjlvAP/1+H+FwiwTUeMT2/3iT6i65QRYGVXTRIe5K3xqGbTQSceWzM0Ef2y8/3lt5
S+au6DEDd8S+ayZooI6iNKRDoV8DlFzkVPMvP3Agptv1k2QkuCsDRri2hK5s3PrvrmxCsTWiyWWL
9/FozuNaCI8+/HK8DWNmQmEYO1VgzZOZlKaga1nrdS2wGfyIPSr4k6bLTXOBL7DDuUkK/hvFdhMq
nu6ECLh2EFjuiYnmvsqC98p0dgelPwDuXBCs/iqUZ0OMo8qZ2cydsfewbvHb1rqye8l8LXok6wiZ
U+Si60NEH4N00nl4GftbfUKvE0xm0y8715REi932VNrPtPeZpKOWWuq8BUOWuj9/fUY9YHRDje3J
91wVKsyZ7dmRqrWIEO3SJ4OZLchJzxx7kxUmA6460/BoVHcF/ZEgHoX+qElW8M7Jqc28KEmMPqSe
CtxVZn52u7hOJyRPgTxAg8bEdOa+z3z6DhgCqjW+rpb+11CTjZtSoCppJ3sD2CX0pPXfi07TRjlg
MOa02eLF9rmod8OF7Vc6TjkxfBCAcokfUGkSLn+BkGmfzjvjBOFc5GIGFMc8W+I5FzdXEOgFi62h
+od2OO5JrN9rnYPKuV4I7FQmknNuSkY1SuUT80nBcZ7q2sI1D2s27gsYpkbG6QJd9DwNYRhmmwYT
KZMGyheY+iS72+2SZO3cOdZh6H7pqgjrLQ4x5G9AGhzwrTRXmERcE+Gb+pLk1l1fQweVqJfGXckc
QjgVRMOS6szlXElrBXtsn6vISIFmlJ8OG+ZFesk7r8Jr094ALAE/wemhYHWOCJ8w18se07sUcHKE
JusTRdK4ZNReJd45xsssGjb5COtr1YnQkzfQUfPGH9S88IImto+ABNsOim3ulnlrhnfQ8bI3iVQW
6sg4d/3lQKm3fhZSoX5OPu6AyNPjNj4zxKY1kb55gDIXk5i1i8VXQvX240ZpV/SUjUhuPGuCzZDe
Cl+f+9vfXGPLnyAszN2my9oJLGdJYDPAP50eBMMfyTQxNghw7stMGgxjizhA4zdgfRUvKMfqHZDl
DfWToVDY/YrVgTC7ffgmswwHGxGOvP5kCEWvmOt3DjMtOVuZJbcMOkrQHG4GbH4YLMGqQyv3YyMV
zLwDAMnalxe/invP4zeO2aKjD2Ec6aLjZCmkOskmlX7PhanvbJlfG8NIkRZ/fOTgS0sOsEVIFRJH
XhvQbGXumwFp263TXMZYvtoXbBPbTvIOaeJeaEUltrV0Oit0W80OksPPsGIqEZTPQLbXP6T4ZAjz
9Gph07WflIAKrf1zGZtsG/AWPghlZ40snCCPUlVrEKhdUATg6gC0C/8iQsz9H+OAAGH4SOB8GrDB
4bFWdP9K8SBacYAJiAjUEgmInpdvBrx/x0p/3jZIhn/9ewkhbXktzz9fSZ6xvkzvZG6KWmgLOJD6
5tuV8EiG6CXT82LjNj9nk/4sWL2rejJh8xyfkvPI7FNG46+EdaHfUg3eYQrc5+2YvBTkv03Vd//6
RJPlN/yhSYyz9ywGkg200BSEIQjkDybDcjbvDBVChDOFkwpQFuWJz3Hq2/wqVqBKEmU3q1O0iqE2
5qYxTlgWWYfamcxCH1fnIcz4OZ9f7RWy6fqNWs6erpNy2jaOiMVyyc5aoe0rs9ycpzgPjUVHbPJf
LuBDxIGf0zrp8TkM2XdIPxcPS6hG9PdL7G1i7TknzqewhHNNvwg+O0l84tZEcRJRRdkRLk/mykCJ
NBXHbx7JEfyjF3Rqv4/0ZWFMVF0Nml/uOKXLTmWjCKHuJcsrv4kFHET9sEkdPFRJeJZQqVee3UIB
J1VdCOYt2k89K9n5WJqAIcZOr6TGdWHdslUerdth25DEAOw23Vc77IznqcVzZiKeXNx+zB2vrqpv
E/FqlgZaMUPvM3wb0ho0i2q5p9kA+B9ZI/WVa0Zuw6NFrtjLVrxC7hYYh+8PgYtNZZhofa/ZcarM
ywAJjrOCZDZkvfvLS4w6gmZgtFghcbqUK6ASa0Dw0PQD6Ev2W0g9ohbOQ9OCdAeqFFgG8/P2ba/L
Qoj7wJjC7lcGFLTJXCPjnQh3XeMq3o8YQweg2b5FjVZO/jt8vX0vDPTRMqazeqwKvk2frXN8Dr8C
oEeBoHWCbTnEJVhzLwwx0RZ/0Fco3ZM9WsKfMjO8xFEfvr8NvN4nogmHerKtqFLY4Vlld7rX+R+G
aU3pG2zPx1R0z/j5EoLEDwYW9qCZ4JEwQrHs9grIqqXDuXBJ2HHlNrjVuQGciw4hShIjSmbmab1i
pCsPtZ+HpSkefXqXR4JitZjOUT9CfOE6iXH7Jh0IAeWW6+JjXekW8Wpx2wEgLgD5g4nzeJOImPoH
HS8MHEN+ToTDYZUC8HsxEUv5400YvtRZNQbXo9Y4t9WmDwAes5n57/0tTcGwHovXQNjjXva4RtU3
3a6hjp7c5KoryRp/SMzBcjy2LnKLva4Qt9w/GcsmUkiFV4MRVZf0iTaKILuAuFgjGrCHR46MB02J
J7vOOJbpuNUkctWMkZjFFeFZaQmKeKLMlz4umAK4OMApnHpeCZFVt7z5JM++Nk6AdPOkHBn12eVl
kWcdULRLj8CRGQ/LYUtno7SZxhbv8yO+aiTP+WbjY1SO31hR43kwlRpXCLhuKnBk8i9+OQuRbQV4
8UxRLmdUtGZEePUoLh1xcYHTKQTQhnoIfblifBiThRzLGgmIiPb05UzneVgbVo65rcod/MxaJKA6
OJpF5gI3Lmz/k6X1kr06ncQH6U82YCQTliiX++6PcX9RjhdoNgaW/sSZdzOajlP6FsiQpJjckmEF
BjmCEZ9aNDg7QYunrdmetwdD6TYTBsYys/kYclaICe1HHBNx+rXpft3dgYByBAvz78mhsHvnrdk0
OCV42AsfTTPSpzFtAi25wRuAQH++OnqUs8ygT7gdvkCIQ0BhjstLdLHDRVFhwmj64VsU+Axptpfd
g7q21uvJlnnRettOPwJyzTAG55N+4SPcGu9+5q3bgoiPbhdKxJ9U4sybvvAf52HQSDnXXMs1i6kQ
9muhvol79F/0Gn99ywvn3bjIReF9APUXRJpjvpb4QRcF24LqhJhJvY/VDoXch5hMi9CNsR5MCTJ2
R7wP2Q3RTfbPRfqlFidbFpuRP+YeCUQLLud9lNGkhqtCB5W+6KR4SU1yK1rfsoui2l05XskEh/Rd
LP0X0fAodkXwFpXaN/P501ADv5w1GK4si4iImy12OOGjmfRzcye0SEBq3tks1MmOBLHqDzu1O6H3
URp+Bcq7TjK1HFKelwA+jgY0IHt9M2TIz53eA8DOfLXT66uG/xEpoh5tRvwzeihLvJZYUxKmzR3b
gxuqXWuLl2opekgQS3P8GwLOIW/2J2q04ju80q4J6TvvkeoxIwAewVwNqS/4co1IytfI3mbEG53n
r74QxwQ+tl7OVDpdDTP49IvIl3tsZgmid93AMKxXVaUoYh732AeQOYNjOLbpdwl4nkracgT0deD+
mch7mVFbT092fIXxMmIuYA0NZI/GcGAJi1YlPMLhuEVz2tMrdtHJ6oRafDPst1L0I1N8O703WuEI
KrciARCF8pDduo58W544tjEoDYJxqcWKBXMpLM8BXEOBXjUnpclFckisH5WZxhcrbJG+S4ZNNupQ
r+SVrxY4MEzmgdloHFuaOvnsSk1thnX/u58INAil/LpxE2bjaui/rjoqrF5+lSRXmW6eTdKy+RO/
cXyz/BS7bjD/vur7OKNonReyVhv73ERyWuN0oBnzt7E49uOVjBxQibylwl/x81Bby5xG08IrBzIZ
xbYSmohtImrlISmvsEQqf99NBxon8MpGi8kshpDUIXggQakNr+x8pLog7/vstLmVNrxFhBEMzsUf
M10qmudssweKONkp/Rsh5qux4aX9E6U6sUhvSGK5z3xYyTzBHkQNA9L5zisp6WsUye3kT70wP4Sb
E2N285/j6VF3DF76QMbo6mZ6cZCyjOcpmZUaGEJAQKwXZFf6XCkm4of7RLX/98N8Fc0uhofnZMbB
zX0W7JWS+LUBno59/HKEXWDQ8dxaYP31mcT2IaYFIEc/mChZ18infP192r9ZxcHUwbmzkUGCvD40
XumqZS9Fd8xbp3kwzLbp14NPHceW4MwIUGO07XHif2/iWr27B+CwjkQ5MTH/6qg/Nbk7Ylstqems
87Qe1APRzsFJ9n3CNJkwvat8yfOlcRdz+b5kPyIgrp1kn5eesSDZ9O40RYwuOfGGD2PvrDPRwsIy
QZNrOo0beXCers1Jqmtr1qwW60PGvR27FKq08/OzBpouZTmsfTXaeKG5KCXHEL9sqC3CDN/ldxa0
SsoNzb/HY8HsEZZem0+qFv6HKKUnobJvYuWZH9LXRlwvewM1loiEfJYAj4HGih6Lp5cTmvwi/2i/
4fosviSSGjS29aeG+q6SbrUghYvzYU2xiVUviJxFlHnaTlLoCShqCmDKhdai7FTPTjT50RDFHNzw
NmL/d/0FdozDaCfLBn3zILB1pt+uCOzGlJI00jBbR2vgWaD7vqjT+2dtRWD8tOyOl3gMx4i83sJd
CtYjv7J5rDuedgPC+/0JZ1vTgClEPX2c9pEXTUgLnvLGyhGJjFHuacSZGBuNh0X/loj4y98Ce+Zg
Dvt5YSJPUZS+s8Pq/hwwpQqPKEKzGFKGNnqdxaKe8vWkcENq+tna5RSxmB39B9aV48Btr2jYik9x
NyhyF7Y8Ci6UEKfLIORHxoikNFThr5+smFnMifhpZw74Kgv5hKHSYXfZX8/aUMYBNFnvDTz6WKIo
hk/KDiN5zsuchUFRLQhnb1DMLcP18+KnbgYJxk69qoIgnxowsetsVygMeH8a2KM6IP30x9vVMaiJ
bCauvkxF56LsyaQWleUwTXNx+eZfsGd2/zxd7erEs5s1vxisrN0197qIbYGNAvrxFCeFZlAu/C+z
IBK+iLSielfGNDzrBia0tCTa/C3qxbypB7LftkFW4h5j0mngDOWcAw9qkA2+CvLLeGVdSndcfwtK
vZ/M48Gn6IZD8TwhxapY82R5F4Yk50LdrIiG9CnLMQNMWf+RRnSN2zwdBlCCT6meR88E8OIltN2d
rZFiodsiP69GuX3Gz2j1jDF9bspxr4GxAR0k7M7lNFAQt+FzPbHyZ9SlVK6vCUDCE/fxGIxLX62J
0M0h731tK7G93SCMV79mMHMnNcbD7x89hWWfEJWJIe5e0j00tQnvQ4U+zOEA2kUTkBZR66hdV/KY
C+7oCVl7Ky9BfXZYMZt1rl2n9Ob/IWCwVjmc9lGJV5eDzW3qM1wLz3KJHm5FK+6aRcGSdy0VwJU5
A/8U1ODuaJ5sy2sfOvV/vUm9giUyeykSQMpUwj8Rk8kvO7SiMxu6bKC3fTV8OlNbSuDYMcMnlfB/
fI/WfN/ffOtG2FAdCikLcmXW6GbAfVd6d2/PGx935/YOwPB67/ywrZp8vJiNEpKZRiuutbzQ7V22
O03y36wPShE75AfpeTVBMqxZ0T2i6HI1KYZbaIbE56rc9wX33fxr4xw0zIC80jxFY0bjN42BEnyE
0/ctpMNsbYZNgbJfuTXzFhIiZV6JjeRpnLTKm5kDj3yM3UM2O1GFrM2x4+oiLCTaleaEF8HsuaRd
aXTuhjay3XrRJyL/hSyyatVmkdkIaPWMW+tt5cDIDz7s1Cjp4DK9BeMgATfT5lKTlSQsKB0pKNwn
+iARBdsyjWAAjcOwTuEySbzYltv86X4wg2nyokZNR0PwiJCf4s3f7drhW1eHUT9FlBNsxV/rhv2H
HXqOJSJhJH1JGUPDb2VjsP2h6QOKEyqAtzoMKjS1R92h9CgC6oJ6zIYDa3JM7PHq7nWlwj1aDXNJ
Aai6YgJpjZMc+9V3DT6lQzeW8BFM37X1XFWPY9nPIcq+uBito7dSRimN8xCfH4ErlPP8FDXUq8v6
uji1exxOmvy2csYXsJxDVfm0aJ6L+tjntgUvijSt1r6D1FSs0KzYoBUAAlcFLu33QzEvx5fouPEA
9rRoZT3gIm9l31R9lvjpb51i0tRUPqnYn/dqadKY5g6eobgOuoTZ2kQYatzXW9VKuL4PpL7W5t5o
k/EL+5KqlvLyZjePINq4x1TnKbNAzbUEpcKnKE3iZNQrBrU3uXTHlr4pf0qYe1DCx1w+Dv1pDO2A
iS/gjVWR03QR8ZqXjCH5FcDPrz//oxFgn3moejd5bmYMBYa2ThBX6Rl8KnET7DJmSATQNaFJdXRB
T1Ym4bXlg9Qpio/mpRSkQEWdjwgSTScWav20FXTsxCSMqbgPQBnm8ONqSj/PYiNEVcjYAFubT8PZ
n8uw5FN+CE/9+5RZ6E5oCoL1nP/ZTcKKdO9Mj616kTqfQS3Nmb5svhWzMzeYw9FWWnNr3wDC3/PG
wSSXQg70aiqic0ECICC9e5TuX2yp8iXH9eKTSpB4qBGOCsniwJ2QQOMF6xnuM2MxfoRYaSHeeBcU
280FoJoHWn8H/8gntlpMcACqHdn58axgExwFuDOOb8kpISF4TLH19/5hqkQqqCug1ZGRQQJRPRGt
n+1srocUGiIg23mqW3eu9mHMkxzYSJm/0Fud7Y5W4IIZyfoF+hse3DZLhbNVwFl/MT+1zsSugGfp
Had1la2Z30WyyHsSMfFlt9FTrJEDbzW8xCiyvdK1q09oB06tEr7iBYWBASNc+xkMzcIsaCb07HPs
lcc5lTxIiKktaulSfHcVTzu7Y44kmFpADzmvDJc+4csggVWCZbwZIRIAx/nFg4Mms14Sta3Jem2P
d8aT9bCqr0Ma0/u/3DQUPt5Z5h+IV9mDJm35zwBVpMisoikVSYOGjDvtY6VxjhhHR52WWsVNQg5B
yq5lAZndGv0Dff5ZKcANWQ7077gD7x4MqFoEalwnK4PIao5EALg41w6l0C2DBc2i4jXrzusbcc9Y
5TGEHY/M+z0xH+jjYI9URpm0YMJuhc8zLoI935/3tXWCin8pqabt0InkQ68mUFOF4h+bs/FrN6Le
+vsCDcVQUIaLhy4lZgqlVLhGhDnuaaFdw4jAzmZN5u8qXxR++L6FZJieIwYVPhFPX/ikKUnICdmL
YzdnqrUAMMdSdi0UZDM6d71GZiPxElQiXVeieDE54jT0PeBP31hngTUZoDkUHcLu3cf35fqU/eku
UmCd/yPJRbuNqp/0czD4KFj/sA/j+5DaaEMXDUnF5FnlXbIoxL3LlJMEKU3WNPfleb2LQnVR5q3c
9pfw1NegaoPnwOwVXtTJ0RqOUVVY2UYvWk2v3lEp1kHVC58GW6cvMXvO7Yt+4lOEotfuEFkvDPhe
dMBFHp/E3F0I3H4O4I6udnHs7kqlqMZd0+UecQuKaQjADrfy6r97opszSn1r9OHBZsMOTw0Hh1d5
YN64BpwFjq7aaVMVCJ6a5HY9JIspfc/v7QnNZJyk1CAaARCrCwmIbodRSmUvRLFCrvb1SnMiNsLv
cSyyZnRHG1OfUN5WkCtFbo3UXg1qNjyT1cLVfRik5lD85Rz7BvPc9e4pG1D1hM2lr2etwSZzvO7l
N24QOyTZt9CJ2HLskCBTzTo/SLBOOjf7PhXnS7+Dm4Dg48Doyird2c+6b0zK7e/+la42lmFHpR6l
N8KJdmTA2VADtCpHoUaREP0BeWVadGmEvOEscQ0KifjqXj2SDXviiUchcqVKGwCQ8Yr2qIZrd4sk
bhMKw7yUDvhy0TSCejF0oANn/DSgq/ye+YvecpFIHn32ErenV6V1cbQIUPwLsdwvi5qcvPXAiuKN
IS2OJol2+NcMb77+nma70fqkAbvNM4AE7gnej83qwpxnJIfyllc+V5xmh+iLp29DXPqe87ZHdTC4
7VphXA6IYN7RHbU9hfiwZSnfObVXN6tX50ODLEHdFaCDgsOUeLQlC74QRhgVIu3Px/8SPAwSbacq
vHiZmsyjXhLgNB4tWdLceeeCKX2SaWTFpMjp4B7QDX0p8iye81nmYQWEO/uBL6bZVR1Eo5W2HvMf
shNNroR0XKtJVIRVKGZaUrdNoEK+NCvJHDxmcWUhO/kJ5Xcz0TjcwAu3vAHq8AqjR+CIDmFJAXCp
J+0M9zLR60sfYNmEY5Vd4/pvW3YSAWLPJ1CGvV1Yd5piVpSlfV0t3UM99BI0MG2zHt8AmoTAsr3o
MGT03eA+AvJjUAR1EQNiqdtK5DNcuv7kq8BFxX51oK5C3LnXjRy2cGy9eBOU7j5csYQRTm8J/YyN
rVmPBJKNB6sZyOcdzP4J5NT91b+P2NWrB/hSKAwgdCvnMIdaD4DekgDIU4viHRLReffjTkruHAng
uoN2H6zbRzSNaZtm9SbGq1UXnqsCfNhjhOYwI4WX6d/mTZRucOo0g/+TTfEijhEOYLAdd3pYtd9r
THYrp1AyW21U8qKqfg/okiLZCm7CFDKzaKjuChUDWnNTNEcum1okbfLBDQTkNyjoGqS4SE3Tv+A8
MZmyMfIoLRHBpl568p8/mIRdcKZiT6+lfeYKIq2N6Exxy6fEHTBULI1tlNpRKyXw1H13WXSdus57
32sBWGglxAu1B4JzGo+iMWnpbndO3HaBMHP6gmRLTxL7L+5y3uLwymcj5swWFtA73PRu4O0cEiu0
tpvwxwqHcOeXros57GMxkHZjuLHtvvbuLJSZc0v6xVqOuZy6GWQ+1SOxo6t8wVxnaeFxIkZMv26X
pAq8Tu+Y7/YHPy1fhABzk4Uqxp0CRaiTr+DPh0g1BdUB5tzxbM1k/2/jSqmNcUGvVuOCwjFf1Q61
jCdv0819y0ykGrJI8PuQuqrE0hVG13KCNc8m7Vf0YwdaaCSq1yQEjxPEX7IE3qCa0Dx/VXTINUDD
2B89RUocZZYve+htEqn5YYf/cygX5Nx/KcNEJcvVlNxHbY3+0a1+ZqdmUYY+MXCxIw8hIZQ8tnh3
msPg3YH5s5bxZvRCjZWPIvsOEfch8jYEIulmgNisveX+043eMR2ARDtIhmJHKVQe7Xwya0oaOPKx
7DOLV5+X19QiZ6kpDiCgQTGBxwt7RH7Op9G8hsdB07wDeaRt7zgKbJojJcWz8yvXRM3xDQW7YX4v
5oaydW/XwJef7aKoKIsHidWKwmRfkF9Yz+OI8uU6iUaELty91BLFT2pD1bWM3o9gM3mhDBCZmbvN
6XUdbbITjmygtp2L1BYb9imGgyLcVcFn8uAd/Wl8FhCQTAuX8URFki5Bv+cgI15bmZw9zG86c8YF
PyBSgGUCKdp6q7RhAgbcuIxgZsaDkGL5IsvmZwdWnEbrLefd3vZAIe6El5rD6mNM7niGn4AlUtov
E5deeusoBCnFfunixmexBxIgGdAUbnYX5nWniWa/KK/n5hjlC45kCMODDoTBqVY4oea7u1SzcMLJ
tLzX5SkOlq5IE4KhcKAEgjs+g5hSTv0yufNLbXBBGxNXVw7Mhbq1cPs82CwvGyOCdzCl48GDxEP0
WZqfY0U9/xrUCRDmcw0EYmcM5hFzjjzPJlVB4UX11JkfeyjpFC3YzqrXgSmzgWAr8Mc6PdOLkKSn
o8VpuESw/fPEgCEdHsAWAHRxnkSFpAuPTqDvftgaTNkItBIi7zyxQsDf2L/LNXyeD+wYY6eZm/ju
4sej2yucPC+wn5vlDYehMkTmcc+B4VSSDjIgvWonISYGG/aM7Qh7IXg9YbPuzCoe4IvYsSBEcnRy
ViYtRUJwtLV9JBOqlzQajEHtvNeEDfmLLFsH3+HXKoBSR/NMRQeXZ7gOlZR+NczQhaP0fS+AHNjU
w6JlxXKS0roIXtdcYbcIanvnnalF0KV6XokFGFohN6eni43bDJHEs4rVgRv2jSaIGICUsPkPyCrv
Yy8P5ymoH3c4UZ7D+xTYdb85dMbX4GvernXOZ1YWK8lII2ox9Gfe56Av47xyaFVvcombyA4RLbO3
kM6H8u1WExXVvqpgQO5wmBXpDSsF2EMR/MSLMN/kwDQqaBGQC/v/ZoYiaRkP858qhG1yZeOxg8mB
YSFy3LHvW9F9i7SP3MbhwWtyQG/uiqy6DFAmmzOxP7cvWIpsu+hfJnF8fk0Qq/PF7BNElS0R+t3l
K70uRham58EelpKiNDEVSsEXMjP53jh7JfqOaBZuQfBxHFpUHJ7XS9CzfZCnI9D/pYihQKskZisi
tz1vqLpCPrnmv6jP37RvZGeutRuYoS/qwbGfVDq9zAsRjYV32HnFV8FSJeTf8Ir0SJWzg6mHw3jJ
Fpe3GzDmfF675/Y3IdIMUe/bTvM57VNZ1OSadRD25/H8rN7z1OhMlebHYZcvU4QMSJZTmHfM/zl1
Z0eJ5R9HVFl2UUHNCQRmCscp9ornjemyMlNLOVGwao7jrbNZMGQ+RkLuUoiLFigNsFn9+kuc2mIU
AE3VHDXr3COtOMhatDdDm14RMwKwYN9lk3jMmqOogUEI2FoAZgwXirzrk/ejbyfdHBFpxjy2USHp
n+UjhfNBxcD1Xw2KO0Dg36cdpUtcdfQnIfIeBMLS3NhiMmaJnPXQJzeDipAlxaGG5KI8V/A3tkpZ
MOG7JDkNfvsiRecbTXDMrx7ns8HGZd0zPxsXTg1wDwhMeoREWssH8LsoS3aO4GOmsYTwGh59xw3z
8An+uxKMm/8bFk3jB1Uop3fysFtnHU0sqpKUFxbEjLC6K6ylSj1VYhnigksnENiQEl81lhAxAuil
RCVR30bEg+IpZ4CPCuuNchvW/hA78LBNpA2hxO3pTwv5jIrjTceBUGTDuASoJ/ut2kY55MJ2htRb
ppH0tiekGK/YG6K5kg+t90B6jNQxIKj62R4Xr+BSHMQncGUtPcYfaNId9De7GRXTfpc2mcE3pCwK
oOOQaeus3lYIeo3hR9StB9+TjbEaxbzHjEcES32GDCHilGjTPnAjqhiNUqz01mYaTjqYnTAn6oqX
jP2fy5+pCcEL9UPbhZ09DpyOmxdojDIRGx6uMtte+mGvixNpJZvxe+/CzGlTi4jUIJhQYjUlte96
Vz1hNMPkHFPrjWg6Ow5QatIA7VpKwP/IZEGuLBKy8B+/+QVg47crJ7aoFk9I72CftrRwNZfGiAHp
BAYy1WF18AX5EZduIcf3oEKGnk8Un4OMBCH7StCyK0kD++yim1ydUhUD+SNHiMmtFeZvZ2ctgyZN
wk+1B0FbPtmAuvYIDfGxxFXp3oYyeCO01OZ4Wp6EYmgxGy5j/fIRMyThOwqCnMyGZcDKQF6Dv/Dk
pQMOu4bbqpvLHeMMncdQvveUR8li4e06sehdBjm3HG3Lyit0jgvCxzL8xtQ30IuUiwUnkO3lAr8B
hn7S/BZQL+HdCD/gxJ4aqBlI18EeZZoeKfRLOGx62RJdAOy1rLx8f+zdkSXXcAtvvPslyMk++6Nt
Q9M+lTOAJabTHkBUDqDKq+eJ5gV3yjutsl99SGYs+/Pv2YZzGbt2euPW5xuOg6+QT/BNR4cEiqV5
ZwjwUUk58S1tbTGdTcW0ikXZ/smmj+/YH5T6kxd7viGvQ+cPHTPxbhwZPafYBbe4yPbY0QsgAflr
pEUhr85oPkCnxg49aNrdYg+yQpnuHvziQHMEk/sMcwXxYSTcGeNmovwPp5zbLPUKh7qAoTNTtysK
TR88HkBdAdtxfULZDlICHYJIFAJvWXOeCc8ejjBp95kClKK6OqzlGpgEsB9dXAzFoiE0Gn3zZUyK
cy9gr7RlDdFFVWNN3vjC44jDYUgoVMseYN367chg/INd59Rj2abGI0OOd6DQbOEcWUsoxGhgCatE
epO6mFEBmotAQaxNlIxoHs1+FhgakQniDsdp2YQ1F7DhPdfm869iqac1Vrw8rJFvitc6hSsxwIvJ
Wx188qeRkssPXtlv2vPsTxBK7jPT1X9+CIw7JdL9n8yUEybogoCfmgvvlrT5SARgTEFuBgKuJMTf
v0fByOwyQc9kF1nVXgrQVEstg2vYO05017smlC3z/tM2OJdYxkvAfPYBDZ9jhZmEjiYkx1+ydKAG
wqMqlz+6YsBulR8siWWpYOwJ6JOGEptNE23Ek8SP8+zVRNbaZlQi2lp125K4DxJi34cT0SJG/GT2
coEbkLYiulFoGBl4vAUlGUJtP0Yypyd7QmKhE6gNUvQDrTAlDsd8/hGzJ1qcA93nJA3S/q7rehK6
WjpUXWfCBCvYdiIe6RJuKzwlMMWSmerh0MC6XZ/wjfn/im1tAZ29NeTHHtbHkpLifkBgFKWY/qaU
uE95HviwrDztwWfdouCpnSzY0FbVBZiKoL6H0LncFdBZqOLJtu4JoPX2/0fWctMCWiMs+Q2RVku2
ZRt4WyJAnoJkEh2KJF5cUpAemYk5Lrpzoe8WGWpHzbt8Tua6P493r3QEAouQBlPFBjqirwjP2dGq
+aD2d7R34i/LZn3FcyT8dT/0aRtUD8STmgYZv+uzukZfGRKnXIBi2JOc9YgVceyxkqUqlqptGOPB
R/pX5XQHwIpuIS1EUzNSk4ffr1LwZnB7M4BhmyYleDpTv+bwNaNZI6EISTXBzKXHnT1XxbVOVC9v
mXi3CX7Q9c0FDbJibI+EhRGJh8Muc3TB+UXtFhQx0QFhNRRHwF9jdRsipwU1o3hGq1XORoXBftNs
B8jn+ohCLPEgusGj/yqZdwkAtf22/FasvFXsKAvC5RBNJO1FD7m/TatHxH0MwV+yo49oRyI4SntK
CUYBwajFE81P1dwxkweueXgKI0y6DK0IOnzeNYKc3icDRRSbWgOtXNfyx8ccay1gewv170c25fnv
v4Mzox75/JePFqa1XVgnrifKt7r2SLvFuj8KQbihqHSnAjcEG55SMxxFCNvrJLCZwXNjMivL1f77
RJnm8bOU8OUmBB5uNWM5bsvu+03Es6U62ki43qICooKRakQ49aockNUcgqbnbjb4+/3g4Qp+bk19
dBa4Bpx5uDv0/8ufO2XuUBVRHut8/iFUcZGP/PdBewqVLWt9IDmND+qsqEtCSr3a9vfNfVmTWUXS
Mx9o/mqtxK8ssQD8guAdDER9icQ96gNbf0m91KDbldYchYlyaqEG60VLCOwxg/ubGDWlZGAI8YIf
BRML3a2FE0J0JZjYBcqBas98+gc4DBfROJPlWJwZnAXaNz+ro1p2iUOEtX++v9s48tBBhg/Gn44T
/g27Cj7ahVoMDZbI3l816hVA5/Q3Q92yKxXDBmL8rmr9whK0+vyM3s8qoIVxwU3iG+XIMsWBQUtK
JjOMzHAJIYbwi5qEDYfzi9nwgGszKurHhBsci0PZplsafg9zdtZVE6pWPIrX6e/wFLOEd7Xjqv4Y
thcLDQGBMTbXlsHR1vJnR5SrfsSY5/bsJqOvawfAlbf0HC7TwZ+oGAFVQLSEcL9R6o6dcoTUX+JM
pZ1S+5rhs5Yf/aHn4QQeeiB6xxdNEPunKhgjbbF0HUpzUds4oa1/Rkzm/YNf5W+4GJNKniX40Hkm
hLXCijk8PLXrXRHAM4qUJlcHo5zN8joXa25Bf2q1ftyZsbTAH5PxN2e995u6F3ykmggaZvZ8lW18
xHNp5BR/kqg8er0J63I+BRcNmMOfyp04XI4OTgvYQdK1GgwxIfbXZMWRrNDnAuh3c7o8CFHYnObH
wOuU5dkREl6KY7eyzhrvZC69M3x6D6IMp3qQAdvfkrynTNoJAGKo99FxhWiYut0ot9vORD84C1+D
OxV+/iRmyANwrt9qng5xEDe8O3a8Z+w5U9rteGlYWi6hYp6Ygahp6i3qVI0liUNNVzaN8+Wut2GS
vV/TQxnsDBcbc+8Kq6vlsyZizO077KtkrUaXjRE1/O6wfPYL7kNpnka3ecOLkp+bSfV7RNAhEXvw
XEoWL/vxZQfjI3ZLj31ao3KhzYiIhE8v8ucQ3/kt81FRABFMw2EIc+VXxiUGkwUB1ukb37CSbxco
rB0MofN1a69wZOEYLd8T2He5k0lpOd/T26wxtYgFGCSi3ImlGwfCXLtWKttF50DNHIRhrsi/xFl5
NVNVyOnQYNLOolLul+pQb9Gf5iO5qv0GiSdoAfpP9EOqpwZKT9ATqlwJ2t89uY4hLzWxfaZBR380
iF1mBSUd/6cvB+Hk3o3L9DEQMFz1vw2Xn3XmZpzUG0YYc05ChgeueZKL6LT9pKhqjeixsGM3Yyz5
DIdMy9r5S83bLphRIc9d5TvCuDQbNE5jx5Cy8C3BrTTvaAXlwOhof/6166dNj6Y/U+t0zUcIgP/5
jyOORXmcwg1TPvfR8mO6/eRcG7ZhaZjwhtgUJriZFRFlcbXnRDjX1tMF4+PjKJwYSUL6yXMPC+le
Pz2buWuY0kvp9eONyf8tdCqnJ4GXs4olEQxV/DlQvttln5eOZKLGWnQQ4JGr+zZX2QQsRr/vmkBr
i6xGA/8lYCyFwgFKrn7RdXOVGNr5c3EYwxKWK1Hqj5fRyy/GjeUeL5ys+0A/AKaO7vYee0fK/6+I
ixxRKwcWdHSU3//0Z5bYF9Ju2WaOoQuyZxOyFnoRbD0SjYtHWvETPquDaOFdY/6xjGLE/SxAbU4E
XabBdP3Skq0vIbaGHdTukGP2FN1COuYbXkQy/pzxzG3sR0t7ncKHoo59e/29cWD5CemAcbovm6Nm
TrXvMXoOjU//Bqm+i6yW5JVJ2AMzU/0a35Q0n3+XyKGELwNIGgFbjJXWrD7lP1Iw0P1X8GIoPBWF
97f9UmJmelwBBSIuP/Dbm/FM24o/YTDrmg0stneIH7fgsTHa8+d0oSQMvvye9cE2JFfvIiQlHQY2
0jMusBJw5RzQfrxZbfxaRTwN6JlIFztgSAv7nFwR3JyUcNCB2qtLV+tZeyr7SFshTKkRvvxEvyJ8
DONlAygMxeuGfBt5tHWNsvrntncMFo8pIcFw22tFndha2gDX5YmpnkWq4k749kKZzRHGH1bNYBMX
0mIP0EQR3QxQYCKarnEbBy53/mdQoND0JNPxatp8FWS73zykXoQ3ylo+rPgRYPgfsSRS1ZGlZQmf
H8J5y6y5RvqFc3tu2xiF8kd3LKlPvmls2wyMBNuo2vLze4zvRN9Xe/IbkItiul/hqkzI+6j/eMfy
kDNN/6Z+UWByIsW7coat2R/7updAtrwIecqXhPv5f/iOv/sXbKB+8kv5xdy3xGFI5wqkYVA7UNm2
hdn0xdqpzWDsU9LDi05SdW1ZTcL+q2+LJ1iUfHZ4bd4jpCCGqdnP81U7+k8h6vsYR+RD7tsYsg3G
4PqGBuv+Rx5Fo8Ffd/nzzudsY4DYIGNAbyqJZklOMzvOxE0/BIovP3GXHWQq8aDQQ/IVdn82T6e0
YqkVuosJy1fy6+NxMf37qySbvC3NLBMqSKFTV6QbmZPR+APy46k7D5wy5vNIfg/e7m+vFy4IGMnw
OJp4cMwvJpxrjM7WP8jiSqo65YYfHc+olo49d0FJ/rYesO58RLDtqIZnHki6Kf5LpTt0Y96x2xMO
/Y9fA42oWQJA3bz0jX4IvUNO5y57YLaOKMSZqGKfRBb49N5dcHGFEhaAIz3iru+ttWe2aC3p+IZK
ZiMh7sZgWz9TxBI0xtoW9pG83zxU5V1MMxkG6SsNbubWCcn7hQf0E1vXTL9u1DgOVSKU5NvYEan4
u0D/x+bX8BycCgOQYa047mHud1DP7X03bDLiD397Hv+svELKJ7Of9CR3wpIF9gtht4nWSHyI0XDT
TK6/X+FLVUONPjvPOvbbyYMlHWbebBC40soENcnFLYQt0bT7XZtCRlpKRViLFEW3LhsFiqrafQBS
o9q1My5dW0gH59XB6ufc4hivWwmZvk4KvY6ZteCZqz+FtKGHlngP1kfKfWAPGg8xXDSvDoKokstr
XtbLPHHVLrqmAlbM/aVCA7kuYLRqsWNnDdqlYEFJvE6A9DiX084InMbIWQsRXeGzUQ8T4fY8RZJW
jJsMoS5+2fb6D7DJ/msU23ri+C/wUF3NECveNFJV8UiMkoJKnWhgh0yIeTnTmh/4f9hVTEFfHSX1
gL1360xLEGU/kOod5OCrT6J6TyHMRJzxr6cnMsD7Aracc0u95VVxKDoNTKxFVlnVTGj/3hNpdtgy
2qVev4ALGdfJ8wKlRNsU2b+1RJrNC5dncsUN5+tXvdFP3RvC4gmu4beOouxYrb1LjSmTXT3nXhQ3
mTDKXMjMF0cpntIUwAj2DbGe98Gzi323OUW7nBqAAqaatBN+qUuCr7ITZo79ESh9JyvjQ6ZOeXu2
zaeZ5lpoWZmwq5eUAPqysL4kyhpr/teFG0u78FplxNUaYzgZAmQECTsDIozTaEsssKOzSSvClPIF
axDIXGyByDj0JsbCNqnBF2CY7lLiu/LhFtOh1dpTGcM2MrKGb9fGQPfz418BaMAY0ExBS5716REC
YDm/c99pMAZq0jZX4WovTjrJH+zzPhBYQhMpCj5PRndFdAUmS3kPcMZ2ogqS3+Nd78j8v1iv37ep
vMsR7ULxyv9GZ+2+cvm5X6bZKk522Te2NQ/FuWxd5Xwnhih9duJb45FUvMwuA0GSo4F5qIS91b5K
/mVDfeT2FXu6ziY9H8GtcHqMhksBduJiThPN6HjUgcrruHVUZkjm8gzTH9tnpBv/bVlOQh5as4go
dtMHIp/RxoCfLclv4eEK3EXk6eeP4FBjkJlJHsGBc7B7wv6gjRi6/Q17OQW6P/279OqoPNO5qU4x
cjKnVtFObooKcS2gF/OSZFiNYL/H4c3H9FghbHWzhRzqnAmnvBE2LM9AVpD1mAcl90AmqXCUr+Q7
d3dfUAlERrPESuYdkX/HI/zKGW2GWtTjaKyuDNJNqTSJAe1ZfXYWuhCHIdzcnRdEJbPrV3P7JTqL
lqedTeEUz10caqUDrCQbQ9IvddXXXQGad58l+HPGpMvNHXTIL8M5gCiXaoAfLkt9vt34iTC5Y0CS
7vNJu45qkSuJVJX8+H854eheLrwhRvDnLp3NEQQfGxrE8wAsZNcESyxMZGqK1EllVvo6K3Aezst4
uxqUELfGWpDP+h7M1K8q7HjsLEA8ZB3HR/TWE3VlfkfVl1Kiw24mR3EHMhX/IE8+Fxn8wfGC0ISB
iQ5zwo33ewLzhJyEwfmrpvszzCFX4IBXh3pnus0BU6ymBfCLaXwAHvoytsc0VMpZ/FoaRd+zjZSe
JmjTDeOhqSE0Ll7GVITLP3kD/Uns5ladmnpDFtAdK2HZaJ77UatDSjPbnhT9a4HrI7MznSfJuhBw
y2xtUa117/QYy7ELytodY/VMX6dc5dxw0CYrkpta719YiIuaAUva7RzBqlxEg8UIQRXNRLCxCYTc
4fWpraP7IMn8xfjYYDSelVaFlP5sb2yBvPdgzh8YqO2/IMUEzxA0lR2XKjT3Rm9z8StDtvEpqpLm
EvNa7/zI5PTh5VNSSjkTUGBapPJse4Hb18x9xrbVeZnS2NjaU12QoXU4B94ivCNUcKqESx5DGGV8
NFZUieTQlf7RReCC203tmYjZLC4HJQPFExtmjcgozg4rJW364PVyED2YtvmX1Ibx8Vx6y910cmUi
4hKaQuWTx/4oaAVxefW+e/3azX7O64k5fQ9o2m7b3lZbrbgHrVmAogAcolAExsRqzt08GpRr+fTR
9RrrMq+d9oqYA/8bjK4P3scV1o7E/c69/MKxpvLoYaMQlWJGuQDNPEFyGO0xPsoCiNu5mncSbArf
rnqMSoPH9p1+lN+hDmWgk/7f5ZyLxykHepF4XIXBCUHAKvlYbTW7XoJD5KQOuIqZZ2n2kAXKNDwA
Z4/QwuHYa6t6cHSnpC7qnGSAcUSbG42+XD1OwJnGLnlejaL/L/Gky+QWKQNg968W8p9B1iRfdGNI
Q7CJXOXJcJ4z9kwK9AnkegTaCcx26FXwCAXz/Aee6wUoGX+MmQOy/V5EmSXmb8IYYul6MWqVblAO
ll43bAZYnF3wM1QowrcTgE+6Fx5kHl8SqfNTJT4bWsrZtkRguRcV+J4l0qOkq5Umx5BMV4bIYl99
RbSuBzBwdrrlUh8tZBB60251IgVejm2xn44aqh0DPJfxFBGUDGh/76ripYeRw0Zx1OnzoMQgRcDC
tge3EE+x0uPY4pWSLnyXx1t0Z6xVr9R7hg1cufRJ3TWoAiureYs1aREGlv5Az3msHlvUlwZdSMLx
tTjBK/7WfDFVPPQwvVN/lunwX7xLQJoVEQe1aAS5jPA37BewSTGNpWpJEOxJf8T827tZbOtN80Hv
U6T2/t+uM/Nf0wouVRcH8ml7C10qnXrpNp9aHt8pnwXUkIferRCiGekfaat4uhANZkxfcUceN7/m
BsfSRkI2ZD2H9M3RpCtF3hNm+TZbmF9UTHaxVz4+PnYKQers2cBYGogrvwcCRIrkU1QKoeC8TfIm
d/RrkgoGaKPnttPOrp/E6KsUAGL2DGrej0i+56KHJd4rHwtKFnwAaLJHSF2VfwgokU7owRukOzwe
am2j5QO1L7jQmEEb/U4cfeU1BXKtHiRxmHvL6F4xKTBvB00CeN9nGJDiju+xq7Ar3gAMzd01Yhej
KMH8H0ishgOm3B3esNjwBER2JKDcVhHZLgdmoMCjiSHwNx9fIrGCUcgULk3YD0adMAkPFKkNIuby
XbPLlGXxlF/Xe9k8tysXSUuaBuIpMVj0SpKs/B/gDxVAKCvk9aYvAWGtkK/grAHdCLBNi0Si4a1/
pwVkMcuRCVEG+T/2aWxF8nvxqK9cPg6F2KaW97RHzjVUQ5GIVPrGjkDvrKvsKaP/F9wgn3tlYjyI
QvnfGHOhdKFiswj+kfL8plEJTEG/93lpV7upKowsjj6za/1GI0AOJeBOoM5V9NyOoIWbSFSdWGtY
p+Ze1O7ptds3YJJPXhOFu+jUAvrlFSQhJPrp9ZtboUbcGDmQK7f/npYoXwI3XvOXhqe5WcdqZj7L
J/nmW4X/muhrntgVrJaeUbXrXiwxz4LFwRczKRGkfCvlRR+FK5x8J/PGhZ1i27luqIq/bUtsv73b
ug96OHi/2drxzlKHvB5xXQYcYg9/W64k1Jk1+90ZN75fETwoQFSO6/PIKM4R7sX0kdrdxsDvjF6O
fDVsnRPJPOTO63UOE34EHAbKOYkrSFOsPuS5vcw8QNgNmdKPqUtO0DF5MbCpBDukAf25uLQ3crdL
KcucCsM0wQpsw72gb7l7W4bUh8hr7lj3GGVS3vtXn9/a93gU7Y/KchNgQENUkZWkaq1KBPPU+GhO
Y3JWSAYDZYDtajTWYFoHjNmjjp6uocLDE0P4hQdLFd2wcAev7CQ/1pHdtV5N5bve3FSLcC4hgqGo
AOEnWbV2RzQTsDqqt9jR9MnarFUYi9CNkqCmSTHSLyx2AC9ei6P63C7y2mDiF0ELl2WQn2gHYnkQ
4UycTcnvebUVKH7R3HTQXQQ+eeffj33OCY1DRiSa7ZgDqsaPkxkyRM5ptEdmkPDBX7kGJgKaEvOu
5WDcI5tjOUB4PYYyRdIyb4ZyEz9F2Fk6nisI2Zvckq6Qhoi4MwHx7EMtZZyOOTPNEmwI4hVDmkNv
OGllNgWb8Os2jW9QTxSk9je6qoQFfWo+ILNf/r7+CvSTIvinQ2Ni6XpVcVoQTw9ZgSUcOeXrwkYG
FEup2LgGcQPFcjUCvW21b54g88ErXQS2mhueIbnMUMlRczZ37aWHnlN3ocnHBsgMsxzQ2MFrpJ6K
TXfSH/auuXz7evf6DnDkF9j9hU+q/xORWKMCaoytxBLyuy/SBWlOLj6LpD7MS4zCnm7ZMn/9ttji
IgeTnCtKdaTbNV3BKn/5ZWYOpa7uySJDa4rtwy2GYXVrg47DEj2sct55AqLC8N+V/4JMvyH22Hre
HyskzCQiQN/Gc35/R6Bt5zCAEkK2S/pxrTx1tBLEyMr5rpfEEJlo2bDtJ12JCcS68yiWdR+BtWVy
o0IRWbXY5a/k0+3SqUdM7V9h4W2A26VEDx/QwHFKhsPfODJ/9F9bK0WmuqVu87ApCfuWiUSDXnLq
NisE7z4IH/nrAmVbIBvx2iAymL19b2kgniILsa7YdSHlSs+gftroL12IlHFUwXqxccetDogI1+8e
1XjpbRJycZTN5DikvAPMiLmid5MCELBfBaWSKbordzFDVfN7zDrXO8tLwKn9mIpPYzH41x8EZH8T
n0x0Vf5OSppnElY1ByAEaNc+AW/7sEOvdhWQKYRAQwAACLgj0nglAt0Lj4Ld661anjXCRMSMgwSU
GxrpNeE7xeMJNekw5GTjwmaRTT7L+fg6sbfi4p+WGn/xnfCgUtATY9KBT7ZRhwsX7VrzhGaBwwl/
M5AxIgzyqgNvGHHiW6UdlAhBk49NPsHUW6VUI8j1vS/TfwL5eV6d01VFq2mlbnJHddfWAQzJ/zpB
YkjupFyq4x6nVsXwEGNzXTisWgX5P5vrGyQrRq0qLwAgzcG5pPJ/1GM8TGTC+BVtlbUXhNA7OCJT
wSglrDDKnMZv1VndhxNbhEBQAiCtSmHJ2Cd+qtG9QILvtMF4zCJu5Q9p860uHZazb4tlQuLcHq+B
NSDcPrlaW3mAhphmjLErMYJoeRVwbPFBMDYuXCNH9s+GG8dMAQdKB1CO9QIcNHEb2+5pxlE7fSyq
Bzh5GGHP48DglOoci6zbKEnhgDYPSMQcG/1y94GgmGGi8tTUaUeqYJcYFChdo1ymPH1dLgqdhrxN
UVUPXz8E2LXccMi7fwz0+CY0ilK3Q3dmIiyL/ByNOgma0hmKg/Im8h51mGQLTe5eZ5iXAuSw8MOb
4QkP2FtV39W8plQudewAaNu1gyZ8gPeuBt92/BndECJ8prUZzUmZ8I7OutFcTJZfHXJmxQOZy53U
NX0aGClYGGFdB3m5uRuz0P6ak5ony+Wa/WUs4+SHH93QHYyG0vqKLFAxd6NEQqN8fKE4aiokFaWt
OwQ3q/JrQ84v/vtZH/FcxfpRSIZVVlmIQA/k9rGsKKTKEz5JLEZBLWm44rj1kMK9kLGGsn/TzBTz
NLJTjj89xbO4fMCw81WknjRJxRMNjfc/bTYXBnnKY7b7EI/XYg/5Qa8mmzYS5M5LArGgXXymZhv7
olwFFR4TRqb7qOh2dM9cP+hfvyttGyCntSPPLAZUweamExQPgzn0OJtZU1ALQ8LIDQ6N7utPVI52
05kdkaW/AYdu2CKDxLT+SZvlrEWo72S6bUlT7ADC2TdYh0AfOODzj1T01NaiQ7UyORzYuNmevydV
VU9rRYtzjQik8NTKQX7qza4eoaIr6jHjJNilCHoXoZEiAPCSPk49VmNeAoLatQNKBaPZRaB5rJmx
HIpH9J5boqN/xF/zJtA7FuwUMwdXF+oNYOXkxqNNpLY1XzIY+TxAr4Zygde21fg6M7mhcT1SjzAp
ybt11fOvZCnQdR4Vru5kqhKmH6xWfSy3Imz0/yHXnOBILS/vC2lbNR0G/r/vG8qVzOiXoj43Dt+n
VaOJZyQNFJ2EOQjeg5aHmrsOw/j3HtYMYKsP6yw2u+ImiBDsKaGbwiNa+ENiXsZiZKmt/WX8QQIU
9yTAw8vrjXRo9h+eiBAsUi+K2iJRcRVfzUTPpG402ZAn2Uv5a1epFa9dH/uK0ZwhFqMDJktmo9Eb
0Z1BWHPH2ioM7f3pv+4JOcTKD5ByXJB1kO+O1oT76AwAQrZLYeMLrRScOdiEtu5+SgTLGHapaDtc
nK+Tx+UbeZf+6+MIBCo2XN97TTbC0XQVTkTRC136g+bZGuPHZa71NEHMUqmOIZgnBA+4y08ug/S/
SRwsy0eDjVwmQYqEbIMlE/fkh1mwLXYl2r2lw2weMwbeeNKBKlWxaldEuDJmUFzW6VohO5OG6SKx
3KzF6SRZd00P4sPcO9YO9f8DlVwfK2pAHFeUBH1btiZGKbttamdLRfShnNaW+qWFdWIUNnzunIR/
YVftGCjzStBSv/OPLPTZQ3uWqZX+bi+mSjXjiJaIzRoquhj5DQ53icHUfyMX5tZDxJAshP4OvOYI
t+c6u0C5yohAOOxoxIwJicP9mI6KW93iV5aIsbIajWuvDwWpDu2HNQ+BLsfI4RuevKoFfwlxYGtt
//oHlsgTwyXjUdIFKgaer6j6RCLKORB6JswOVLJUKosje68VdhtBRnTXgFF5DDnMe4coAXukLQCs
cINVzvlg+BvtEkzDZmCY5i2CQrYMp2AYR2RG74uNqOyHWAtAGfX2nsvB41KQ6B1cSlbREv9yA6bW
uTgTlIbXiDOIPlR7+iWteI7cPp+fz9iOZrqJOjEJAH8aHGX4s+hYMtuc4T0pqyWcMDbl28byPZhM
cBP7wpsD70Z1QaZPpDbp4rrKQX6MBQq2Z61VF2690Zpt1lsfDKxvEoNC2Mc1mOIkrpWFtZW81hGi
Zi3AvoIeXpk5NIrpqQF9bUMQJUNo00oLNlOMwZ5LnV9jTQs+yQzbq+DYsqH0OsLG7rwcchzF1POT
ICzwstGixS1kXUoNGn80SgruSgssdd6T4IFBrWKGu3zUa1Mh1jdeukMvz2hV9mHIcFoLiqtoO22Z
60BMgthx3CMvpwbkrWaAFgmkKVKLRumCd7HknHrEfT7aa/r1AWnYmtsAKqeMyufSuoymWZBUlKqd
nOUjq+Th+bUK9LwQZg7Gn+jpmr1yA1wmEeXNFYjHPyCVxUT42XnC/bWLjtopV9mLvfNnXF0cCnoe
PEq21gHurCOh78y9g7PdL8DlQGbm1ZtGhu2gSsu/Hi/O9fL+mV9YTKwhz7a5kZ9uWugyj5XecIiO
gqfp6kGhfANNtoxiYaXwKo9mkIOWCL0Td48R0JIqjZtGeL5mU43VEHWNBhBMNRye9BLDA5sTAevz
lJx9+i3iRi3t9o9+WszoBr5PkrEQ4YenP0pKQaykxwMyu7VmjMGcCPhNJ1579g5c/q9nvXiyNirU
XjRxGmImPH77SLdRAw3PChFgXz6iFVOERgk8DuntwAhCftcacNm+pRffXeu16MbuCJEWEVP95Pjj
O3PY697sXhE5TbQXvUU0i5GAQmX7NgRfng8Yrw8kO7RZjhdt6UlpL7EVwSC7Etu30WrXiMHm7zaA
kQbN9xZvAHV060KC44FnxAq5ZnWh2M+qtfc8yKDhgFDFTPVQns587cVi3JF4dR8H/zNzVjwO9hMt
Ju53Nlvq98kclHhbHl5zX71+sxKyOHxhIOv1IA5zp2o6jIR+fEHuGJl/OC1g+M9BII+4AzNxpsu0
pOa7jwfuNxwJTNfKFD6/s78fgZLQ9vY/McAf2QDOmt9Zgqc51yfbfOyHFpZlocwX8JRiqcpHuVUS
36YX9WXg6z/t26hyWkLh608QYqS63J7Bk+FO84BDq962pFrr6DKe30pbi1y5NAbzmZu0HbHVQBra
NaT3yyLKba5dPevI1Ik7bMURWf7qq1+OPi9ZRuKmns76TroqZK2W2bIUBqBnTWzKsTwtSPNCrkeB
f/184QrzwJuF0fRWmEdotafH9Ayht+9TNImO+0W6FNsKWDzeqe5hGRvsO/yqarwBc70hHwLNZ1P/
THa0DMTbWxSjXdPHxjtESCfpp9LKT50qmtwLlnZVHeoJDnDLw+h/uR4nXq+LX+2sdA7MvjLLt3NM
H13PAPikDdtaQe0njbI+LR4/6lCSBURAV7yGEWelDyQ0vQoZMz7uHOKZ1laqbgqfSUIhnOkdHc1Q
A8q8DZL5/E6QlAIS590VfaSJ5oF0eCmJvXiRzaqYE8uIuPoNaTUfyYIaMGa53gOiXfvKmYJHp35K
4a2VADWbeO2XVk8qKQVUcgwb1z0iZ4ws4H2SPWjaDH+utJih26TPIc6fc0cmejo40QhzwRS/5geD
3w7zHcZB7MTJ0mAGw4NX2GjcS83jPcl1Ro9WHPzCx/ug0wIAzzAY5FpJs8BArUKhK/MgOYNrmamQ
YEW4uSJ8u3C9zX5GkfS5BNNXX6t9yoIbltzKuMz9p0EsdMyQKzTLP1sL6aeZij+c2motu2jBrEu9
XuBn4G9rVciUiFXJbOvTP4bikp1fm1XO+PuZElVk+UTftWxaSYofmvT6wGUX8BJL2rLeS3YpZsGl
yuln03gpAUpToDBj5NbXtxxZ4iAsc1Tqf0nlP5q7I9mXMajIurG451+RTkFxmhZVoLgDeYtBz1Zr
KkeQvpYpJoNiQ6zwHL0ZDFPPlAi91+1Okn3OrGTykg2wFeBoJE9AomfpFGCUtK7BTvx7+0Ro86sv
zfCMAUDxJQrfCu2JwDlpJynXGGduJAg7nQEw+mDfap/LNAPgsDk7rI1iKC5ZvVKmszfGTZpAluGR
qqKStxA3ILQR9Da2znfkMZL06ABC8aVpQzELSA3069BtiX7ocdhwySu++j3hI5WsvTGYUSUb96ov
5HM8EH52tde1FcPJyzYzM08NhG4FEWSaFLi0jC9m3hPLq//V8G5OX2syqoMOS0ZxWgz+umZQiLfR
c3M3f76GOED8NfcsYfljIiydovw5BbpZr6DII3rI/p+k7ZOGHwwpd4MMK1VEFMFlo5MglHrWA/gg
RB6L9OOlzwN21pjDo8DqOqBdI27Y+ncQd9qN2Sgihc4sSQor7ViNqj4Jas/IVd5cPYqK0NIck0lj
Oj+4OzFDNxJpUUMPFJ35tw/b1XPXHkLWljDceg5vg+Hk8mdqYRdFVDDB01ACvL+vTnZRfJ+JrNt/
6Gdz/B0l+tbyCZHE+ME1QdcBhldeJ11pfqs1kfe25eIm9jcWQinlsKubsYRUUWYs94mNEOqgcNj6
V58OEp9ECValqELdc2pkOgdUUmDYY5eycIB5Kupk6I5Mv8CLDm8gTO9/tv50jV+8mfrVehMPC4T7
ULqCDwfNLShwa0lIP9wwQQS/cHafPReiGnrVLAeonpDKbA6MgDtfZsOkRNYFR+1eELOawets2gAI
HkxvMnBhReY/QM2sSk5CFXRXU+1f4b5SLJF3dYI1vFx84Ie/bevZaAlZEs0b0wvvPuZQMXCND0Q2
HfanKYqUFT07CuQdLm/+pC/CfB8BauzDO+ey+MUPjFsvBVXhyA4IS2bVK9zG9ZLY+U6rDoRGtpjH
2y1C5D1t6X9sHBmBzi/DM3oKe28CMPxhcfsa8BTPhIcTzcf/nxhnZ7U3ydvVKn5z48c2eqJq9MD3
Oc1IfFJTMPVfyq7CPgwhA2L4rQRgQyfMk2eGWhbPPVwK2QasVJYofQ6uol1vfKk0TS3W7Uh997Ts
aFL3FdUxA9qXe9JTiiVRg2nJzOpDIpGE2lPiWAIz0N1jVEZi532xJp9HUDJ4LlaiNlZY8mGmdSt8
0kEygsIkAMeCT3eh4TEo/aMx+mv8dddtzhpCKf+rQXqgcloJY1nOUIZ2vXPaDHIS7P3mRlsjsc1c
TB02MxP/yaIvML0tNYxIGhMsQHhpwyKAytvIBIHf7eF869erhRXW+WGC8NOG/ZY1VLAi6mlxJ7TH
sthh7RXyFAYkca6W45OYbhTDs6rks7BAuVEofdyaLUtQ8So/4KNJiLwO6a/jzj75fzmuNPFeYDt8
s3F70UX5IAHliqKM6K9xrighv4Pov4+bH3ukA6UBvCg83tTNjUu6AcIsmHlKkMGPga9hshctvhLd
EeZC2UGX42aEiibzwIu5crl0Gu+bRf0e6nKy+5RnCsHHJIzl7WYq6mlFRjTHrgQPGk1+yUE9uE5C
gbIfmDeL7JzI1uLSq0HDYqNgBKvELFHQ+RWikSwNn7aZYL3uyXzlI6BL5At0/VsHA6JAIwXKyf9U
rtN1YeEzK2ijQoArNIfyncnmzdXl8yIybExw6eZ/qb+UgPelCjfpepWnhNdw29KlJGnz2GOQrtL0
tVdUl/ddufqywcCfHu1qjGo/WAFxa7a1ilJdaoPWuTYsrqVKg0ZeDjkfOyTDCZUN3n6Mb5E6hAdq
al3vtHBUSlL5+s7hqPSWdE0kzaCBb56ENCSGwJd5DEuk5NWQiRVFBiVL12mELCvw7YEZ0gXcYUlX
v7vdUodBEh5tXSCJNTy8Yow7Low0VZNA7I4bdO4rm8P1RYMoFAPDWHLm39/xSNChphRsZhvPQ7+f
xvFS2auTaNAR3GLhsa63qawuinp9inPUgmLcIXDc9vT390xBjEiucteRbeI+5g73ZH4RJRAVHyB8
TvdTXpfZAQgSdtrV1i81q+6eubtkXBPSdEP3O5BVBJ6fid6uoMODPoQKRQqXwNYBEGn2yRUT93+D
cWIowUxB9FmWkUugpKZSJbyHcZtavg8lCTBUuQXJO+zLWBjk4vGY9Ij/0Zlwu65Ha6A1SdJM8u9r
QHLEq4cPknXuH0EpGuqnRi0IUMOhc4tsSo2pHKyJg/fp7TRswuxabKkmTDOlx19zxXev45auMQYf
xvh9m88sSHX5ZhZ6RgBmBTE6nzWlNSwd3LL525qIzPv3WuaRHwZMB88m0EKPhk/qCaQ0qXTHgPn0
WqMQ+wZwKgbc7s+ckisI6mFJjjwWP8w4Pihn8xbxZAaAsO9BY3mVa1D+HJZWOGly6uHrKtEguh+A
ENK30YYH/sKCoPUh40NsLxwBOMHB4XBgk1KJ/iz7IAzmpGf41FjBoejb6ufpUULZLwEItwOCpTwR
bOcvUxfd5hTAqseOMV2xDzcmSXtGmAMZug5tItv7+57BLncV0vtk4/fIOMT6MBNPulcHOOlo+/C4
N6zZ1bK0LlJ50lRU4mGP8CkeYTV9Xrv6QAZrmWJ+erFyV26qb/x4tirYIB8nQiAMsqpCYPxz1RUF
e+nc1H8EzdSgQ+o7whhzsjRo8SQwH8+Aycu1K7IkkhQ2IwrEYjXT9MDypAj/2rsLnVfOpGUu5DBT
Oc5kGXdGp5rXzCBb8Ytm9c7vOrHet/fXsZBw3eCsAnB4enQZrlJTe2XvP0d/tWORc+t+vYw95din
Nkam22QMI+qeOg2tq2A5ncT6927q1RBw3WcfODLUOz6SsWT6hAQXbYIYDP+AmaPieen9nkGvK6Q0
KH/rSBI1PEKeUJxSC7lo7Q58K9DVtNTrCvpyf+HIBdhAuDEpWBfvqilzDImOEYKypyAF1UYcf2GT
pwot5TsEKq9Yl9IX+L0bQU1KTX/Wt0JakwlJrbsf6JDg74dDoeZXhfANv16X9IGiSMWPA51kNHY3
tCbHZQoNjW+wuyFBEjbigpFADYWMXnx79EQf2dqKaX4gXfm2zkYoFZh+CF5EaNKTM76Ect0wrNJe
KedI2tSGhW+mUGW7XNXBfW2WghhhJOglxfdDjCUN8fOpMkHwPk0grJh64zjhOpJ9fGusgVp7kaJy
akRaZ1iscWDYonMOpTqqpnVMA+12aB/mSM7NHFCVPg9jUYJBGxZL0gFlJVxj3SHrIF1FJfOWmuV7
cqDOS+7MX0pg5E9J7FMwJ2efA0WJOTU6mFtf5+HP5+V1+OFlKQgoGosLIwG2pwzHvS4XkrZcdPS6
cdpZfmqvkaDTdlkCl0wwOaqTMhQoXDgC4KSkdGylc31ya8xHGF2FtG4bzOigE6fEO/KrzFEiFKIu
ZBTKpcpLminmmeK5mWJLf6WKf+DoEWBexlqCNuRTAeg7xujdaXRHve1qUBK87OCPmdGBNsfj3R/K
611KFaKthalsHvxZedkv+L09tMokXP7sGV6xXnI5Ww5SU5r+mdu9BRmqLtwpoXzleLetsddvhAHH
0O15WYdbiqbKaGzFo6j9JTDwolKjLVXgV9IrG8AZ346dIAGhqebrWKHusD+z6frkuwEHgNeFuGW3
SMdl6wHAnBJbelrMCILvgN1EL9gOw4N3rQp1qcGXfAAFLAFRQwqbQenLC4gedLpH2gePrUG2NWsM
fo5UZc7KKciaKHZENOeKaYf2C6dGaJNsD2iqKbBOZCbvw2kz87fei1U7v/JvKy0Oy5hvHrQ690qW
xjWSX/v/BCNrll/RZn02Sm/RAbfra/lY7RAcRI+7ZOMFdUBZgmsKeyWddIJJw5+HJnT3eQ8yrNyO
lQzwrj64Sdw0rVWcFB6GPP6BFZ9AQiC0b0QW6GCdNwecn3newf5eVjdit+XmT4I+pFKXGu1BPG+j
dO9zCi/nYxKqYQuOM47i0B3FrXvRu1hsln24K9ipQYncTfd3nuPeOPEp716Y2ZpQqOizV3Ic9Ogy
sCuxnAU8syIoRYe/zkQPeKuwf/VG4aytEyQlS5VmoCea96YlNkldiJaZfxyYOPhlo5MOQBupObpZ
mfKV+WPzeOw6HT+wAn4gSucnZ8aJs8ilh03wN5LajuFappjOZ/1I/MlQNJAs290y/M6WtprtpjkV
LIynlVspCm8pGNUE3YjjwFOpJ8GmJXYrKWwYtwG1W83BNbKoULBwl+Ho957ZcqK+0D8gtI8dv8Mz
/fDWMpeVmTD8WNUM2mNCHaD8wDOdF5mofG5yuXaBRzEwzVy4v8XVbGM9upoyVM9ystopFWsA3JTP
RvnHZrfn8rJanSyWn0gVia99xS0FaKn4+4f4WG6/tFjD0b8QsinPvauW+RhTbuAgVMfuHDSx0d5s
jG+encZC93wQxaVBN3JP2TzZ5z1yZP3exwtevbErl1l5OnFqI5+eFJkCMAdjliZpXsD+IRnLtxiW
dTIK0FGVZCqWJR4WX16CCbbfzNo5YtcarPa/SpiLnuhq4mWnHcTyurj1Up1KrMh8jIAMMAtd2qgT
98ZfrKxxg8v9iWetcByOn7UZHfPQ0Ru3dsj2OnEFqIV56qVem6wZkszWJk8pyXmG5YnDd+Penxpr
UaxTFEs5yw8xNUKT0rKezuYKGT8xPA2a5uSw513OWVT3MTbreYd65UGmKZZg4hSTTrjeqAGqdaK+
Yw5+vW4+tmaGyi79eR9rhpe9hrm3tcRYxEJGYBuHJy5pWI0xZlfSYGNVvtjwTnc+a36hEJlpALsb
tlwGMJ7KfX3dEZTcQoeN7EoEK1GEZNh1lM7KriUvfFPt0p48WZ9pm611p8ejJMWnfPc1Q6gCDfD0
NHc86rEZ+15AD5s1qqtfbW/nDAGWjcfKDfC+T/dhD6iXu7MvldSkbz4SuM8YStmhFBk0C54KKbDb
Ieuu583BpRHeW7hIHxZFCP3+8PsD43AdfgBLOav9MAqMyWJkT323lFkMVNJHYffSmwq0WjVV41OW
8Lq0KryuCAXJRpkNB8IQQzfG1X0Or9Ff9YpY4aYw+OCpr7ef3Od7NYKvBMFlIjT9ddZ3wTssGA4p
YZnS7BwTt4ffM6oZRO0OjGHKUr77iwf2PHwyijDnSaUDUX1+Vug2TP4RaZgQXNbJVf40NftgfUvt
sm1rR2EerCCMVc3ZsctFK4KSeE7a+HUjIWPXOwNguk9VbHIqaeNyHBxqxHlDmfDBABRUDScDrosF
sWzZ08wTPsmwzXOWj7m/tcgG1cTRfmJOk+uAlL57w5XbZWbcqlJ7kOVc9BusILkVTtxze4ogxC7Q
NC+87t25nlM69StQ7SPkh9STbY0qPpbQuHBSo4pqqiA8qjPiFCV07m6HCWiuPBzSWZT3zYXZZJdv
VGgw+NJbJJxhfHdKRL3XNKKwGajn19vAgrpEW95o5R/MBbGmnaBjVrcveNd5xtHBEo6TgGY89VOV
VSI1Z87/cD1NDbILtuUlwzrxbC0VUVrhSen5T66KFAegBWtaSioTbMertr34Z1xsrLPS6J5ptkxH
/TO5+NSGf2SFBNdFV6X1mqEBPF/k5vXvYpMBUnb8bAaVXmm79rygs/DqsOHWxpSdv70l06lY4Jxd
/74V28ZNkMfXiiyCxV85NGj4VBFjp22Q41TvSRQ++Vmfw+vGjZrqRLlFpnb74Jn+APHZpyRsTm6t
VkWFe5JgKhNEMesK/GXP57vNJUboDhgEqt1XnQY/2gFmGS+RwySe8FNNUbrG3OvZ2rgVsdGTCEsl
INXqYeKF2aH1v7/fcpWthWUBCfnGnWlbbvduOIRuRnIlMqNnX1xg/ETf//X5Wpo8tU7d0jiZqLy7
4F4ioSmCBrYJb6hIttSUFdxDD2lgHUK4i3/cngd1LPQKIL3osMPOK/v+QGRkuKn/ZoqBRzqs2Ma5
WZuzoNvzoU60ALzVlrnsFPgSHtJ7jjl0d2+ImcWJBD/5OamdDz9kcOxPkbTBPxa5QUiZt7GiKqWh
tiR/ueumb1zfK0uRstilNtb8jDvUaCspxG3s44ooVvGGZYRajuInClDBOMBj4HeNUqIYZLgqGuWG
ZFzqyO3EUU1pCIcojWxhKHe9KU4uCmzU10J9OyforQwf7K3RNnF5jkhFMfa/CVrPuBtQr2UeDPv9
7NML8MBANMJl5YZyiGAQ1MljrUxrzJ6ag/WK0JzLqMbeXv2tT+G+oA6+IxEaK7F8vn75M7NKFm4t
na5c4x9f9ujjfE+W7ydm44TzhnhTUO5ptrGolp1LriFG5YZ13lBlS5JMyjdFDL/3zOFXHi8uBGax
/5vo2yzEJFzmJ/qhzHMQ/cA+1w1oimtnkURHMnOsKS3UUPWTU2An1KQq7VAaO5E2mB8IDpYqV69Y
9ZlSZTQ73Nalofrl2oYP0lro+s5t4LpNI+YbU0ZqEU51cT1r3+O7kHbrytu784mLaY3S8PoEbE8W
Trx5Qn/EsI8hol9/rcZIxt1e6nATG8QFcbkDOBiuKQjCvJ76dmRTaPS2+ZGfI6ras5Azwt+XXanE
lFoO9xcjsUNXg+FTpE//e9eCt5SsMOfELBDnuQA1rv1YH8sw1pBi9WxHF6F1pmuGzuWvfli78HVv
93ws5kp2bgI4uA89XLNZ+V6a5N4HLPTE1DtGib1DIkTIWxg7Ji7xSqdohr/DcagYudO5wbpj3Qec
Sm8TT6QhEFt1nH1KORSPbp2r26fThGuVjIF54c0EvDfs7blc88Bvpgfa6Gl7mawJucqxNVMfmBap
+4NNWxQ943yqT8B0MzWWpiFSE8/6OaTWZj7C4ZlREM/H0KTZfYUONLc2am5Lq519dMCmBOSHfyaD
zWDtV43tPqfT8zE918uwP8I/a2Gllryn1OxAsqMtJr5Kgq97UywwcalFMvbHe82Vvo8seNXqx5wL
uEGofNOTU9hszZubgAHlZS/9mSdV6hGiOQuNw5pTAfvtimNx0nFMnX8ubtbdDWAi7L0lAPwbWeLh
Occae1U+qyVN4n389WUPth4ciEsdUXJVDHEn8Xv0c7GtzvvkrWh6fXXmBPPkBCYFguYyRjm/c+E6
+VgfQnVoQ1xmSY47yDzmkMzc5xvNJ9osK6oUpdxqXHrb71FcdLhesmXXrAgwCQKrhA9ihfYois67
iyWTkuTzPPZ5tggvdctiaZ1f6MmEcZXbk0AKH78BGo2soQqtolVfSnnDkXrSkpZhhSsdh8yvzARI
bTFHbabP4oMgHGXbE7oCPbJP7TXIXHAzS81yqCS2pxkr/aStTtQCtMlURNCwV/nmKbxgSbzwyVLd
S7lkuWTNWKpVEehx3IFdNT8MwKaBRTQIyubsviyadZHAUd+65nNQgTIkOPbt1GPHZZOCT6NebIuI
7wzNnMXn7NXT4QABLCwdFRL5vFCLtKY08MPO2qPxLmTMo9tyQfRTuFqFHumP+EVrF5sg8OrnOueo
PUyJzjRsXn1Je20NcoPblhmV3hWK1RjSckbhHHTVNFlAcIhSC2kbV4axstNfSNpYqbaPbVW2jJdO
3r9rCLppg/zp2jxRAX0W0tEedRp+3oeseBullN8ZhPKCF8j8AYfN2krkKFDcDloayJ5ZJWEFSFlL
YuHSrmHM4fC0cecIgG2m/RrmSxXODNlTPvsXXNmcxG9vy1wZS08QiLF+FBqlg+j40ShdAtOvwnUG
cq5SyuZXsKYusuTwSI7CdsMyQ8H9OivlJbzDrN7z6BDqAR/YQOX5A9wtY+JFeTzOWLYWkG5XMa/s
2Tu2QiFJGEz1zMEhln86GQi4XHoTLSePYG3v/EFfiXLnGZFpF5VrwpsgIULDBok8lpMVzMfRXpbO
FRm12na9JHiid8dlmYx960CU4W4ZijKXeGtZPJ6SQZTprAcF4d19jls2Q5+BQG9RRQtLoIdBZl/y
g/vhHdnBETJOAcaQ70vuWhCD/UMjoAx2ENuT09EXn/H4AKlMp+GqWKxxcqCGpabMCgsO8Po+0cmj
WIxufNI8TVb2hkWm5wmk8c4lUdjsw38bqswYvyin7hFCjCihAjWUbOc9t9c3cHkIhMaO9jfUOdRx
HSH6jG99VagqNBuIfgVm41s9Kj8or9kDWRBtfSUdNNMdoWqTzdERjGjWzFOFcsGRnwVWrspGBexD
3z0IgPhHqBWb7Q8jnWi8IzIVh/BAicekokn2tQF+IzC49zlkYVEaFvcD54vSkaG6lH/dDZ7ysI0m
uIyWcGmI0nhWcpzpNxqwi7eKEEieWDG21HlO66nZ/abNpjQ4rfL8+YRCr4WfOfo1+Dqm+EmSq3aQ
Fv0Mou1jGNye+1bT3tMEyBRHudNlOVCbkgUY/cf8XDyT73OAO70hCImXvLbKNBbLLcgUAnDzhemo
ODn4/7Bz6kOpOM7ZDdzMs6WOzrdSIdH36ba0gy+ihKbNZg4+Ybik+u4YryMwSe6KMwCzQ0u2LDLM
LttMjDZT7Zb1f1Yom0pTEZeFsjXxXfLz3ccezb1LVLYTo4dAK9esBa257IP77bdjVTntDtzccioT
Bpak1AttFoO8IOAexI1lw39dabQ0+NND1YRyPn94RzibttvkIKPMnSkG6XAIsuUalDYJypaFcGMh
ZApmOE2Z0gM0fQyv0zkkwknDfMJzmSj+RG/tRE92pbwrY+tFyT8itRW7+H2bV7bUzSdUo6n/cMhS
gAG9thF99YC6tLqy3U75HEasvBAjx0KC8LSv7W4NNSDVxarLvco5YhXa/tA2YaGOz6HagKkiUDLL
MAJUQUS/x8ax41ve/OYkMi6oD/Sc3I3EAbJArcQAPjYnc8Uj0uRIWKZyMvzvUJhhG/0MqB8u8Qix
XX0tlkatjp1hBgUtIyiiMoJhEdFJEuaP7lv/y5iOcIWzFGXSS1t1AitSPu2ZANebeGSzoXIbEF+a
sgfdpf10Rh/j5jJJxTqbA1DPC60o7nhsDKVeuUZAxntY9BdjhHaGl2i/EfQmjl/BwY/ZlYtnAITS
sqzcPNOE6sl/pQaAnEs+r0su3H7ro0N9gV57l4N+S/Yf9TqQUAjoe9x9OmAf8dWy9XxcRWH7vLQp
9GF6YQ+HJWVqYkEULe4ClNFjNKnHj8RI9sEekMvRPxbBznK7QthA13zWVK/L7ZSVlzmEy3lq2WfF
WYwOQdzHQAENqC0SpGNlpe7CaAu4uHm6YAsNZe6JxqWIB+14kjXrqjuWrmc84tiRfXcQwjgTR/wQ
gNjW44fk0v3AvXs1YYGA2ln6uuqDXhlLgujHOFyvLpwQg0FsbF94uMjCdcqzZ15WNZkfgETbyIUK
Yc5UViG+yO1mPotKPcd+3cRbRWrADiH+DIoqI49eo1WDLnTijSZ7hJq2Ll0ja04KIQWN/J/z3mk0
pCecZUZvDTxhb2lXy1UcJP0ZtcxxberekIClIZS+8YwwS5qApKu/WES9czOL0elW+oBeI3kKnh8h
8bZnXWeH58VUCE8oSxKzP151jQJ70dAE4uKosEgs7qBQRCb+nlWokhj/RpKeOWaT86i0p2iq5oJF
nOcf+hrtkgFXAjiixVP72vwUUNZpsug18IZDKIB57qJ27bOCxdnlcHrT3Yr5T1PmQ45RBM97afbe
wOpLF7GpCo8+abBswYLcQwE1hXmHP/7nSFp7YhoR77hfyBroDm83hkjw1ecSbDVve83062yPVTrJ
RQHGc6slTz2+gUQ9VqXOhPfbzy4xF41PmV7RBF9BGA/nn7Lv6Ual73jRsm6z42kquZX5LmygQZ1w
QrBUxgY7pfQn4lKgPUE3tMKmv4r1y5YDpPGwXKG7A8bKan6wzQn/Jhrqt6a2eB0vChNczGwaoh94
NYlQPTJnzVoYNaPK4H7hGFFNZuX8yW9acHhBe/08oZfqi8M3TuR7GwDqbRcLWigSXeC6dKoKM/FP
WSfFF2grCC5u7s14jvAoEe6hAlPiOL3+RSEk0PdPSnswUULgpwIHkhdb3RVVTiwLZ9KZWG2PG2Ux
u3VyJR4yhc07lRaJO/ig9+Py0H7Z1kuFVoLXQCqqImD1+dwqhHBqG45TR+yujMA00VQ3QBhaykHU
hANJghA8GDXPbqfpNnEOjEwr8HnKE335lDCDyJXeMprUHgzKwk5V1QgFPGGtWM5w0N0NMpO0U0g/
aZULeM/OOnoVu86uQkulC2DsV6wWsnLTi5hHroC2FshwhjTNbd+6/nVPSQ/zMxarx3kep1GWWI9B
DLLt+c/jh+Ge2P13/Av2qrajGW9ho8saXz6rS+OKV3Yf50lDzbFYF5qXCNN4wzcSShUtPBSXw7Dy
cnfSkruA2lbt08T7/0FtYBJ6H12sgV1tpUPwiJgoK7EnGUKJJFZxIvt+J9kXxVXGazRjmoyPI1dI
2WHDxj29wjLWr9aEmV/jRWi0jS+tOYgTjuaypWIUlbJJVZh7cd4Y5rKlNLOLLzeGDdJ8KTf0aWVC
on3VfE4SYh34++mx3t9285gu+psP+l9bcPlg1PqzXdhzf/U5n8f8COjS4JqJ0WlCHXBx3XXq34Zp
A1Lvr/K7t5WBHN5MJTqczEqjA5esbQhClWVZZBq2QxAkTfWXxwpehKg7+Oqh4aw1WbWzuYAbSGFG
ArXXCzCYbn9mBnQmTcz3JmvvV5zLN8T4iE+evZNxK36fucASAPw709gYJq7xjlv+vKlsv0S9sUiY
QcFWFWEk2L81XmWGvkSPONbzTVaYR/bOsLWS1TOc3v0Ks1mCFjwfCkFxhC8SzUxjj4hsZ6X2pcxr
GTYCZuvV+Yg1Ozb4efILkMLKdnLGWdxAxnrQGAQl4UwjU1gtEkfAso7nVFabjHr+fTw7RGdqj0TC
pAXELPgKmThehUWzd3KBMWIy6rbPy016dPpzXawq2oEJ/dqWUSTw62bnNTcJXT0/MfyaP/5ErLTq
QHllNIIn6jLhYgxI+qr3HLLxiLAzbGou2WheMwxD0NLIk7JmdVItwdz8F8MIOC59EqoTVSYKBl+H
JVihZoWtSQYpW5xLAxrsxQoGbHpxuD0lBthjrZDoXoa5WU7QeAWykTBOEUq6Us9esKKgXBn23SCv
J1IMMXOGba885dy7ymGPKZKLLf8Y+qpmDL5ff/XyaLgGLGMF5MGGtH/fXebEKVTrOiOIyL1zz1IY
BfgwyZNTb162dqGmxM0mOvn+ivbcqZak4GG+4slSpwwvP+GswIf/NKukZH47t0VKe9hrSocaKpEf
UiKmF3dOks1LxNdjrxQkNv9wmunaQD9kbfkXx1ZUHoUJkydktPe1e5osCcdvP9JBEo4I3W5dyTul
ERIKAnJBkYaDdYTVHbnY3SUPIiH3kTdvj0j64mGeUAzRpMtr/qX8Kw4IYWACjJUN0ifIamsmMCx3
U+S5+oc8B83q4ThDyqGS7D3bBexeJeLlpP/r3wf2hCnscbJE8WBOLTPkMFqoTzBUKyOd5qWWJxgc
S+PmQh/gLB4njD0CWy5K/WFkFg0XTBjPGayf/30nyDy23ITWcYz2Tb1Kk3RHcFNo6T1P4VzEqORp
GNv4eMUkX2nCSFxyf00Hc/x52lQ226+7YxSvbP8pJkRbs3q3tcN+rztVu5DaTW0dVWvJu46hsvh9
1qtGixhX8b27DVUvAWxlCBDah0fcHRnP0REXDExvCn9iy6fHzsJIJWp6OsVTeqMYjasl5R2smLxl
wKiidwaVmgyJA/awY2jhk1ivYQSW5U9BCDib9kTcApI2cOrt0XIPb0YMSbVP/fx1u/Kv6CKit/U5
UjKNuGnO3LKFp8F86BLSIlaooqUjsNwup+ZtOcNclJcUehtdvWkyWP/ZAKnWHeH+OWwmB8sEgMeV
12867SxHYq7wyyAqdrI2KorzW1ulqKe/Uipu2Z9XWc8KWBRWkgKFhdvuLiZkVA3ekFRrSrKqP0Qq
NxDbJyWzkHWlnPHmi2u9+eEyMObeI/aGQb4SclUh64iutnow0b9Yd5QVfBPgvGgd3IEAMWhvtRoY
ZqfBFsgx+1dxDQ1Xl7J7J/daRj3tx7sghdfhAnInIGzYeT2TaIebdEML2xEeYhpI37GphdI0yYcg
h9g2jiC0PtupKF7gmMPZfCDK0VRRmSTY7k83U2CrI0sarmKa9jIx8xWY5FAw02VGTldavTX4RXcI
IMFpXlrGwqtDLyrZrKrVp364arnvM74hN/mM0LmoA1yGFzc3K/9nS7KIZe3EDX/05U10aV8EDbIR
RSGG+bOMvQot/xXJWuogSxQeKiu7WkqixBenlsldXDssDa3NJpoPqInewQ4OFi26MU28epxiCa5O
tn+OxS5aeUtYh/gXVEVXjoy2JZboSAugh+Rp77BVySoi/uFrco5W11k6h5NAEZAh0mixrrI1l9Pg
vv3nriWa5akzjln30MwqUsFUsrIpAvPRFZfBlaUcV5i3sUtPReY6TxusE9owZ+s+9jgO596RTmre
gHlAFUWY0IJ+mL35i6GFWSmPreu67XWuBfX0rQTEN4Z5YgoojqGbxdO+urQT8B3/b8Nh0bquFm8/
ySsV/OtSzxX2vF1s15PTKxjeUi9wrlOXf4DabYdxsU6E9afleeWrNRtRA02CL9kW8krULnUBtElh
9l4S9p9jY6/sVLNu6OdEXKJcffE+ljhRXL4OAqBhfUjwGaEoQhV8R7rspBK+wwXStxtGLIdgYJAc
BuFFu/FwOFJDOBDxo6d7MCW2MhOryfPDcghrfOUfvdKw7p4hyna7fAVYwnEp/wqtTm6LG6GSdauP
/SpWAyDaEjZjGjWRvNawHHuuzsGdkOtXKvGCCFjYlaOkLBGlYLS0PDmQLXO1IZl80sZwOWPAxIRa
n0QaPSLhpwvHAMG5s93DGQnmyYfPCW03CPxqjEsmiG4skpu6oPOnwW3JXDdPVtAc/VQcole/nbs8
hO6jaQIFSqvHEIg96ooQYTOx+o9j18D4Cawj29yDBJkNSpLZaEJ+9Pvp+E6Ca4x0XZz8l7923FIu
1t2+cB9E1HGx6uL9hEvEqru5e1LXY4KiDFi86dP3FwOtOEqIbQzkvfdL1sGyz7+x9bN73zP82L6v
KwF+f2PFOIPBhdmGkUxiTszm0dYETDNrxIFYxoNq0StyJqWVBeZtG833qrsGY3eH3svcZq60neHG
4/nwarNs//q7bxXPZhnt7m05q4dhV2YEF+DoptVpe/LY58OKoOMQRT+Q16pdeHIe587JOXsJutC/
XqFTLRjCoK+vOjtux+W06bnr9VHQFWCQm1o8qPtNhN4bdnI+f/q8nq3hso0W86pp8N1TLXtEqiPO
Vmihe8y9RXM4V4Hu6PtLpREGGlNVZpDa/+gmmFNh29YykGhJxwIkK4zLLPsXXVekB73VRO1f7+F5
aNCz+XpgZ+MVYyuMpN/7VoalAXdDMBmOvn+UK4KEpd8tAak+bw4T1Z6Lp0/R/hKA2Fl0H0eHk6WF
7Bne2Wi9sNpjB8KkJwJh2bHLYedzxW/ZpLIv/hZPWlj/Sh3rPORxfhaCLX2ogazebFs8H9lWnOMh
YhD36llcFO4FlEJey4oAIdJc12eanyLagrbeUOO0WB3MrYMsCWekDyEvJKWiB9xBv/kMLFYP9gep
ynNYDRtTuj1U2gjhA/u7w/kAdpK7lwGJoJT+c+0a0wQH+xdhQKl9P5V4dlPNBaQYhGtEXkv931Yo
g+M9Lhw3rpKlgNTKqHLPse/WfL+yHBKNE5GQOk3qK2KFOMUq+syLfRJTCnYEb2qiDx2PwsV/0GZs
Y2/YPqP+nbhf3YHFYHyB/l+1hGERZ/LNW6jrPqZiO6zQgTAyEh+PxURMC+gbLhsguUCH86ga76br
CV/okHIEqSktpdh3/YnDuLmPvEmzi7sVfR2z8+bIckKRf6A0NnULCnQU3wN4bhsHc+/35l2Bmjgw
3U0lMnZ+5aJth82KFFRGCfiD0K/0cTg+6uJohGSwSGFeJylNJe4KsiJGQLZnLHcQackhjcXDac7o
VMm08MPGPWfiHSa9sU+AFgIHpzO2UsiDzxDovm0c1Bs9iHdd7SitqQwronFzSyQeuz3O1fTJfzvu
spar2LL8F3kr3ilYvwy5r0eTLflxRIVHRiYI7LQNyE13oUn2Fe1Tl5wsqia4fGRGG8cb+7pqtz06
Ns6/DODl/Gkoj1rS/aNk6TQpPV74VIg9imhyCVaXogq2YqACoxnzSZP24cllW+makteBM9KRyZDm
fW09BKGVK9EqMIzu06YSpysDOrvFDueSKiCqjUPM9cjmU6roEogIu08l/DxDT2V0gfhF1EBQsNqs
6CIz+Wdljih9HiM3SVB5sdBLZg5oiHJjofRCiCIykRhSdHbNdlaVqp05cm/hRPi1SSEnzd4gr2xK
QkLInc+FgVCX1COwl04didud5NpCJEyrMXVYFCG7UzyWtxdX6otWBVZlvu0NCrUV5vliaXhef/C8
lsGHAmL8CoHDyvhT77FydAtFH/ubTm2e5Q7XDxVufjmBpABaB3Vvk1HU7gHC5rtu8JdxTz4mxPNR
4AoHLgS+vWYVY0Iis5ZaTmXM57KFABw9heAt9aE2MSxDyh685Yb86/lZg+d5vZpDtH31Rn1ZPFUm
t3CIBrnZpeyDG7B+3926HLfDRh2Dh0EC6ZYACSvyWl4lkYPZzsCosaDX0M4CNESXYPtGw/u0npTG
R75E712yzegDN7YLvdftK6/BhfeX13FppWwWjvIpcxZpPVzhLOTBC8aFIbw98wPgitYIh+UGSUP9
Jp5ozUBsZax+L6zLIPtCVBV1F1hcXa7xfMyj1i/wz+yysvld40SQCcqmDMqC6TZNG529Yj8qAkLt
pQzE9RVZ7Tgx/kci8nvEdzfYKM8Q6APMPeYYTQaSe6rqc4nDmGUNkiurkYZ5Z4OO4Fun6N1bIbaP
+3hsUlzRrb9RZ4T96s390WKd+57x3Pd8Um7AnMIljL3DRUyi0EFxvW8kDHJiHs89SOAEHidJPflA
235AvWBdKbTiBdwMYuWKEDphcc6OMpu3wqRqbGxHrUl3BsCvRL/DQhvacXVEp1xgsC75/p46i6Kx
tkJ+1YRef98N7+AAed7PEtd1MW/c8oJZgjedvFSfGB136Og5w4X3TflMq3Iw177athHv6rAEbyZ9
gWHsHculcRMSHJ63mJjfT/vs7xTX8DrwrGWM+YIJVZVYPLM7DkJryuDDFIFtnkogL9hTlbTcwKNh
0ovdzned4thjrxAMBs2AEiqFTQbN6SxXhDbFOR1gFNrVhJkeMggFmGzfZDMTpHzmiWQsqmONWLKP
TM7uBKSl74KiMLHM85E+Qut6qvu/jGx/HUuB8/StDFfPiwCCIDT4psLotDrORAz1sqhtJOghdqNq
PaOcDoQO07pZn+BhiTbZjVpaYZHPh27ymkoYFdsSA2wAWwjQ8IM1G+UD+EU4xM6ncTeLSxndqDxG
JF882Rk0MRmuEe+FhysIPe+LbGMccOiEzALQApsJhz3L2eyYJaG/ZEtQA9dFjUxRtg0RXX3PskHQ
6QM4el77XQybdKaogwJyFkUrfbIO+wqvAegkZ5cM29twgHL612yNTBPmllFjXpJd3nau5WoO1T2B
9YY/CKK5GChmdA0Ckb9fgiy1lKXDFDbBo1slgz3WSxaJaA5uDcMPDA8ToD11VrafLRTlcQCqCJsP
tDMwBB9wt9ApCQXgh3Fu+z49i1ukuYkjuZtUVOT2s23QbLa3EMEbBwmtAdZSYqgtvI06Ton+7mRB
ApftNltYm9AZeQfTczrYUU2CW5In2tp6Nd79mJfMKnUfCWVaq70l65gCiuPKidscA6LAu4K0s5yx
vWIxccWSdWxSo672giK+jmWT/kii19vJ1k4e+roao1+Ux6kHRynBN+QKJGsMfYO/W/3tFTK3NTBT
rol2CovIAkiRgh6eV3lP3CeC/3MuSbe21oTok2wHLx6gGdCxvE/wZpTKXwdZDXVg2xHXMVfeKFWE
3EywrzqogozTb5wHfIdxDnGprjl//XmxZ6sK0OjhDharjjMJzYKip2MSghhcqAQxAc/YMwvMCZR0
QInJjjGWdahOOKvUDInyDXaNpSARV74vr1vqUt+F4e9FcJZwF5nZkancPmD3qioLV+1eKijFt/mI
UQ3QHuPEOLgnnMjmJVaqvlVXGl0uHGGue3joFtpeM15Da9zB2RtZSIGICt05Pg4MsB2L0MQBctNG
BWhY5uH+AEP9I+GjxyZD3gQr0r+y/a3qRRDXiqxwJk1p7HhNQIGffJp02vBisQ3qqr5QXMuFT2R9
QwTUS0GSeg/wCqUPKy0NRnAhpFjyPYr8IgFxOTOS7FchJfbGpWXAAbqcrlCGWDEwIracdbejIiOe
JyvaZ6enVpTUWZYYBq9c9wRnyIhQ16PmvQ13uScAf7eUX4Wsr4yYcB88tL7rPrzRyb/ZEvOrwc1y
jUPU3JpMGiIKFUiHWpPd4SJz78Am5MzjKBjaO29ICwIN7guUAgvFjno2IP8PN6MwJLcy8wlu64ou
RCy3HDkCK6Cv7WHU1TlvztEIVyZ/mjCNnZ6xR2H2stkSZXs+CdkdR0IkYp6Io6TwHKCGmC2XSIs2
bPU6iyZEv1x3rP+MIXQYLcgfv2xfGw/9PcT2u5krko26YkXplZc5t1ksNHedlcZO1qIOmmGt7SKS
hbaIFeIcGGv+Cc5vM4dWzvfU2GUXNN0gRtl4DJST2uUagi9GR9naiM/Y6+myps8dwtEysL1XIFXn
gSWPtiTaUfutc8NERy0JENX3jx2+DS0GwEB1LriaAJMuEHmIZZxg0sshQ1YIuMavLWT0V59OK6k/
AsE4tNqbE+LvRC+vmCLu9PF/cBzCtAGQGcfA4i+3R//FbYLPVZZ7qm8w/oU+pYZ/qED/qtTK3NWe
DZ3gY0bJVPJ9lSlyU96r/ZgKsHIuDdd9aUSf7BYPFNBQeEk86BQXQ6W4WMgUyN/fh6KchG8eY1v2
3oTzkzcf8grlsLcbTkTQ27utu5wkCu+KbYRD017x1I2XUHZMpc4ji5o6rixWzX/2Zj4KvpNXLihc
wfOhtkY60Qy4sWPnTO0HdHI1EBuf1O4LjRcdcrozIhptYhOVz4y5LeONRrw6knrR9Ygvy8PYAOhQ
vWcLvBHvrveoKRYw1RTXjtgxUiLJjhSIKXhTVIGFb70ApbFQpvg11stEZdTRwFxo1YOULI3gdkqG
jt5n+OXjiAiISmBwUYQzOVi4C+9wMDD5BRU8tMF3iKFqEX2GxH9Itfo3PQVBWDc5TvTm6qvheSLr
CKRhgi/YA3iXP+sV6DqJuD1bmN/uPRyOfWxpgqblMwGkTEL1SV/yXoqvmP5T76rUUm/1L34zKLA4
ye72bACCHCuhrv24DYgJS4PLHH4YQN458n9KFBbTD5mjJcKkbjPNpK8cz2pnWyKeP63UeH1pAIgx
JNIPyLtG5sOeDMMasIi6ZvEExtccFEPfw1CqSo85dR6VviymTZW9QDvT5qxIlj3DMKZJUMmt0eWf
29f7WNHiMtzrJZrneMciVOPqndx+3Pv84Tj6SC35hm3wcwPCy4X1nLWhNXiKGKx5k4SZi5d3ChqC
7DL/Oy1lrBbWfEZnvBroZjxgYcV62W+55dytOU8Dq/A/O0UcM9ZqobhVMSxKzfApoX0jsa9tL8jO
W05ytB0SrQAGzZsT01sdAiQidnIt9Im/fYihqXrhMHf7RVE/VclC50iu940Y27gkYy7tZLpt7PSV
AkwAnvCdl7+LUQrm7pCRJzQ/uRqnUAVypQVMhh7zbI8Kiwv4B9pCnOY5ADZrN5CP21/b3B2DSJym
4B5p3MAfIn6f64YSkQSwRA+Fd9Ihj7giV8fIK0XodMZzugTBBNZ7K2FJZYCPhQDrOxYsCqOnsZ9K
3jxxBUA+dD9oUFZaGg2toAw/gDT6jMNm4WSU+lTFvkDYdIh4t0qEUnDMk+tWmKDpARewOWGL+DbC
O5TmsZfuur6NmnHLBnigae29xqZ5Aa+UA8TbpYfcr4uu2dgSIgiU+j3R/bKiHZBBNuUxjHXKT2U3
GzHsvq/R+YFY4jHzL/iOQLBnr59QHbLGRQCOdSWX1wO2q0kBbaJSF7OCKmGc/UrCBJmOSlag3OUt
EOvuzHagy6RcmWtrvy2k8Q0sqYeW/EqV5sKf4hF+Od2UR4PXO7n4ermlg5F3XU0qk5JMf8bYzaoq
K/l4861H/kDkCmzbKRvbwOoKadwHcgK9Rv2yJedRq+HbotOwSsEsnv4PO8uFP8dt0I0XNLTW0aeK
m4TVdy3zJGUca7vkzVo74eXfSGpRuTRllNcw8V8h6KQhjMv0T9JRLSnCCqGZpS9sRlj5zA6nUJiN
3uHaRf93mpQonQy8JdXZb0AuqirwfmxWWvoWZPwDriBwvNSQICuUu9zjFEjFhFQRdJcPBt8Xi2vb
jySxIgsDCbHWr8tRwWeZlTmm0GZhk5XCF4bnmkfb+VDAoCUCLHcJKGVnqTx5/Ciw2UyamZgclxKR
iAMEC9B4P8Vv4eaF91walApiHH4X5QTvayblZ38mZP40AmEX/fiSWnimvUpQBPvzX1MB/eBfxliy
EqfIlDwEcWp2tnNa5bLQ7fUvma4cahb5xoREzGwEQEuN6jgJb0Bw5yssOxu1/ZM+eVpODfdaxIn9
q0W4BI18A499DskJytxqRW6WkpTD/dgj/UkdTMp8rig/oY/iuWfMA0thDxNMkaxkyxBitVdcJPAm
bY4297OH6VmT7XvgmBZe2JZU9AUkeKXhfJKLg7WuXfz13s3ch4Ru8U7yFY32Jk3E25Ac+AoRPmRi
qVDS6PbmBo22iglCVUa8prDGP4fPO7ihqbL8iEYKHo3SuLnkEL9KMmf/5RzANTEDnZHq8uaAcr+2
twO5Zycm+dietYNWwDcjnm4cyrusG1YeErH4kItE3SS+kuQnKcxZHQnN5oVIW/A+Hmj6AK1YqVMS
JllyIjUTUUQxUcAYrqCtrN75HkH0AdS41l8TyM60Qc3D+KQlbr1cCH+uM/ekOG8lscDZ/pXNbQlV
FGazpqitYdfG0LtZc9xLzDU2IIdFWWBRrHjv4aBcA+iGS2hUx3Cnc9UUoa16DraKZenxB4XPI5NV
LqSbZjMdZ7VkoTMSqNmdZohYsouxFVnXKZfOyRTDgC9nBVlMWv2R6fnMUTmk+yMBVHG8WRbSirux
A16XxNhSC8igFVowcElyGhH4uYZ14942dPorui1/ZRH2hN9ascK/u7Ozn7mHQIzll9JCUgWbt8y5
BulHxVOfMSbrtEp2JiIPyKefHcLZ5SYqCC3dX8AAnHQ48PQTQEQo3rpsnuoV5yT4wZX5fyDDBNiH
9f54Ig/wNKzMC/u3Y3D+U6Pnhwi5WSsEtfyB8RlSHdsVOrwvZJBKLiducg4lBa/q0cUxna9xZYq8
cnTn1+QpA5txd7LtBWeZivWjU62SdonZcd1cBGvEGo2Kp+5wREBan4FfyDWpB46wlACj4yL0Z82r
0eMvR79x5n9Pd9crSyCJA8+2eVDflxF98dh1F17Zqh0yqEb1+2K2eXOZJ9duJ45t1MnZixNiVnm4
a8Q9CeznVFqPSko2IkFIISOaioI4ERb1OiLL4UTB2CjVzSLVMO1oVAFZ6WXCvHSvl2ufvqL6/g2i
C2jkmaPAXEd+nzUGgrYK1zz3/pDChG1HG+Y3Lfe70P+FsA52ryEg+hjQ/86VcwSvcp182EjIKGFE
WmKgiiabqhzdDtFFitTrMYfH7KNgX49l0/jzaoSVzlzWj0+SioeBbSF7x5Ll2AuarF/GFcWSCkaE
q5OYnJxAGP7JAvwgF3NeghJfTeXfH4VmubvkfxI6IqFvZSedMetoCr5aOen3IOP0zqklKPqqGufZ
8g8V+WF4bUIrit4JA+K+o789roT23OTi11479VhElPQyKeHWJAHLf+7ahgVoR1Y/D8WtO8k+fr0U
2uS2ZHsbmWEB4mN/PW+eYK84Mt6bwv/w41fL145Y8y9jFtO16QNF0zLJtKGgbsMa4/m9R3EJZCDA
LZs9hft2SSB39dx7+NFFhfpRtk9R4cuAYWnqNI4C6mIFcwPI1HGk6MyeElrGDuebaxCG8eS+ohDK
d1U05Xy5hMMkTVlKXyN/EBgd3SwTTNZdKNZt/Tfh8mYpnGgOhNIJvADcMe5x4yAV1cS8VsORX5+c
jQU3dF82FKeniE74TxiyfK/avNPbizvHfBw3/T5Xzw2SYzlNguMXcPA411XTBj6d9ehXaDWNHm1a
T+Jj5PRjgHUQaSCKxjgyKwDnGM0rllxxkdyJX3RJUqod16++pmYDneZSQxmNTFo20ML/oJ+VIRdQ
R4ulz0gPCPhgj0oUAcUXfIJkU/qq9AbVC1E/iNZUJbTUMVOq1uhF9TyttGkDuRuiQ4iQCKQfVem0
SJE9wp6N0A/ZtEb+1XBiuqajSWuQL4fc0nG9xantuKv/nnKCXMrs43s1aJkg8ddXjNEnmItxxgHT
huKDL9O3sO8Ak1WtrJufVXA8p9zI46jsA8H5mhym94nlOS0ZMQG8FhWo31NwOTiJePyNV7plxZYu
DRbbpMX6r5XHtohWLSfeMj5AmOzvLbGNzCqKScNQhzaoqNQc47rubYh7ngFqmqNOmURliDDcjBna
9qTtOYqL8EpKcPDK5OjJ9ZyP7SofwsAZgYJZSqRWPXxDEevw8LHTV0uc5gSp9HkPRzeCiVrENT7C
JAIHYXbJ/9DEuCMfJGPJ76XaLNmpjUlU+CkfCJtQicIGLqV11+Fr7fBVpvJR1pI+yOmCuqYGvGv2
SggimRXvGP7p8j7fXkLcfdcql/l2TIsUCi0pXAka+a36g9tbXpSIU+J2LaZoeZqhcXuFtm0K41Dv
XMBU/8NmFhdqHLPF9yOKd5h+kVZIukBv0W8dRbnZZ9LDvOjMXUA7ZlTgqCgHn6Cqu/C1QQxWT2QX
Y4C3MWjNmf8UE+Bq5HhQzen8cI2RSieodJ/t0GRUmZkjOcf5hFFKxC6OvDf/6lB65YNQUkrUUU5M
s3c+Sv9EcubNXNn4jk+hNKlk00n97fiMkwI2EHkuEuUKWHVWpvKj0SlHv6OiQ/jicr20mo6uneBE
2EtOLGLTSH21knNRdPJsBmAdZ6JQlx4IJcCoa1DtgNbqBbCdx6Lw2Otrws0eb19PXLSZcrHOitRl
BG0ys19/OMTK46Yy/VOE1b/0g/gm4N4cVo5X1HQorN8nJGC4OzuYKedGnTD00FpV/Ye3LX9f5ply
QFA0drjsQparVZjRxLJRljSE60LiuIqeA/oHHczeNNAhUFLMsozaSCSDQl1Pr7fmIcd2nQB2YN3e
QZO2UZFICIoO3sR6dxp2nY/Jrti0+TrG+mcht7fiuvwsedSbMbTYYeM+WnrgoEOY8lj9MdqvRxPj
Bf2xXL1LkfAZS2Cn1oukoqwk7GKMko2SDPOzkHz4ko9d/1SigKckN5oF7o7s3IM/0ZyIh3Mgxszb
HUtNJEc4Wss6FTmOR7mkONhBQYTqmV2zGxy7PPpLC0w0wSpqg8ZkMZsCYana9+UKWlecobdB4d3S
r4K9A6iP6PaDJs9Eoa3zoUl9buKU1QOs+eYm8i3LZ9YRshjl6CgQPykHllbVw8724ZkKrUBIIueo
i1a3CwijAGKtHNTFGhCsu5tnJpT/FUsC5SjKZvTlmVCRRpsw2cK8zh+PT6efd3f/e21fyvLdLyzJ
2aD4cUy7uAgiYjjTYptSMgEpJyHn+BNHHkN7VJs3Y52LnCmEFndtZC5RjNH6XLMzNxwszlnVnrla
9+npdsfvshv0BDDN61gIlVC/RP1yi5d95dMQwsMVPEEnC9gMib6A2ciVVKZuAVNzO1W1fte041Gk
ZxVlk7hP7mvP2Vm0fbUo91hO+dSAwisd36YYtweEkVFULbMV+nI7XhyPU4eQT2Sp+StO9CZrdRlf
BROQBNZcehRflsTf/DQSrctKN3fpGnr/tn19zwVBTWQ/fPPHTfr4drPR/Yra6XdWJNKfAbzomw7M
UUsDmwciQp6/Tnj15AlZesRzwXbOr1HzqRgY696zAjuRMWkKXT2J5o+gEHahVaajTqpa3JMQvy/L
7H2TRA7YerggSnQccQUb1pA4JrwKCXIvDaJRMB+9fLPilHuJ5dpZxwEYvdjsPUnINf2BssJ9g073
BR4zjLWUkec/dhXAUR6u/WKJOYmM8Ujz2D3LlfaVOp8R0QanogX3T+8vhpyy3OinkGqPJuFWmcYR
Kfs8wv1rJOELIfMQs6VnAGlppcHtJn/ysagQCGG+UK7lE50W7JRLuqcLuT7Mf71LymaqQcAM97pq
e5ASvxDQf6jjlHt2kBROk0WUH7r7FeqyPs/T/dfcjWl83H3sotPap/Zv8dqLaHgnYHrGn36c0gWu
+8lfTOn4t+6SD4sfxOcThFzBhg1QQRK4v3pZZ0zkGX5Js6ztGreCMGBVMWsnZEAQ7kuMkZQXi0kM
oJJ6zD9B/rV4cS5lNMFmbI1v6nZhnfgr1D9CHbz5XmeioVaVYVglFw9eorLOcYheIfHqVw/Fsw57
FZArLkDwx5qx6i8lV4xkGHC1vAZro3lu4r6R0Fj/V6HFN5YDtf6rbdcDbt09jVdBmwX4sFeta9kJ
m951xXyKkhzojsZzfe+5GJRlPPZJnnMQkzSvdYYXapH1Frd6/u7Lbyl9I0QBOSvODcXCMVS7T9YZ
f3CZt2OQ1NsZ9tV2lBjANImsxM1XTaXWf76CtqCAkIKS2bU9f9KAurML9ISpyPTEe0KkFCEjU3ny
3f/cGEi+GBuGdbhoVEG16yJTvTLtMZ1YI5jiRGybOEgN6fHaoa/RSUjQHDoAxQpmfx80BHsLUGwn
kBPYF7uZfXIoIOVAIZp5TM7Te7/M9Z/aN+MOtLMBVE0CVbc0a8IU85XMWBgRO0w4c9z7iFO85CPR
5o6EDtVHwSmmrI8C37wehiQZ9uPAJYkorGcvQvIAC5c8Pep3XUMDYDua+y6cILBbTcFi05orqd9h
tzpVvz9BNryejtKvEUReFSR3g5hl87LgkEyCN7IA7ZzKoKYn2hf9LymUiR6C1Ua+jWv+KIRecuxR
XnJTlCYO07RVe1ENRohTqEaTHc6J4XlHcUEzLmcpySsKDweABWb5GeXoan3AfN65f8xbeTHBSfR7
tLLm5t6VCc0zpe0kK3oq99vbSfqEIzMBhtY3TRazo93O9BrkT7Ey/bpQuUpbA4RAEJCaD75toBSG
Gk2zH9ygiFkqzMD03lByFlH5E4lp/0PBlRdkwOdu+PtdeA4dSfLvGYWPd01CyRe6pkJMh7llV26r
Z4XWkCuP/KZOA86UV5Jo3KlkwaNFw/T/V5xcQXsx//UOjKnXh/Ui2l2qPZ0tQzDVlVJRAftZaBda
FhAcnak+GJvHhmZJDncaVssY90h0gohvwLfywGI10hSktr7vs2QM0Cmxr8j7EEobhL5bpk5wHJlb
Zklz6dbcOKaW4bkdG+ScYykV62MzRiGPi2QK/V0Z6xSHZDJMU2h+2XI0qv31tdIZLA3fin3yJbts
y0/8AJCE53nLCc4eTBicQpncgl9bEBaBxw9jKYoi3pJELrnSd5JlUST/D6d9C9Hez/4+tDn2zBuU
tBiDTiW2B6QycAgmp7qgYGkIxG+IhkDDG7VBWqBqS7DPn2KeMU74CpQIV62v/99SDEZxpSuO2TTY
CuKHFpxQScWpIwW4EMQ6fSAZkbNyg55UyNn6S4VAz+C9QZUdCfdkufsUHnW5LnyRM15N7LgRykUc
ZkLRcEjIcGW5XWFhtzdy2NHG3xaitftxv2NuCCIsCbKEy+zWeUz2u+fhfM//plm8rkKrF5faAnaV
ZJdFVCDZrbXbmDMy1d2qJMTuHIZ4URoHC0tsrviffWli/rpUJJIjNE8YgS2UtMRR6nu0zuJ6JQhj
z9A6xMfjjIwTRBatLsZ8UgEzaauJ/8Nw4g99B3Iq+WDDWq8/GxjnobKHyTFjHJrYJ3uf2eJAF7IW
exxoH3Pa3C80zQwDyMvUUdwLiTfWInuwJhv4UZhLw8GYEa4DzYrvyCdZGywxbb8BdTy/pIotPCeG
ec7noUqx3Sjfnrq/qcC4NGu13Bh4TZiZGBTDdevlaiPgB8wSIkee6oclKgOy2pqvQzRHZloehY87
3IzttaJ9gwWV5I2KcyPmBgFWvO3RrZCGOfvW2/M2ZCTSq15G+8F9MpkkoRm38QG4NYLwvRaKSVYe
WtwH7yX4rGM/M5ZPuG6GJ6Is8rRjxACaSj2yZY3YFsXeu3vSSfmC3ZLbwIo7YPadwfCmmYC+RUF8
6QtK7ZHoOXOZcfA+Y/LgIelPgqHnCsMwjASZKr6qmkOx1hhKsOxpZawYkX5P0pOBKqfnrgPY8SIj
hJlELD35Yy2JjlWieIZfcP4RiULCwgDv6xvhMPKBZeNv/g09hiQltp9AsEGMNOAh+gv001hS8p8P
ORHsXed5jjsfncXkRYxCoBBWLNnWi5uLUWAyH/fQHIIIJO0UL9boRN2NhIkdAoBE5PBfexDSmfbM
SDvebfT6XmxaR0astYLL3sOOwij5U2wB2KHW0OszB8aa+hutXUgjvGGiB5QD+mhqPBJtsa58OVne
v1aziXQ+4ANUp8M2PLXwXuWaT+JquOqs9RS010Ft/Bh5gZr4hg7YrT62IzQYq1ITwSAMQ6Iremg2
AIB4fcHFIXkzCwMhYyP2U/L0b3CNqLvZMu1+6onG22m8ZmOlkphR2Pv99KuH0Sk+JTAxMlAWmi/P
pzTzJl5l+uyd3QC8ILkzq5WSnLGL8ZYcp49WjcSQH3lCMSyzbo8Fpf3Tx5cP6my2qYgjoV4oj5Zu
RYdzHlOIHf7Gnnmgu6165CBvYkrpFCPIBU4Dnx4Z2SZP2xGfAIuQaCtmu/nrVwXkHTlKl0B6GRZO
UyxX+WIgZ6aez4ouR8gF0EntZw/qFbtv27w59zdJzsqByeo6FpOwpFa/GEd9ZVGxvzoIyEHjdgVu
DHeuo1yq8HAcSRvFs1eT0lxKYze0KcidcRS1BtduFR+5tg/8kq15RANd26pdisZtzCVSgmQjx7Tb
CiHxiobXcqu7AM4yatBM4dHXkXt9rnSQxsGnyNET72oSRdaEdm+lNASzyWVUW4pj5Exok8IAdlz5
gTJfQJx6F6rR+xCxHm9CoSq2bnapBFfjuVZsUXrYNyIVX2UR/oAdvs4vp2wq9abvKzeMkv6iqsPV
067VeshHt8pKqfcISeSYAyW17YXKhXgSxJiYlhuqaaWWWNSRvX0ZaKn8L7eLSNkFREbRMlGF4xsi
0uYjKBeTzbMV79VnYtlIkS3Cxa6KgTDGkUEFQ87if1EJaoOPBdiYKhU4mc70cdIrDfUt64NHpu5i
hR2SQhS9qdD9fOg/Pc2SHEErFZIE7bJR4iiCRSoqPz6r9qTK5h8yHt4vQG2KZnfu37IXhbKxh0Zj
tb6uWJhXumlXSf7Mpm52zDdiK2MqAXXtPoFJbGJ/tVbtV1ud4/5o5sdcgXDQQwfAVPRz8kbOjO30
xITfJ+IfnsYZB4/974kJ9ienFs0b1cKvdNAJUjyGsEcLwp2sPlHo84C1JRDrqfWM+qPuewtrYLUr
MmRin2562DBogQuxWc2L27risJ8yYLYK5yLe1xhb/kjq1zjJI4rWm8a0aZgGVcznK9reqh5gIsbW
gyGjRo0D69+DFp2Ze8YEfVnflvT08w77NFPRzsfMUpCdsbOPvqLGCBkizbwSjcZxAhA/s4VyJ7V8
sNjC1n5WOtuhYFqeLzkAUgW1ZZeBfmDvysy4sIUjUMUHpIcnC1Y/23qlEGYBpCFqPGdNAWLfnn0e
YhTw3VbOxhK4I5t9ISlTiwARKcOoPlr2wlL0HgoIlvQqgiCAD3nkrLWaOTNTRiR9TDeyynzCn/JW
Xwu1qwKzgxTGbb1JrOYwxAz9CoSKGdOjcIY10Lo6FGBarogUt5OULPsJ+HN4++/dKlZ8D4vqXsdv
s8wA2pHemfJ7i3KwCwYJea2rHtnio0KxlpGWfEImUCX4zUSXkVCek33dkJwVpV7YsZI0nXaauDNg
eDHSJfQMzLB7A88fd/eDKLs4U3bVaJNyzQ/AcLMsel28xnVu7l64KzxNl0fPU5EvYb0cc05283VW
FLLJNXgRa61BtSgcI0IjzvUP84l6h0M/VTat0IQvcgvAaMcOTvx3VS2lgndtwbBDY3cwlElbKR0y
s7iTmqlzn/5Ua7c7zCsDHaxh+WZskuDJGF/pIirkLXBrMXM0U36xwR6FZRFl4VMKurDc8Zi6fpKn
tV8v4BUGKZChlaqljA2cQ/kl2EyYoqYU5xv44toq5udcr77PF0HCLQQPKJo8Lfzkcm/g1ycKVFTF
dGFrfKx3XJxIayK263WbgiAO2QGf0MsS34hI1ZLcYygaf0YoCRTaNiy0QFOfE8WRpOutF7wfqNd3
Dtd9XkCi9l1IZrctiNlaKtvzebzFrAuIva7BrzRx2GqpGt99hZ5U4LYvkal0wKsXj+WYqm21ZDY5
9brHjrNw81yNBezDHn0YT5607Bq8aQTYJ5Nc77KaQQpHBwJNTlEqLaRX5L2Dpzy9ku2C814g6Qxj
mNjiBSXptAZh5ULv9OH34+rkp3va2xAEjmmw9Z90x/AI+YEwnPhaTYH8yvVY5p/nNmaQHKAokDd7
U7pqhtQTH8mru0FKgWadYPvmhMyMWPATgf1w8zUTF5W1JWRwumqMgsqMeiUcFeTE7d/LP+DjNZIA
W2y3Vfk3r7IpKNFXkXEPJKK6kLuqTZk/p9yYFdDP9goFhIa9fRpQGFO05208pqI9sKHoibf4RcJ0
5ZzkOmc0CAO70ti8PzZm0TUMsWH7V9UMWEUwJlGtAJlBW95WoyJgRs5MKqrjWRhkt7LUjLvGzARd
RJBmcoFv1F7Dly3+q3afYYWi6JlBEmAS1thSVMm8MM3W/Od8djV51C15g+D5sAVUfP9h6itOhicj
XkyCLWh8MZjok2eMbDMwGPZhOllw19JiHr747mPLSQdex+Nbts7vhVCOW9JPIY2lgX58uNiuX6c/
X5VZlq5ZcV/35OAylMSiAKNi2Xl1g3Hm2MLHSZYqxYlA+V5gkCLYmcPLQIg+Q8EE5CoEffMbI+Ml
Nm+Q2Ex7Oxqyg6NtV86bEw6+88tlR8vkpVspsPq9ZdRinhOnFz5KOgYnS1Q3weycJJFi0TlSmw1w
pAq1Fn487CQn5rjZ/GVqgqD6X64TbasjgdzHCOBn5gy4ZaNOm/59ZGc4mQm44DyedPYERswLXWHc
45LRW16rlhLNngGjhUgwSc+ITD00W448Y8sfjYZ4EJBk2FMvCqQnr6ejiO9T6XgDZ2LxJZTbYfLx
xbx3ZtcUQu0u+hCEeXWX9IKH1OOnIZUTQPgilDJeVMbaEPZ7yHknPb4xZYl3wOlBdDM0a9Uyvv3Z
vyZrC4w1FL4fQE0zhcLx7kuPNe+NXFMLLTkdgUzHgvFDWWkrXr3y22jyq+1dEJ72W/XvbI3O8n3F
PBIDBTP+Vk/hNSIfxUDpLzS1ZhJEODnEtZc+oFf9mtUvlBsWHEpaMV5+i/k2yyvzge7zgv8CfKGw
n5wWLs4Up/+i/uzzIJcuUk1cKzKise0MM/qxrjNCOXrHLAweA1Dlb7jNXIsTb4YE/+iIssOq2ory
QoK/OJR0mzQkNH9rlVkGZmjB/R4c49kisey1LJbx1oQuvU9YVXCsCm4nqJVUBgb0T1yDoNBm7tpR
sK5tc6fnqamxDDTnvfobL/RYVSWRlCNr7t5jG0Vuf+3Gst3q6SqoP4Nsm/b+E9ub7BNyTxSupO1t
NCoKsYj/K9R1gdTIq1l8r+kEBzzp2BGLsAG+c7Nrnyh3u1ua3cywEvTdeWIVAfMhbOHAG5rc4hFk
sGBYYOFfRTaj+NnOS9SDMg98AgmxzsSxCw69bhidEw6VbseUn/wDn0ryn/uyE8WnZGA41OLMUccv
D5sA4qJwBExBp2XVa2y14R1mGAxQzOYcVOdnvln09BQHDyc5vbgFSDojiCInevdJg4eoh0P2iNcW
KyfYsmQR8DPeuJPfJ7lT26cuV1lhv1N/AZ+dk+GCMrCGXaMw0V5/6C4QsVFmBqsL4RrvsiXn15MO
2acFEyu52spNIb8S5BHxvwNLLAmGsNYWzy2ohEhW9nK2fTZMKAy5GwLQp51zusZf0dutmzvr7X4y
NgEbx+cfg/tl3Eci9YkWhmo61felrYWZQqtLmB4R//hffxX3GOslvBIZFhiqY4w8C1PqCL2daIpL
PWewJSqZvwjX+gkyzvDlfPvFAToJRm+ZwZqWahLt3F3kLlsjwBsxeraExITRKcZWnDP6WNJs3W38
be3oaxXgVk4RhyrPYd8INpiGUl6oRIhlyGwRVADTzZoFieXGi6NIO90pqE7vCw6ZXKNh9TYQS+Ak
rj0KddsNi19urpD1y9wb2vPxyI9a+6aMDNRMj3MogLlGUbL490FBFhPWq5H1t0mlhC0/cqOlJ0H1
aLxKgZHjOOCQo4qhlBWfzTq6VOEnaU60LIOXuLJ+vEzAHtx/aG4VV/O2Q8XqTu0PsDXFwfL2SSJb
Vg48P00haGiRQFvWBYm+Fcpx9uhgmZVgE/6NBlIw09Ai6GuZUXkU7OnEhyh/oqqd6u9eA+qAMcM1
Qwd3sYI1L+9O0N5i3au033CG4aC3mkMrItquwKRlUnUjmDzLgDhM0423MujVO6UDfUa0iy79+bx5
HRd4qWiPcwUPRovePtrtTpE3QEGpaI7GSvajJ6eISBdFkIRGLBoV+a81odIq+SrqysDL0OVsDq6m
6ElnoliFpgVjSkwjSSpdrCWtXleUMa2EJbkAikDWAOzqQgmyJKb8AqHM3+57Fe+BUq0n9OdumVCM
fXNwUALM7wuoDgDMb7akomnF9PupAxlDHqnvk2vX7nIKR7Ume70jw9kKf3+Z8ofWBNd2O5AOk8YQ
b1vFu4UPYPVJ0qxUNjmGtGExIjCD9mbUWBmT3xZkG3ZHbjYX1r9fT/nMstXc07xzAvdbp6ivkbYM
SwtyMrYgUh730xZztQ+KoYaKFrGOf66OGeruouCToZBuRT1bU9mlWk0tFOiFNNtg6q3jNqs+/v2q
lKFSGjMJVO0cLtvZ6y77p/46PPz4itWIyTEJ8CIHm9/F38y6Cpky0N8+bOD9Ha0w1wEr/SBLGKt6
g8+OrgSM2EsNDU+YeenmrED1fGrscZoRwJw5VfOWhNNSj3rAyxAWgq0vfkAk5C4kmGkGdZhPFaV3
SjZcP/2c+uq1KjOY63RIguAcY8eES2dMApadhFd6VoI8Hz8K1B7jM3tcAuti7pCK6LQUSuACHWic
LJfXRCDR61awoi0nbPbyLJvoUdUX/ECnlRK8PGx8VQdHCx/2K2T9rEKH1S6ytknV89s9ofOWFVfA
Kd2gssfdTWun8yH+3+405Len2qRtZbptKZV6Z5V99U4aGjs21ew4VoQY7Y2I1IkkCx3sdMY6cZS3
jBO+0nX6a4IDAzuY0PAk5W3HRbloZjXlJqDLqIKa0r3sNmXB0U+GD2DExVagPdusFr+OPcbvGVOe
O7nettAXUXSMV5XTucv3D/o5314m3QGarSLl9nbtUGkzsHPer8RkH3WcCeEVM2W49NpYWcE9Hirw
KpvsNjKnk9nUisFgxdRwdYMgw11GB1EJ1jcef1L+myovgp19fQLfCfJ1XnRNQC0k4N9O79w/to+A
cYZkq87DjIez9jUmOutiN/eXfIliveGbJvOQliMayY4Qovis9UDflYkJC7APcKfwBULaYivF+xYT
XTiYhDxKRW8FVlIyJy94LPY1hogpoJ5tZVpZFiK67/5Y/SIwWv6xbnFQ/dFZ/UVkoW934l48koL2
xu4eJFkNpWl4NpJ0gP8/SzdFkE+CLqhHhkgc19cAEsaOQfgbHqNGvd1OIiHl8BKX624UVxVRbNCj
5imVEVe0tzNF5d2u9DZc5i7SEgQH6qJy6noj3aZUg4D/l9yZ5sB7v7a0N1nMtSSZleMFpw5TVi46
XPJszTui92yUf68WNTg4pNGu8Jb6JRFKUyjZPvtxnETxbotcZZxeURT2bm9nj/msJb+XtiJ7KwBu
8eF44KwM7HdUMsHtE91attumVFW3UquSCgIr3bgOPU5ZQheH7IEmI+50lUNzDmujd02GQ3Yj6SC3
TWhD7/Qqr0xfYeoAH5lU7qkmuZDBUP6h/kFA5VWeg3cyrrDxTnzR7h77sbfOIbI/lMDI567rDoCP
OCOL+x20ZNTNQvJPYaxlnZihuSjZGFNtqLUUJGI5Q0g11e98gZdBJhKdPNznxLUdn1Ebj9vbBtRT
GcJKS1FvTPcKQmg7sTqt6YSaDXe4LxCiJ/1xQCOx+z6mZZi1+Kh9trqbsJLWkvZi0WriZnVwqQ0D
9F34w1TEZioRQkjMP9eRpTQbkenRuwM+pFB9rgKCitPlcI3IX2Gu+KHfsp+nEaPSAkPc1gjEy5dn
a2mZD/1foQ/V7jFJpHheBRoxy9jgl9JlWbTjTvWx4zVCLxoOKU+IsHhMd35yPjMGVXFYuDPfXb3b
uiEZPBrh0euitFY5bUpCpxVHsuJwojtfgWWrkoreLYab+tkQ2ahcb+K7syfPhTshT9cFi+5si6UC
FRQtXFgSpWka2oTKbov7xIoCJqbDIm56xcmSS0MnuPkZ9QckDpSNZdEU00yKHaEcCaqQJJmHw6t1
HO0k8au0dirm4NbiGRLLT9G25AtMMJ42tZilb4XENv71ruF/EwTUurW9o+Z8s4SFNx7DqgPJ6pMG
Ny2gYjJypitKTNH20oB+1s6DvDcZT4XvAGkVAUGuZ7hunEHkBjK50Gd/MAZKUEMSPLle80OOks8W
/pOj+xi62BaXhOFWB+l/9d18fpqru2/rwBGVbNugTTSXN3HeDW3PO2vjQ4/B9Am4qtskEFJmt5da
algz+cc9JQZbwx2G8w2BU7+LG/jX+M5X1fvY+8XUFEDeoARGcxqeNu/tqhsMxDLfOr0jNs2hdV96
1GewVrpi9RAIkjWeSvXuoLRajarTh2uCVO675E7UVx/AeFjo7x2rGKg0Nca042HzBpagBQJ3N4db
XfYiL+jsv86SAG0P/mJ09y7Uit53Fsyll7y6h3rHLVkxXIpZ98Yi/0kBqXdFGfE7M2S6tPj+FJhs
CQlBfz42ykvA68SfudHKNNrWUyeMbbCxRAGRKlcBaWq/CwKjwL5Tws/xLNGXYghRsqFcKGuD1WZx
XNOdxFaRePdUKZNAXvSfuUAMzVODBZ0McEQe8w4jxkTwlSJW/8iDwWLp/W3Wz4olq5pu37O8b3e6
461tjPu1xYbrvV1OZo46NNzEBSARTeKUSA8lDSARhL06qNmBEGtpE04JhB2JxLhzxLSNxhaK3Eie
91ORX8y8sPtbkuA6spiV/ypwdHAwFjIoUclbluE6hHEDY1FvEBuP1Tfg9l7Mr5uUQIOi3XAeeTXK
5GGn+W8iMUhRD3xko+vMGV1hOl70b03YMh6p5zYzYzp8HzajeFnM9kQ9kkm1Xg81WrNfIrEW5ADy
sH2k8Py2nXDHJaQpDmK4/Q2iOXco/Fp4S/ZU7Yz8AeiE3uMo0ZlOgDmZDjb7/43HHnXr6YkKVzbm
BfN+YNNns6fAIjQB8PJQWEeHIsN06HmYmSVD7ai0Tj8l+Q7YII+w8pHnVLGEKMR77UVb+D+I2fw0
17BPSA904Gd4bwItmwWD78FukRducxx332dPuTARcxQkdoYmIvajEW9seamr3NUGRR4u/ipnjON4
2iSxQI9rUoht/OmHWJrO1LpdLM5aAEb2RWtfdcsX+YNwfejAVU9QH15x0CazEwAqTtli6V/s/Xa1
4Nb9aAZxxYw3N42V0zE9TuSMx6v9w6QxTnL0ofAZeYwHawxn+xrXTP/y3exvZfcnON+Sw0q8pyud
JTmI4mG5kd5k84KEoVTUVCtW864egdOHo1WJ9Be5S1iTXNIEFVJk2BlR0JT4mNgdiG9pBa5fT3Up
nuknB1SbZXv9OeyvQCP1e4riR8deYWZ287YEwyRsIuRB6xiIyrkYY8MLGo997WZeFWe0RfKjghf4
UZWxk3dGt91/cETi2r/Z/ZcfT7Lbwr95OLgkPWCB9mLaj+/r2bgGFZDnYup/07YLwloUmsKvZb2b
cX86hpL6DNPjd8TG/58SxSLBu3bICwCGMLErnIvCksDantHX5rdWmSrX/qN8ZLjH+EvdVgJxOfOR
aJcl12aD/Rx57gma/7FsA7X3C/nMsnqv0KHXHvLhh4E0NRdVHWvDHBkUtA9K5IjHfVW7Keejo1RG
Ks0r1LGGzTLOsOAo3qZ2R8H0fzNOP4/IT06ksvR+PUsVOb/OS+l60NJNbIooohcNAKBLlOFoF4Ei
Ym0ZFzx0kZG/cGOg7xtNiEWjNczgom8YX8htfp5m1RB5SqdWN/WME58l1UpFy+NkaCcnvg5BOkYE
BXibwSDvXV4Uzyqf6XcAvPip6f1TQXfVjkpycPe1mx2ADccwPgQ9/51ESvJa4/ZWvqaQLV2TEXnH
dGk0kdPu+1YmQ8FDVSTO/7pavE8xgTqg89WhcTnJezQzSgp0v5PERCAhWCFTGrHFqBIe/t6NIHD9
AN5w1yOj1vGSUJCaFhy+wc5K8WRl3JjffloVZm8Sphg3yhBZVMDdsVQX9a80NNxDpeNW9UKD4EmZ
w7nZ9mSoapFKUnUzdGwTnqzyO7V6vHgeYc8CvXLaHBDlVPT6LViu+/OHGv8uN/Wqw5R/549I9wi0
W2UtCDAuFhbUK6J9DWPcC/ZnhcVO+SXrTst8D1lkAlGlpgWRC7Pzb6YLhDbW0F6vNjTBQNbCnNc8
52P4/P/VNinocUG7IYdHI/XPuTz7PvEQNOsLqoQKrFTpc6yJmzyPJLTbmZRPs7GhezeMO5M1FtKh
XWRlVHtgoURiwrcU5gDEOe31ctrJzxwbDC99qd+Iz/8m3BXJUZJ6Py9NNJa/rE+xmvWW8Ffmq55A
gK39qW+p2wP0st4sct5Fim8hlVB9OKnbwVa31pDR5MbjRb7rTOU0aD4YjznYwOM6IB0YzSPutzhk
4RXERqkUtW6A/pZeM/WtOMKZZbEuHsGpwMzZ378Xin7zNkEh+m6HWNe1TCBOqu8lWL6rblvKgdSF
FVB3IH+apB8c/30+bfHXxk+smzYCKVPu/9CpgmItOAtNit9s7xALurV0OzQjUINOwavxuwmjLEQn
AJaTQTUzN6lYIQih7LuUhDIzEEbFiXQJE1Fk0wD9vVLgXzSTl7Z2sW/zmVXqmBHSmJ+CrUEClP2i
q92+jWGAy1mym2LbaJH93HhQHJJDCfNG1z5KD5WYi37oMhqoQvYeMQN5FutSFRZmxWkPFXF5a7ns
jsAySMZUYimrrTmdjIzse6pBUFboKCAL2FtuQQdRUXdMmNFgpw9JBfnJDMY1CkSW/lnZtiNjCaSY
ipnHiKqjC7oMcrJLtXm60yfrHLV8Vbcz/XwbZJCI94Z3CqKafBoC3UaVyLnxCQp5sr+pOUx2S6Ua
gW/HOWKfYysdC3VZMJHzf5MPZOlF4GVbBADunpkPAP9FPJ5SHxYaVi6QioDnV54OQsCLwme14cPN
ox6PjqNjvvqZnPLd789X+OigiLbmRQAJpl84xwUQOGD6YXtJIxhcxPnZE4zAghWpYnoJJA2uf6FE
T8B80j8gviRgMJampVGxVFokuIjBI2juESwdq3PF2a8FbwTiPbk8TM7RKtq9HMT8JLfgVX9P/e2h
qk72bAii8NNLw5JwE1CVvgiSNgj5jLXbqFqwOt9D50Usq7K07t5lN0bYUAK8tVSgHtDHJ6vtA9y8
1OxW8E88uS2DeCkiBdxOKZG+9KkkQYi09GUcN94Z3zsux3ja2UyGWDf3xosad0UykPuC+c16Cazl
Rqv9NEo4xlPxt4R9iVY6MIeNgux3Irv1eQb6uBZnjhz105aIBqSIk033OWfFf0z9uEA2GK/Z3jnf
QZy6/IGh0Fec6thoOKFkoVj78miA4xllW82GwxYafuwgvgCl0gJkjhXLu3yQFXrrJZZ0v/8gdTPH
WpkK/JXbinTX0IIpreOi4D8Z6P/dLk7jVjY/+w/KJDIFVM1DuTTHMYeYgtI3K9hc7wr36mi/idpc
dsvmBJM9Mx6OmOmglksjZ7NAUm5j0NcDTKX08Wov3l+pWBpZDgUg3mMYI54haY8I/QwV6lnphT3A
hEasCZ6iLoAPbJx+bSxYzwqT3PoHsd3jcgLinHNsRJ3Wc4cpxxMLJuxnLdp9PLGe8F1AYpA2Nkyy
u0sTx94mU7VLxCQcqm2s8MWZAsT96NOP6+4YQ1/Vtzf+VnYi7n393/xceyze1jgkn3jSMBY/Mcql
e0cMXQeDvro1TlyI8ZUcOSabvaZHesByjEK+ACQA7Evo9mGqDSFMIQFO5wo01oYb81PoZccSVWag
/16hvDqHZXrBz38jfof2oMYMaiz7eO2JBpt6dkIOeplqO2WFwxVsdZmZZMEYg8/YpaTIpXw+g5qb
nDr5rI2VF7CU6/DHsXgRNg5AQK4ZYhQICZiNi83+DilGintXSXWamC3jITNzfippWSalbZs7k4bD
nbMbHgo8dkrH8uOm6gBSqpfm3W06IPlFfICnaJVKGroQVqrC+Xr0plmjfrWSCYwbWfVpOOV7Mg4P
UFWn4CTNjE3rNSbSl1i6Tw1y/YRc59Wawsxdthq9LqDbvYfyj6i33XEyqTNu5OIFBlYs36v6akV8
joUz4V5aMWZ0npEdoeXY5bUptv1p4Y4SJl5icMIIQ6gcOQLUT6pS41fwJS/h7g50MvIPcXuHllVF
4ytM0PVvx+BycNg6XqjtvLljGu7BAR0AIs3wgcpj+dmYzaxM188zHIpER/Ldyipt6sVGfrrqWHtK
qAx9qXFBUQpGcXUIjiRqOzOgg1CaQhLtvBIK3CuGupZnSIn0o2XfwQwKguUCINSkCP3BzOr970nl
p7uHUC05dkyfKyeBl/ctL7LNHbfk9/cF+WuioiAfjaifJQBYdT67b1Y8H4OnLaQaxPCehJHm1nhF
D1q5iLrHj0eGtDeW8N3ExRhn1/yl17U2WMKh546v5Ly7ml25WoOsW4t1GcEDE6kANFymqDJm1cT5
DWVjtxtlAmBMUJhOk7EMIEsifQxsSZ7ZZm/CJnl2vvinbF+1G07/h9t6EEsA/P4g7mgHz+QwaabW
laYjHB2RyMt9X2bAcwXbtLR1pOlFbLJcFSbsLPrHFy7cDmSnsWS64DVYJuvjLlhqNUsTVLt0nhHt
2To07xCN4He+yxXyraBPd0tH43rTYyb32hVhL5vT1oVAfjdjcChs6EXVMP285o6qeeyTAh8joCDD
e1BBPxftjOc3SVUVSg0bl0bE/IUqPNtw6uguS5KA2Y6vuCgP9ZQeI5WRDaac0fXVUx1KSYtKeuEV
ZeFLCKOqlsApwbDK+t53BVEUjU36xoJ6J+t/z7LTB7ujZWhtusAe+oP1w9Gsd8IvrilmezgyanxS
rNkBPdmDuvoQm39UzW/PkCQICmY/E/AjlSRHY/LsnspJs/UH4D3RpC9X4a7IgwWeJ64a+7MumiSd
qpikU4pt7dm2LSb6GJKzBmO1VhiGoAuj9iKFNsw0c5EBMImQ1htlxYDPzF+DWjSqCgflPW9/77zk
s9fZD5/3W/llQbK2xQ0kDMuct3HX4Xj9xG4vi+Iqvq4dT1Bh4I48MnP8BkHYHnPN4aRQ7ukf8a6j
odxNbrxTV38TIgzDqtJwLLkLYaLBK0JRVco+B3Sw/SSrLoP+aKbUXiqVE779qX+33N2nzqs0tdVX
BpXCUd9UDjldC0TEUZzdddU6DhUQieaZVGQiX/MxPV74FMOSN/RIx60ZsVTEXbpAPNSJKSBv/AHK
/3Ur/BmyRI53gtUr8VVl0sjb6TzDNbnmFxmUtJ5a7o+TFO210muJRHJrotnx+qZkWa0gh06RFOVb
FNmxeDonTVaJzEInuaCG/SZd+PcaXlW4R+wfvi8J/iBGxdXTzp4pODroyLiDmmUBFR4lNPlmAWT2
ysBKr101HvLIl6OkXJ3SK84VknwY7cdAfFPLvMerHb2niIsWLJ8DTJsBgUs4NhLAlqAVP2TS8uJT
H0LbjZlCRjraLMsjpRL92VkrgCUDoqVBYfaPfoJzVCTOOeHxPUIyEPyaMoPqFBquFxgVsYwgjDI3
DLbCEfidPGWfwcq6x7mufxgso/6pGY9HozYbOGr+zY27nf5qkHvrhfsl1dCIeY8T4+CQNx7fZ9w2
XL/x7GdYZ9yfQCFMwoJELPnLBCvT72j1s3hg2h/SYMb2kvExYeqFugJRLG0vZXWuYRp6WszDraKD
AilxJKUqPWQHq0t8yia6zwH0FX6BiCPjm5qbiVVEWxsbQxxVhWAD4M2DYZiMDhKWiv5CH0x5JsQ0
JYIAwQ+IkI4QQksK+jJl/0UIWVIBJzRR0fkCAjbUqXwP6c9MvUi27yrEYgAI62JvvJYX5T0KHDoN
GNvw17cu6ZnCYt53V3PF5BNigG6JSarbViIaotUTzhjCzv9eVuit5VOU1K1E5JKHk4V/XpvsWcY6
pnJkPmfwSU0dPebZA+glHYv7DSfC/VNyupnnw89md8Dk0TtFW5h+IGN3dsHKQu+THeEfoi5tPdkt
qJJEf6ZVAM9Vp3LvZLJd3462+1KPZsn1FZ9Q96xe0+M2bWkQ1hL/oK5UUTt2EjEHOKOe6ltcYbEM
r0BVOJ1+02Be5Bs37KDHsvGxgCHN/z8QgP8LZsNZXq9iTix67K+ZhTxYMzvryHQphKps5rJgYufJ
zZw2EKgLowoP5Z1va27Qvy63jj5w/HRY+4/azIMk4fNRVC4zO7rvzLciaYQz8Ithb3Nw/VkqzQFR
cPRlDv4/lMX8Et9GDLTwAxqLcyeQl4TbCtRhW4aTQ/PEswPqTJRBg6CaT6603O45d+fA9ivcZ+A+
0oqhR7gg4z38ZVXO6Y7vUXAuv2G//sB1Ez+tZFEMG6s/qwlifz4bsjHnUitkvNXEfbptpzFI/3Ad
UbIut8/hKBVrjAbYps87AcDzOaNIhVIigmWeW3OwlaBBjxTbgr9qSntDVc/i9EgwapmbfShZU+3k
0kS79SbQEMlkqTiA1PGR8DYYtmp4Qf1H7knKWYpZq6uO1CKk5KVOnYmC/1y1l8kNbUOhD8CZBFdR
TjVD0bEAhRuzZqws9+8v5uV1W9FpKWCmqJ5Yk58sSJqWuwwx+ZvsGkd37gAuncynI2gYWm7N96/b
p15q4bTojluBzrZaJgt7PZ20Yyi7V8Q4eiWIDK918zHOwc5OYhPW7wrOwXRHilMkIptbi55ZwLMb
E/CO5qa4Uul9DnqgHw7JrQqEt82kzuyodYQYyh2GRQaPkgO1/88DsPPMScWCJmZEVPJJceE8TEPo
mpmmia2yVreIR2jko958t2GeNlB5xX+1JN4VimqPqBm8J6WjFrnF8jAGBXIyVCKPFN2tiw1FcD27
pXYuo4C5h/jCNeIkYO+mY65nZH2jLHf88YxcLsOQbYQSsuVXFzwaeey3CWExL0GzLkdKM/za4K7r
kSHkDQA4tuIpAtl0LOqPN6grDadckirxE7+1Ce9mP6ECd0uw1LYX67bXzo/LJaNnI9lyUmS75zt+
0Q3lvpfj22sITXCLxnWneLgRtGN/XYQQvc8j6FiZ+3ItEIhC+2QQeCl12Rw86L44tisy5g22iHvU
TbjoqOyQkfIySDPAw95fQvoaXC7+QDzyKR0fj386Ow8HZcmX3cLgRrOIlkkZaqV9zwjkwRamPxji
3gTt80j0550tAhhVTvbAq9XDS0bx6k/BWxCJlxuyaVP8ptwNU3uflxtnT5wGgjVqPXbNH92Kxe66
YqgAMtvWfnbece2QZ7xRcN9eN9hK/cZMv3rT+GDafn+FtU06n0Jp73PCjJ05abzL7hcXqE4Ebnew
qhO5Mym/p7TvmhSYpXmSifH2Ls2auJ2LlLPVF8kif7eRLhRK2bMyHCfLlAhSyagsav3MWaOKahmC
Kh4hsCLDPD8uF2aLGQ0dFB58+hl5PtogFf9T6z2PESBG1UChBsW5DY+Kjr7PL3o4dDKaqY/YpOtR
PaVz1Uik1mNxsXEjM2ue4b1tE8NTgmvDVTC+/kvJYaSQK0FZDSBCsuoV81GKUWs7eAvi27BqZ4OF
6a1fVvm5XNsPGXgHsuhX8XF8vyIOVQXxj6tzkf25kqB/1WAfQNXfxpggjICgWvpkstzatqahUve6
DZD8wysqpm8/a/yvywND8HIpT9GrQxoI4mfKsLxmRMBjgl7ysdTElxKIX+DWFsyZbTsa8Tgk764t
DPVLnG/eG+AM3bpQjBFuH1nt03Y/GmqT6dhHiX7WqskofA0NmDbvGhGcEtPns2571QkxmdN6Chnx
nIkuLTpMnl3BcmG30hXYd7NCbmyEP21mHQQkhCdUCsH+n12OZJ3UkMgxNPAmQ84tiN7zp6uifvIF
tK22ZDz/7c0UjLZ1tAYBXHPPj3mpVht5etpb+ECdi7dPPZn5XNHJisSSWDBLd06KNlrWJ11EPm0b
quS8JAE0mlSJ0CB1NsrsdNlv24meBVGFLARUYj+Dt8Ptgm1jzY9bpx5zg8NuZgcUOxk0vkd6DniS
yb9wU3AzwpDE+kkePr0bCSceARFBulZUqLo5ixaCbVJNtEETYipjtP7BE1wRzYIFySoDsZiSlpL4
DzV/LrYmj7EwV59qJ4dLHTK4z+qFanj1qhjxg3P5m3P+fEh+lSldywgq6yyQV+O8f7CAhZKw971D
R9seMXtwdpm1jKzq61+SGuVqfqL3q0KxHqsVpU7C42tPLkP2OseKTrcLnIEf1+B0LrLWldBnV+qb
1C+eGXPd/7+YNQVaFPCkh2OOoTh10ItJlIXr2ecDUpit+66GPf7gQhuMjIm5Gb3dr53gDtbKuR0R
ALgNERkOMOukJnFAsHY2MIZTDABIB+9g0Bsncke0FMhSFpl+X1F4DjLVh0tfvguzeJgrJ5lvoitK
4Uy4rcDxBIIlOIeu80Imy9oYahnx5uHqEBD0OwcOWhuB7hoCIkvM51RSM5xq+FyHjqOfpqdWwIY/
mVTxxZmw1rYqHNX8CT+ChilHgT2r2NSuuPNJ88QCKHEvNfHLIplszhlyhrStMhKxbrTL1SgAh0OG
+phivYHmdEcx0ZkWngeDhs329+H2hDmsVUYzuv9g6H5Vy0bvRsCj4VqNKOSImPikD2w/a6bKjHT5
ojibyRDbICLYIGgbCDL9v0Cjjbjp6YfdAjufwiBNtQEJ7ChvqTMqVut08FaRpJbjKCWajPlPRehy
9GmA27QTZz/PnKjy3O3cv+1neCeBMKkuTqip045xRsUmq4D+suBszgPu2XW10kPC1EoRSER/F7Ml
EoR5DN3LWgOhlfOsZkoBDYU1EPZ93r23VCoHmbCT7r+A0kOIDMKYZCPQpOTZMhU6f5Sky9DHOH+b
Ov2iluJC/tKbdmqLNvFOcv/MNcJVtFX8WPn4dYzAchyeo0QVswXBmeIqVsif7Kbc/UEk3hEifp0T
hO7mh0h4bv0vkm5V5ITqaV3QSjialhg8LFDCN4Ttv0aR2Y3REfrmx2dOEEhqG9S2uqYwmRIzL6B3
ikQ1YwM9a4TSTnXQmKVEVR8PibFyHUEhyp5x+QlY7gwM2Yr77z2JBm2ItiixCmIj8NKEA5Ujhwhe
azW+6U2G4HzT24HRdT7Ez+GBYsj4CKOMsQn5aTdL2EaFudGYntK24mv9NznFLV0t8T3aTglWmT2r
ipOjLP8Z8GAkM5UsRTQzkY5lDB8Cax7yMiJiGLGmBTLq+U6cNHh2MnDigQWKVt999V86zKS7Dp0m
XrcUlR40PbVwFiCVCyPoFE9Qvx1b1PSesiDUnhEoteMR8N82FQAHs2cHF85BKV6lu4GW5UCGYjtk
t/F6RyzJ9XswEIK/cFph6yBkXjq3tdY398W+3+tsOp0y9XXqcR/FjMiMMSxagu9KFS8kJy9tUJfX
RBKTNBxmhcdlxxTT/m9iMJt/8huJAJdWr5mY6MmLbfX2R3lLjTj1IE0QI5aolbP04QrayaV/7vZY
AHP1JaV8DJvkbWQmOLqqWbS6GaIlDJN/F+hfPBpX9se04OKkl6tAR2m5JHFJNPq5Uq/hR0DcvGWA
dB4FLbK272B6zFCc7UrgaL351NCceiGxWem0AVkTxx0rmsXJQzxkHDr0QZxDQoQsadtSsgoP0gin
Ys4nc0StbRUkGOBPHCVQcT95HAJL3m+Vmdz58sE3yWZUk6+pxyybHblHXAFr5vsH9oOuvV5WRe5t
u4I9Lu7qbTd3Z3WyKY1N62xhURo5HC/TCINnV3vX0KMJqeKDVNidXPuKpSRVGi2JsYMwrL9k1swu
/ryWrDiiZKlznQ7i1ppromDEnDluB3OJA6HfYSNyWU9I9I7xQSIX2WJtCFHDA0QwZAalM+F8vD+8
iPQvp5zIlhz8fWNmuVXIHUPAr73JPcSj8vQrWjlBLISt76TmdYiMxj7iLO6wiNWK00Hka+ACKA4g
MxAqX8keoMj7vK7J1Gexh9d8aMiSPcRCikoMNg6QEc3bcOksl14WQvTixDKItQecWFd8hzmKfPxh
jrcX/olq1Xm7b3noEpAh9l5zN9VxpFJRtcA7loG4aWsaQo81hjZHDnjzXFnpKo91qSRVDcVrXHMH
hvyLAKCyAl/xHTtGJmJnOgp9x6vqYXMG6DFrCORsRLv9t+pourWo/YBeuzZcyY8d4lk12KaWfYy5
6yNcF2HG1768VSMSGLw9pP48VV8vslSHs/Vjd/S3wrRGZIk6Jh5s6FdTjpvY4TfvR5Fj6GsDC6AR
4vaIg7XLNtfF2dyeEGFjpgs4yspCie7eWdz/sW/P2ds1YaTRjkH4NHAbWyDJ8xxR5gbp+kfPwVQc
8KSK4F2US/W48Rf3/cflot5kB9OcBwc+n6Tmr/obGPsUBC8Mp2jXWlm3UCgoZMWLLYdHRpVlxuAv
EHk8CThljmWN4uuhdOkaE2s2CuTR9BNXBZO4OGLPQp4Wvh5SVwjc+I2GNF0BCdH8muPtTeqI2feD
j0PVOKtGEiDMIMWMU5J4p7xqBNEkHmGTE9xhfAY/lrS1kUSdCRyF/mbkzOhFaw2YJ5TtU3qd1pwx
bvhWWIWm4p9ZGixMGC6G12pM2U8kM5YD5aKDHdOl78XAwzOcOtWmWHpdPi6Ybxbn+9a6Ot8jPTqR
IcS9OiU1xhOiVG2SoJlzgctfTYr95c3WzhCrnsv3T6FKMiNV1NIPk/+W6LWwAjP5lb9j+kAddK9t
OfWmITaZ4S8mge/QV9a8GcoCurkwQXbqmsw/zc+TO9kA+VV5kqkAi+VgWsoFCYxurjdQ2O3aU/yQ
K+z6J30SEbITsg0lex8PSKqSEA8RS3AI+SuUnghKUuwi4C/uz6er9aFEkXmoFte8xYATdkR43aBM
oLkK2wIcQypT1PIiUQoSJvQjdfYB6KkRGPUUcIDq4Td+9WjYurB9z4z/H3IJvniACFjAY4l6Fw1s
XXj537St9V3rzrEy3Z/I30CXcedyk21vVtRxG/7cViu9/MAaQ100nIhRG2+Tnu+hVauYkZVGERIT
yox2pqIO2U0kviHZWSTE/rb0vYPQmjpIx4MOo6eZ34xZC9y9U+HiZcbHJiJXZVILamT/zPqF1H4H
77m36vgdrkFodEMOXd1TyFDyrkuIltkB1dXYRg0wgS51KhjBvXA+glavzcnFXKWYRXFZpZ840DDf
MIc6Qg44g372y//WfJxAJ/4D1ge5QqRK4sTcn2DC7wnD/glUV9ILvHMRn3Q2MsMVJRxB3cV9JAmN
aWUCa6eYWJ0abyYCQlAIaiBZx0nkkM7MhmnAgwYlrZFlyZvlSSdXggboKBLyNG1WB9nj46NiTARN
rT1/4shsQy7PfZhQrmg5CFk+yQH6Mfgt0GILULNFnFc+5YIYTAa0ig7qgpV7qjxues9J9AJK3pLU
aQeHfFGCknxRkMibCU7cjXo0Fvb0SlqICrhjPVNBciU2lPbDYoLcway0JBOmoH/UAuyA0I3ecDVw
5LTQA6sbhXRgX8+PSx5rY8MRCe222I383cCY+ncUbp3Jk03LvG/DjKqSIGBZG64WMl73YImihmh+
j33x8bF81HHRfQX/en+YrVqmZuvEFTeyQ6ROpLxkXERcowxKyVcwTTkpXo2+YMXV8XRfxXqJYfCl
QKGLfzUmy2FPDet8ZTi9ckTgBrNXuMJvt7pSpR7GoiPgwYpumgFkPpT6IG+7hO56tmVAPnU4VrOV
3XIto5EUg+D45qMZcj6AONkWVSEw0w2dzAU8htTGM/eOwM/RjYyY+x8Zf2I2pnYjTT0uDoDHVVNn
82P4ZLQHGijeDgoEoI4H+1jUmvoHTc69RX6o7UKhUGcxZ98KR/DCGIBOelaFICip6jheeFfEKxrU
2NCKC0xeLkpbE9jhPeFyIiBnhIVVljwY1fNiRRGH1zktpoBcvNOIEKbHDIw/829ZOYTNCZS7EtmL
ITn3NOsBQGQ03ynM7asspJkrt5FNcM7tET/ERJe7qOCQmnyBY6WdOX5tpDt1OEyEteP6KjZv3TVT
p8J9LT63V1STvlkbEaD6I+4yqdtYz1uxzhTtoaaAiSqY0vI8xklY8JObifM5V4UztzzHpQtOF/D2
IQySECaeSUXbYGlEChI8ONRIdPah50udV6qeVFXN8BKgp/wbT/K8UU5StpT8m6lsXPZLb5YwGknc
aArny3iheNMnqHCAhUKn5mypB148Gxdw6Cpyk1rln5va8BWZ5yKwdwavaN2V0AUlyc17NxIQlpAO
VzEXafCDFeAGZCpaiYWG5pv+pASga0qEoRbNw54lBQwrOfmgSgXMPNUEG0A4F3Mo7qvaNZGvm3lR
n4DlrcmxJ6/B3U/vcgrReyhffQNZ3iRmDlc2PBDiqiuyfXyth3ZX66JNaqPCQsEddIrRhm9g7ZCT
X588KSixemih2r+o0VjvZkvF1ymwgpabSJVo1UmMOs4P30A9AJpAWK50+I8rVgEXufxeUI+SCF65
7UlqFjFh84zbgPgbO2VS+hq5eDAj6gb8bcgTivTwNXv8L5LoBpd/xSrwIGdB96/Fa4nsbzbdVjw2
ozeSQ6C6tqMpb+C02OHn/Bj+vYcp6aotoMOMo6Vg/V+ZTfl0nXScBrBqnIIalr7MK6PP+1txWJi3
clUkDF0UpbUcyXdu53x1K89m5N6shYFwk3XIB8PXpsooT0fKVKm1ZONIpnU8afiFEfTy1BtzBRjs
PqWM2JqigoPcNAmm7C95VvnClOJDAkvWXVV5MZOPO1C/5BP+18CaPq24+4AMJtSCHJXNIe0OQlmq
McgPFFsabqFwaNUVbC4x/nKzmYdp8RSqgCSXpF0NoziZ7gK6wzQbX8M8udo8Pm3C8soKHrT9Vf5N
Ez11jJ1g2zvHxbIn19mrMJZ1MQRjkWHjvAdMBr3vNNYR0JcH69m+IQGOteTehQuxVi4Kygl3GHau
1bRng+0RtvrKE0raEOfbZ0Fe8MjBJnbVS8M0F5ZMsk9r08eU4AppMt+sG1I0yceXVBfpZhCZpFw0
C2o/uCEwE5Pc9tuSVMWDLYK2Q7W9YaowWr2BFJ8Yba6THPrBfc/Lgc5IFUjnldGBNlqqcgPAyuHM
nCx+eqvADMZTmHM9QqwZhJwFT0BcqSZO+ffcZKNiFmSPRFBgxQzbkO8KgWrBJoFE5glKzKfgW+ec
jyd2o7dTgtKCUOtIqNowFcwFAR8XA00ZU5Ieu1lJ6c788SIse/yNo+TpRZfFuxh/0qS1QDjIXP/l
rAqFkCLQsPqWFPIdHMrUtXFHVH9KGu9medLFjE7QacJMJBICp4SDL4vy7HmdP2Sy/g4/dny16KHb
spku6uMTh/J3BtJJKWcEsXeXuxdYM7bVEc30dqEv+2/f9ioFSwyHJLjI2lIci9qtebKMH4Jz1qUv
ZdXOQy55hXHjobTZgx7HIsxtQuPgxq1oEazPZM2uJAoErHaAevSdMraKONVgEdWB3gecKaTSqZ6i
SZ7Hcn2nmFef1c559PyeEsf2VISyw9PgR7D7kxamr90oeSr8Qa8PNmiJlxbWswHZk1ehmslXZrV4
6muAQicO0kIbQMg8I0Ehy3h1Av5seh0PUZVUTqfM2QNyKqnthuLSfi8VF3/BotGSkvl5FkM9dniO
7+AXKQK+O/BDQviJLuHQ1oum+rlEMdESGaVuxXyNLj7nSPy/obBQncQHXQrcoM0zBrGmStjXEwT/
y74cONvdfWqFhojYfHCh4Oj+wYgp/4xmOZ5LszwTFpiliQ4MuonzCtrtj0yyRWB3oeqqz3VIVjbu
Gmty9RUNnjyglXlWucIhNrbfb1gt83ZpDD1DzdQrDH5YIHkPiL8t1HsChdDXjtequywnh3QQEOeZ
3CQC0+fQgrQbyiU+E/7w/RWT+0tXwM568chJBq40723fcehFb0OCFFumco96pRvqQKzmLNnDJEQZ
CDGL2NhUxA91XgChQDwVjtvd6FrCKaGQpqQkkJaSNO4T5BrLpu6MPzXq6oCTm+IhcahfL9YDkg/G
gCx9uYA7i6i3y5A0rWRxb9DjFFaa+msTTqXzyTTy7nYB4buqakEtSBnudacbx4J1XfgY/xyw8J6t
0cU7SP6coDtZ5hHGzURqzPzlFI6dJroulti/i4OYO97P4/PkLr3MlyPbNVtAjRPAeH2BcmLMjLxj
1mKbiGASo5p2rESY5Q7XCAFSZ66i3PgjUU6ve5e6Y0JKTQuyKkB+g0Kr5TYosC6bmXM1AcpYPuBK
CpdcrYznhpxoLoGTdubWtlqeV19k+yqY7Ly0vzkRhqXdG6hjTFuieaDp0K/VwegEMk9vEVeQG/Ri
pPV1l4m7UG5Ns4SgJH35E7dyYeTxlNGdxVgUe5DneV00zq9Az7ZyHQHD8B6BD8pmGIMDHKrTt/8j
bq0eLIP10V2qtItXHdkyqNtb+JWrjZ0SXqMiUES9h9iOFhHfKSh9EqjudfMGLYffSRDYOkcm/O3e
yps5U8fhoyzWcmj0O9BXN22QmmX/I4QOiPTPzMeTovV9k2bjFbqgMTlm6N9cX2dBmK7ln6/0A2+S
scHb/xiCEswkhHk7Ys/wvxBiX7lXXmwVfG+IIsJWyRuwMViOsAstqt6mGq6Qk3mucizlEH7mKZTU
Z0IpoCUU5wUbV3QkTEc+Hxm8uaNDAGGPgGQ6K5UU+4OogWh+cio72HJ+0WFsqjWtI6IGDmY6s3KY
ZV7bvvNn6v+4Jy481Txu1WfkAuw4P22JJXx1ei15UpRMWgIl/RMoA8gx1St8XyFPSmtSEs5GrHcB
fl7vwE6ySaKL0VkCWc/YxbR03ZvBlVXi93mpEcUHo0J03zqskWeMWvUXVXuBmqCaABAcaCnYfK93
y9rLNEZAkMQvIumK5RbcwPzQ3xHMpSOe7fKLgSlLwzBzWLaOmbeRr9c0jSTtInx7OIVTL22Jomo8
o4d9ft0EsVpWQBTfy4LR7qKKypHggiO4HoVJailG2SJYRM4qv3GnsM0A+nV3bJj+cisSSJXPXhXT
0XltkJscap6nRIpQ95y94CGzqTAaYIME6FJdiTPo97Lu82B8+yo2fYDt/CVw1dt6tnGiGYEfpE2/
6NcbVhi4DOqzLMPDnqrHl1f3yRRV/NfW7LoN/r0/6E4z4Dvu9Cx2dhiEAuJKIm9R6jysI+nvdzMZ
P/cquNruzZETWQ74o0ElcwdsTH+wfJdcaUU64lRBLwBTehmeMZZVvDjzwXpVQoP3vInDQ547K1R1
UJ03h6XNqemlYUrLvMLxYSrqO5Tu1VMlbBffcIHfBQ5kQj4E7Q5Vv/oR+189nldp9jq89vVGDv5P
edcd+QfbawA8VD0lqila+Km6Zil6+gao2aHlFO1dDw03rY5fBcfTooHAJuUcYtKY4Ytctwzgj+7G
a6nyvqkCFzzxwRDoResEpV/LPb/7qx+7nKvksY2y412CpYVTl8nvuQvr4siekgEMnSny9lKDLfft
17iuftKpEoorA0OBTUrm6wj7PWVKu7knQjhUlC12STP/lB4WzkMIeJJzpNKMV9QUWKhtjcLwivUo
VNUTnmuR5PWH0SgCSmCGYAuQzwmKvR7uZTaT12fJh3xHWJ3TXjF2RXwhJlhXrw8rFDR/R7/VYuq0
qM2au4r5AsosVg9VnsMVMH1bYQJ607x7Z6UxoCEgPF21kfULsHbhEBv6TPU8c0tdAzx3sQKrjksX
/Az22d7WA/NaolXP6KD0JlZzZqEYdg3fFSQYkiBM/N6Y9iwIp4r9Z7K3FXorGwj3L5DN5kFbqxNp
vF2OpBVlOm7INy2pARmWZPJtGw5jgGDd8nc0LFRC45vo2e7+XPVzEG/Ds7ropyDQENOYD8QoEwlV
h6sKmF2B2EBGx04BEkhm/JACXZFPv8opwacJ2TfAyScQlPUXA8kJEQdOp4BHvB06ssN30NcbxPMU
ELipmiDv9fgo2V9R/YYEm5SdsJ1rdzGOQ4g4FxQmjK+SlNEgfmC0mJnUXNltda029jsXgqHjsln7
Mr9ahcTWdJDylk+aMSC6TelR0VT+pbC4nuppnNOha7rkuyCFf2V/IS2HvFET3LptT5sGbJt32uJq
90MpmVUM2cds+M5LrEwajt3hSfPS/cODUAK66+a0vsvNAzG60DoW7aZpcBx+Ney8a4Xc6gIAkR2C
LkO2mN6LDqHFv9i16dTz3nETzsV89byn/I61hKAwSGqod1JKrOT2QhD5sXwbJLD1wgOjV1O/NlAa
3U/JVZKGLzJ6gOWdJYI78SoyuJEbyWkEcdgs7mHXoQfwxiD4KlbgvZcBGTaJmhv/QBQ5NCcbSI7m
gEiftPSLv4zcAr2xH3Tw9xFf18Nhux5HtwaNwRwGuN4q2tRgm7q1zisbtMMq6QrdhwlmCyYY+nRK
m9ErJU+nhom7pFRt3ADCJy9qO+LJm5fReZ91g9SBdJMEQmuaMjyhVgjfrhLCO3C73fh/ZmFtFhm9
tISVBUFIxZl9X0sGkWU9c2PZduMTGDuNFLJCFFVyZFu9NXg5fzu3DTVzEwJrHwmLajwHeC68pxLa
EanxPwTWfHaTCrpC+VykYXkyxfsJrvMeZd0XMe2CHxYwWsXkbauQZq5GLF/iAgLV77d6/Lb2Prku
UiWNg7+QJhDHJrZA3EOhzBGqn7tcFmcWj8L/Un3++C9O8TcDLs3Tw3wTZUbHKPNKoZf5oFo+cvt/
RJ6uzOmnA6tHxsP5p++nHvJAvBGeIs/nohMZgoeGe7XtvPFErPQ6D1kDFsk6BK0UU/X2UEcG4ks/
S6YrDwHqc0sdiBw1kA20aEWFINmKB0T/KKr/tP1FX9Jo1+OGrPtWMYW5/BcKXUAMI8HK8AEliHbw
dKwbvM1Gdh0oGqEb9LSCpaIbSXzDYQ32hJbqcQQj+sjTGTjfdX/QqGLzOd6wOgIs2ybCJMqkeFg9
SjyKRn8T/1A/Nn+heqHAFmZ3/oVCpb7q110q07Y4dBakBWldg686vRY7H6HDf4WaOMUhFBAYk3yq
djo4/MEb3ZVoERY6ht053fJEgV+X35MZu+xqQaxVVvjRxyEVVLbu8NV7ZG4nDGX27a5JzO6iC+4X
sk3BXwqAbubynnzc2jUBCRIF+4LbSczhghGRc2teQkwbFhU2Bovx0QXJx9fNUIfqyHgpVnAzItp7
xe/7uVCgpIC8pnXiGP7LQPhJG6hk9E9Svybh28cu/+v1NEBLF7fn4G2bMvEe4CMLASgJ8HIpEVl/
2f4qYQ5PgHLh8mK/UbA5H4DQUk8l2TgFQ55JZ7xoMK88NPHA8WGX8aLqiRNcbDScGaRE9I2aniu0
8n9pppR8sGJEsFER4CT2TONizANl3jA6JXuC2OSs+gTXEe+swR0Ne8yWqORBpAkWEJa6qMozEAMp
3+oXyVn0lXthzxNDzNMOxYUcO+dMptHxr4BaG+oc0fvETbUHGVGM5EHmizJQCZx2vSmOJpO3TZG+
V7TYY3wvE2hIpzZw6KM+qyqP68QHOEO/z14sW6VBcS2rm9SBgbLHOSy+z3SYBZouzbVLrlq+iwkI
BL7spD3a2tRN6vDLSyCGl/Bzv4fV6wAYNQ9M4Gl616WKzMTyGqe4ljiCAEyigLljGHq65+as0Tja
nlMhn37hAASl2SFt2ncJ28dY4y/dMeGywsZYw4zicXYbzEtyAgcWY2tWuT5y88+sq65Pejxx2tlK
NuKZeG+3bHcoeIziyqEjkXJBQi0DvArrWQU3FBR0gp2FmAogtaqkasbSr/Z8gnOqA5c8rcwGouxi
ilgVVdan04V/RV3Ynx2cll+FQAvnsDQMieBn3b3LXyOOxbNrMxp0Kepr1jJefpu2O8zr83AlBYpw
Wj742n7AbOeDhIojW2NswzNNJKIwa5kFCmFHaBZbepmF6rcIxAPjiER447gE2d1nCx7E2395RJXU
SZqvBFD6sCjMSRKzbRNcLyR1M+MLLS+9tXmBIQjgcBhi/NrQbus5w9QqG57G2OszoMl2TF1sdkAU
2NQo4DFUafpNNar3FVwCHSeoUwuFi0E9E0l6LQiIRvfU6E7fiBMd9HRk2Slj1P0RV/eL/xsX/9zC
7vagr/t5rz6PVx57G/v281ZDtbU6gamU3kwBb0VQw8vOGV40lBNjAxHeUG+AvJOjJDhvlhhJUTTn
IXZ7xrXbjqEU79anCSoHFW8LgFT3Ung9JLPPmSOPAee4/VkpokqHMPcJxqv/Dx8kNUgQk8Al0YQY
iQuJ6RmXWjmr2H+9O1fWTjHZnNFU5GIgWnXGbeKIoBdKtcpvuw6ca6lpykkuzO5hqjEmGqyewZm+
5ZFSI2WRFqhsNtUfIVeI6sgECp0s/305Q8mRihvvYA4sriJWJA+4Bo8EKQ6Tsn2cphvDS02vlH33
5Hu1HpNHHkrZgHk3r503jZdi6Gd9pkXLR5kis7KeSxS09RF+9MHT3ww3HwUDfE5e5pcCM9NRgD1Z
+xqHz8//JsVMSAcF0mTOEAVwnaIm1EEEMo49/ObbGAP6y3SyIgxVYTmXwbbSWLZuLCldXOAzk9I4
LV7e7Pl/YSmh7PeIB9S5Ohg/y6cuW5sv4Jw3QPzQOOZmNXNkhUjn8EQxMx/4QfXMDvwVbzBGStSl
F75b0CiZOR3kA03IIBN5DVkFNPxI9A0LJHQf2hywe0/IVJTevTcKj7IhhZ5WmUi8qgkJOOZs1wsf
FwU8HG9RFfRDe37HA3ma83mzcFzROQt90FEhZ2GaeHpmKuh0QYuhOW+zRnqo02yWjJJ746StDJyn
qNs4Bf6UYqusO9GIlLifLb040KR+qkojT3VIsiWqjk3GEucySFMbIoTtwuXledab3KRRcYxDDVx7
W8YHcmKCBw6rtIe87gw4XF+efz+0SvcJ8TvNDh1Mjc/aYmGJECokxwoXDjHJYdJl68V5n+IpNj0E
Nz9ZHgrFey9h1cAtRNCSLPcQm1rhjmjuWYAfWT7qNOeYIbBeo5rMFm/0KbCPRDkJAzcvpm6FcOUd
FpkEtFpAFx4A/Mw6DJ0wUsJuuksS7nviF5+yOEF19u/cHgTzsjSGo/sRsLwhINrvfTDPEwhhc2TU
bg2g2gUKoGyTho58vLI8ZufJj0QDgjaxQCs0K+nGCC8SiUJzL6+/NGdVbiryuKoiDTbmGxMHOugd
T7kxTCDITJ+gO11v3Y7pCIyaJT6shVRo2QVWhApXqKWEbcr8G6nOvyrxow01NiHpSJpqgIUo+uZ8
Nb9Wx//bVLacPSwoE3/Hb6OniIIAdcjcc2+XagpoJlCEmO7BUtL6/M/LZu3rOyIgkq8UItLhZuqu
ICOmBwmqQiax77UiDCw5yC2QvYD4VdJEqiBQaNXeBIYvnzmNZ6ZpOAEhJEHr6PRekaHf4+lIKZ1f
N+AFJccDSHw1QlWTmXERVlb108C9pbP5WCY0+IT1feeUz6YQQs0p4qYZ842fqjDFwiGBm5Z27uyg
qCb4PGuUKG0+zgkALZi+EzKHWR2oLEnVpP0x0DzaOWlzcgrEqohrmlma8tJQbvHctgMvGtuawz/r
6mZuJ6WOEjT97IarD4gUE8gH9rWxvEOMm8odxExSmV1SU/YtuS17AKUGqu1fLg9eBCm4ePnEywhm
q9f6EQ4+PnKLx+AvCYl8e+JyxalE5UC398FNFqzeWE+3BFw94/4Uc0hWDqKuYnJdI7JFosPivk6b
mpZv4EBicrctHA1GMpW2Bq1r8luwU5zz3fDvJbtkRu+0/JaKI+7nqwiMo+okJNtuL2jYD7TLAPq1
c9HL0pL1nrKJODIub1MltGb2lvdQsP6ckoM77FXyiBVTu79lZi+6ZULjxOUxUUe1IGq3RJF6x772
MpeNu4Jjk5RfCVst8xyuLPVtHttJUg2yFBKTFwfs10v20WkT9sEnJYV6ct8HvvBJ5sjfRMRA5P4g
oq/W6+4MrHj0K6lsoGLlF2OrUB5wVWP31IFRfmfAlskisFDSwcf/OjPizvBjEKQqGLEfJCxdAjPi
oKQZVztNgg+tt0CG33aWDLW+KOxCVLv3gvkKf5CMuSw7m0UN2WBS7wTH90D5fNwk3qJ4T/EwDc3E
vcVbYIqHGQsEwfJaPrvm6u8ospK9ZM618sbB7Tor+TH4OiOf54X5IaRIh/wWrA6/0BKGvqMFBB5K
wh1pDXTKSSvVHfTus8ENTc/FRR+Mz4DUYmrBzHch1i1AkRwVq8S46jFRd7UlkVO5B351pt8UaoH+
El40O9sS/uxJqdM00Pd/NdxRB8PlHAgAdkCwG2CdeljP1YGLcGxJvKMujZ53bPh5c2UmtuB0bQFR
qfobh3qFnsMD8+//Se7edzO0MStw+Ss5u3shETMVnGjUKD/Zb1c+ZNO+F0ppuo2br9jy6MMLrvf+
kkg9dX5Vs5eBCl8Mhize6JflsfYTG0JN/K4DkL7GAECLu77rk7WCgxNSUK0EWfHDUOYTKscPZxpQ
Db/7K0iKtzqpj49X1pkjlRQSO19qQsAcV8Kpj6gM+NlbA0GEEeZd6TuaWwnWe3u1/QNhKlx7MQME
xtmJSsUNJ4qHVZ1riraS5jhjAr/umcgAT135fr8u9cvKugOuA27tOgQZjpPpJepV+OeczWzkuYem
iDA67Qx5I25kdx22cvJ1Mw8p9Gf01H6MAUeGTEPJTFi9L5KQIqd4FamAPvmRcSTxXOYsmp7BRJZr
qGgnm1B21LYVOyN+BXjaOTubCz7kVpqlTRzfJaWvfjfOTEJG4jMyg3o1vL/pwFTouFE+4Hd4G8XC
V6ynsN2CXH039tJl8kxxWyKv+hqZOUt/d+PQ3ZvcJxaMWANEXVOxl/jAOlEaXWjfIDkNfdpvL0uo
8q8JYRgpc3iGq9XG5g4N9cuAWhmf5Ep6rFEiI+QPERf7MGxTLZusM16WpjKU2C2ilKRb/WPJFvlK
kV4iU+JMGId8NId+Kc19/P4ZjmN40zImFfT9iaNFWUyj1MM/5hqqyOEIBzt2Ce5qPdUBERSIxESS
Q1lwl8UQy+RZUZOlQntgOTtmuANES+YtUvQHK9t03GlZP/0SLj/P1/nhHZpHkhqPEtK2H/2rK/PW
G/IODFFPeggXdpGNBTsFoYuO+RB0fgvODalV8rAQI4H3/MEfrEZPxC6laFp3pa9YhcEr0katUKAL
KibViJAkcI4qZFT0UCOkx+3dldiCnkKjLikna3SsovnyFOfF9qe/LNGiP0mKUFZlzOyVWSRWPpWl
vksLp8m/FrQjFdY68oL2wBywFcBpuXoXIcKjN8zE038DPRHgi2hD/15Q1BLt3dCVrKBfFErhOvbu
25VFqn8BMoZOc0dGaQ7xfeBwsb3Rm0DYXKKk8L8/z2jkhZPkerDIjsJhk4h0pYAKXmJzhNtfQQSo
PQBsCrll/xlqp+dxqAGDN0s7Kg1vDLmVLMPrgcoK6pyK/xX6eKpMagmhLeM5JKuamop7CiJEra+b
wLqjmn1EbA/2zpjhSQU/hxlexgTkz922uFjpe81gWAYarq3y1SRGHufBYBwUM+/kmI8sP/GPlopz
90fF642CJEWF/7SeBB65ZEF/6oKPrPXgarItpd4//QWQR+9lT4eNCRLRTpPXAw5MlIi1gW395sM8
Polco5CfEotqVnOtKpT+W1ft8+T+lqV6moeZ8eeI1JlO9sy4kpYzGY0P8wCZzADV/eJcjVO0tpr7
HMO/Epk2q34aW6wc61RPYxTEpEFPKDYe04u7U5+BKpsKmF+M9l7LU/Kd8eozDSf1Ysj803Q0vIef
tfzPBGh/IYRiwEVXvwNgRFo3nscescHUXUUtsdkDA8Cfy9dhE0E6TYSUpaRx3xlCg0bldsF0FKtU
XRZzaiOSJ26OHiTzqTdFu4/fUsYTSgM3MV9kDB9NP0rnMWCiSB1mF8WyjPkyQz4cnyiUtHf4rzR+
KLOpIAgQISSVxLtzmxXW20ZZSjVc9ldufiiJgEN0iIjGeDtykT2jwymH0A8qyDxBpKS1IRhWiidV
wgaezciWIFAyty5Htab+K4HZg8iyHlMvqhCrzW0hWEXZm1K5AQMj+atQDNphVW9lgZ+16FWwk5zc
bACcPJ8HrAkZrcc+oYotzM11612PYYJYEdKCgz7lwP2AINrjnP7kn/FA81E2ybHU+JtUV20ctTvB
f8t/U4jLLaNW2t6SBUInCV9yLLXyJm0cHzFdzSwQUIk/Dg6vMTcMPc4Rt7OFyjE4YU4D6NWkwz6M
IaNfVKwCsxpzLIiHajGBouV9pi/bRvzE4UUhbBgSle0H9Jf4OOfu72vB3CJbRjIbM4olbVmCJ89V
ckZrLSGUNX3aPaDnNQdUjuGej19MzvOBwNqJL01SVXJRaOALugZ3nOadXCuEajrDOgvTVguNZ0Zi
V2ngLVhRFHtQHFre1MOhh99K9Fg+S5esgFH6r7gYQZkZNWARF7zg/xgEY4CJoMZYIOK4dsA8MB/E
eN3ejSV9qWFhAl5Zt9zPNS2dida5LlOdYscSAkm4mxnIBiE+8+QPDhmrw8SW8xl6Lu/98fyKLaX4
QHWCGL7cdu12mbn9eCbldK+7LmXURkte2XP+3R66ntdkFPXS4QqTFrVi9s4R2JIRGSCp61nMIr9P
TecqvD2ZnOoESWRKxWSg1HXAPt/Xn/ptHjbml5OijcepaNcKdoOYopyeDy591zMM8WIf/txM0mhZ
dW3NDz9yDDMzSOmkz1QIYQ+bU2wbGmBbtU4edKrtfCwgLmx2qi2JRF6yT8p9+Fi1HNN3WKiYP7ZQ
sTAV3ooGP/9EoL0n4s/6LAL9caO0S8cqmRibdhTCTuOFum2s+4fnBHiOKx8AmsRHCWiuGr4HxMqb
eUP8sa80+5Smc6LztnWjZmRW2xkCduJQOvV8AuQIb/jS0NMueYLbRE3o4OaH8OFaoQU0X6z5ToEw
O2pqskBCr/wjPWbgpyLlbWDkBDrtfchJXX9Z7CrA9lG1N6A6q3QltOZNKNFgQ5rpPMNHr/hKXTnO
pOKJpYQXAUxBEhLSvesia0MvOjjzZp/VG6RzjtX6gxZQPkgHmQYjGZpgkV7CRsYeaQ2lOwYFcjXN
Zu1qPZnrhhyToo+1N1ycoEl4XjwPmlLzZhPFk8iwXYu/VqPUz6jhAXeyZuYcqOuqLFNo9NMmLy5Y
ABRfQrC51SpWtFfR+WEsohbmEnm+AjSnB1r+IqVbnibYKqEju0itSR6Fr3Lj89bkyHXrM9vgB6UT
lcsizLwy/e4yhFMjw8GuJMfBvcFarrTPBRo+FDgDrwboeIkPuoNMXP6uH+BL8AORZFRTmp2QcnGP
PrIBt0TchVflU0qvbozZ5AYbaFi875gW2DrBLxOzwsSrqhaAlTCdwPoBkSOmwp9HsITyJvGY/T5Q
2rONel4qxQYkY4G/CqjIaaW8DZhP+IjQQjU7uTl+NZUlwBxq0IdoyEDwwx3zrDxvKX5UG8IcLUMx
c7kPYNtAV/yhPf5cB0/0Ads9xOAgBEl15/bKQAikYIn5f1N6JWS1Bw17ALBXSo/7UNd+97fCWnP4
bjBxC8xazn89YEGY6f+dHN0QgnEox1BFaCWlLdGkWbSR7H+BWFuSuCAlHK8ZB4MPq8ptjUOtUoie
DzpRjc50KZsWDgjBfoFLWr2hQDt7OJyQ29fvlGkkQQD+H1yuKGrG34M2stn2yUa15CLkTgodhkJA
TEeVA7hxVOfJTq/aiCoh6xMXJg9vsPBgC/hSOD7qaZGWX9XrYX3xnShbkXgQtMPfvDOWprI5TS6O
do08ZOcG5Jw2aByLuwOfEQIrxC4E18EuNkTh0eATNDYAtJ6ozgwtBupASY/p575jvU9XugBjwcIC
Y/f/eB/CS9ZBDxOb5rNuSSFhj1JT+tqz/Yj4eUbdEqqX7M4TK38QfcUCelzfic0ygLpA6WgDwTHw
XPUNKPJS7BIgQRwdXXIi9rv0l6gKC+kF1pH1+teb793G6SHNX8/AruENKbs3/AgYbDpWneSF3Jxk
M5V07Mmr0DqjEkx+G/ptaUMPIus167qOjCt/DJaxDuCAsylUezSGKzvDqsowyuD1xlZWZUy/i0ds
IWf/Ai6IMT2ywA9MSJ7bUNsjJTC1JlU+3aYWc6fwdGOB0izWKicpMhC3HRJGYzY5QCNWYuXcbfac
w3qBXgYgCb9Y04gg6QhbGgLaXukKMXNmDEQa9zjO0JKee2XK8kdFJrOBy5ZCvgvAbUxEy662daZp
L+rXDgMPJnM/7qDvnosTULf4QzK+KYjG+dm/M4vV2WUzH2dy1Mr+RE1Q7xRCK2kCFAIcSGFgglil
+6GaJBLGF0je7EEYQlbQD6Yiwnu21EnbMrc34cstZlR69VOLMsL3WXl9G66e2PVn3StaLAoWGI4f
rUJf+WN66pva8u00MhHt/T3Inm6Hz+/X6eblXz8EJYNwnQoOQMtat2Lrw2mTXZYHf87L558s3jFR
YugLB3xD9r1EcQteXKfWEfatA/Oz4KIsXQz4/KPvyqmZtVe9BfpxeTRHxua+/OJtqQVWBqdsPcvM
zXyaCCRi5uMg7sbHDRwpeiMgk6oNWUQP7J701ibcK5YiguWO5HMVJ7HcYtFgEGTyK9zxbA6XAT1M
0+2Z+veB9ijJiTjMxFnLSZrDyf/EztZL87WORGDUrkl4yyXAVGfcLBDN+F/PTlT1e9jax33VcSJN
w+e8+6JtMmRhLSaqgHQLjHIgUIEkg8589A8b7FOTkinntX+egKu8QjR2YUZ72X8rjnNO12R4Rmn0
konpMyKAe73lHq3E1YQb9qjGVQyN8f0nHIqLMLEISKWeVKo6xmDcl5pgr6nnYAfd63wGpgppBPzy
8XRJn5+H9VFwSEQzBgbMVTpC1ms4pZFaERxwoysGDMiFuXiA33JAi1l+ZhgSqxeu7wAhbtnYYD1W
jwJ+XvKgBShdrpdNqFXO3kH6Pl135++RzlpKCpSQpYNMkQH9bB/mFkiM2p8HRiwYFOAjuSZujoND
onJQXDLG/fsJ0OcocKwY2Cw+LEa6Q3P6s1Zei8D0Gusz51RcNYASEsRhVXL/q4UFLHXMSA9kCC7j
pnyUs0n46kAPEtBp6ifwIMehiEkPWQagbMdMzAGyCktRf6l1GBMydf30JaKEeusmOGzSaEILebx3
G1LVWgJOMKB0adxpHXxLx+nDTUtAoUVkqW1W2j7HG5n8qbZzlZj2AClxZPvM/FXwPrfDd7ZYU9cl
oVxMMCiJ5hStSNkttJlXEoiOmrLaWUH/torkwoOwZDCon0uRMZWWh1hoNITg6mMvD2wM2gwKwGbF
dfEEpTz00bQT77NNaIycqIrD0Bz0q5z/IKK+z75grbBXQ0aJ8faB7jVoKtY3ENXU0z2Kd5+7I1G9
G80Zi85Exa/V44V4UB6aOpEvD2mJ2ArzWDtwhq5rxWI+tFgPg09kQbGGbglYMoaFkWZ0t9ST5Lwh
JHtt1ZA/2DNzh+sytQTUGdmYWhS/4E/MJxNhob05nANOSM4gHkxbIWch92lc8Y6ta+lvJtwqH5Ko
Ga/ZtY3owCVu9g/uAOJmyUnECjvmPnnsFedFYErxGhE0y4xeGNxoUSBqpkAhYCl/oNu4+POQRHmq
caYy4RDeide2NGSRpFZbGu58veug4gJH0anq1Xsu0rNp1EwatKB7tggvkMTvllmWH5hCmxPW8A7L
Gdl3EyUCmv6mL5cDLP65K6nX62E1p4VjL36ArjJQW6RNTs05QrC+bqVBrVRA4dV6SbdGTvZVLUxK
OXVvRgmxe430lnT06ed0rnS21qhZ7+8MDN9Owv+q0hZHIBaMs7nHCtmRBcHbFNNeZhhg6i7l0S7W
tWiEpHeq8qKclsAp0pkzTXs/6Gfs92irIZ4t1w8+vqU/U18+pqHmURnktDRSxNAmUGL+gu5weglr
6qt3G884mNsQjHcJ0v8kGuYz9mZ4RqDJUv3YS+8mElRYrk4RoV6EctnIjSwpEC2F+/IZZ0hce116
XyVtih2gZ8QTsNyt79rPrqVxbWKUC3oHLEAqbTrO3qEo7igYyCmI+Whoh66AOM1lrZhms6z32jan
h4QRGAAkInApbUixHAJrBqueZfpr49XBaeRTAu8RK1GZydi4QuEwUjARSHjMPubn2dOBdiUzR9Bc
05RJgGTN6N30LdzV2l0TWKFHzlcZW+VXf7A5e8kzsEdsqLTevxOYSNgG9m2tGv+pvNXjcOKj8xZy
170uZDPQyGtrlAkV/kipRcs5Sef7KuPqvVYQmcsFUdpt2Fz2Sb5eQqsErw0ZdtY+KO+MJDBDg33/
EijY7gqj8aCIw8srcUFcNLGvf7GhlTfK7n7veqYbKdupXUE0I9CJhM5chSxuHjp5Pht8LeWQunlG
Q3/1wX8UoFGqogd7/ciyCVLJLTpPdxXd2EFyG13S4YGskQfGa2EL0I5kPrJA7FBh3BTxosCfhTq0
uzeZd8vcwT25YWnpAI8ZufRKG6e7EoqSBHibRgasEbOtyFud5qZdLT6K9L7ORC5+Im2eCYoAZCUa
4gg5HLJFWKPWyaTNq7p7IR+sOUkwnS5Q55pw/j3GpL+clLzxye9X3BeA/ev+tNLcT4BNdZyO3UzR
nAPqp6qvP59Pe30op8TauvuGaafSW1w2gQmeOQ8OPALCWxpytfsi/CR1W4/9lCQdZxUUthTe3zPI
2t0agocEXcO9jn4Kg6/iegJUDP+KztUMYi8GiQb8ipiDFPtXUza9yL4eqR62V68ArwcU4P3PPnLA
qBUpMqyr1qhcXBMSKHkx+S5PY29HonI0F6eUDmjpZ0kVXvPl3Nhg4vLhLy1F1DU0Nh4JMbOtoRQm
SALKIZKtqDof3Xd+8Q7fo3PfAEnpX7PAKSIYPuiuh1F1NcKyOW/HmSc1vy223mr1tRzHZ/lhJJoE
EmSyToh2+PPnvuUqPY3AXrzITqmW/8JaI98cgIQRguNoYioZo6IMj+mkmVk2vouqM7aV1qG+yJVH
8jrM0Bd29sD4RoLsYkerZzmZmWk2cqkogk8rz1GoSnr5jZs6qEsJ9pWwvGDQddVW9KSsY/Dbjuu0
9KGuLzWEZZe5zWaGDzddSZ1b5ScOeBNEtLokHhDf1UTTPFxZ/IEH8C4sDC4O6m4tHk/io21r355h
fprToBvjzp+RfE9D1O2XT+ELmAMlIol1Wpzv6Uj8UcDnT4gzMSktuPAnr8BoYEox1fw1HVMFXTpl
gY1/NVN9AaxErV5if1vhrDKKjO5RWT3+C9rDttkqjPkp9GgXS3Pgvsbcnn7m8C0NvKne87q6d4+a
BnJi0RBEPwt2Zy6ePNAVr5RMnad+Ciyw5ss1vZSelhG7xOv6fBUCyxfOvUgOx+U+xxl18XY6DN2+
peFgoLRfw1EbgP0Q1bNe1SFIskwYxRG4nAs/fwlwrl4w0wgTmN9gOfsQQ5vVw5CUKCZ9hnHsLef6
2FM2tmCktGHhueNGQ9F15Mj8KQE5aEAN31QYfuCr4dxJDp2lLT4jTyYOiOLqbLypN4LRk34UFvv3
dHCRnsXCO6JWi6gf7M0G+YFFcTDbNIvxMVkrk9YMBTlFOjlpaljHcl220HgB+RBjuT6M6bvZ424Y
6bMC3xXmreuBlhZFu6j4mhWipmZ47kePMtXFkuO/wFVIMzEOQLd109FkSPZd6ahLEMs5j0eJ16QL
teJz3K9949mOZt2p9kZapqJKas2MUvyJMGYiO9zWeHEzDJSL6LFB5FibcFOXMIXZQ5h8mYsJ0NzP
mswe/YIrThcPU+5sh/B3kj+zL0FLgreVkszx7ihnnMAKy1o5kC8QAutlIrGQGvmOA+54KWYkx3sR
fYb3Zk2kWxNmErZEIif36/wZMgZDWOpAaMJE7l2DIoGjqh07i8qNTzauup4QKqhPT7wCO7oz+nsf
GLPePE+nepDfoNdIuvzjzWlAZ5LhdtqfNERjo/UNMX2Oyxom/GH+tAmFqvHEiHJt1/nmYDTQ48W3
Avp8k0vI82QtvQq065ZBEs9TyqwxWl74k3Rz8Y71XFX+nEIbIP936d15eS3Wpg7biUl6bbThogEl
WbxJxEMDjztR5dayNyT+TJzBZBnDRdRdfcAwS20X++lOae8k+MPSgBgbjGGHi3MKrMqEtm3lOv/U
d/olxv1hKqIeLHCaH+Vc22lat9znPuygM+Ddl1QGCCcYSuVTUgNBnA3i/FY1tXwyv7/DY+2qGtL9
QRYQCeBnyX3iSE9+12b78BvEGtpB1NqMC4tsqx+oMBtSJ+tP71DiG9Hmt4sgrrk20TsD1zqUcb8B
Zh5MNGuoQvBZCYUqMAvFwPQc3A9KZYJXlbc8nIQtZJK+gdFuItfmKZ6KaxbpnJqILaN9KcHb9ZpI
efgKuT33l5Tj2Da7E9yOLt8mNDmhDB5HnNtNeK2hrUBdAg27T73S5DXvcE3H6i9tUmXtF+nlOreC
ha5SO4H2sOndrwQ6yroJImlYzvnhrB3mNr7tW7kLiTrvQfR1jDSdsXHmgjoHAx9SRvWxdFvMt+FG
WAje3n7EUgXmyoWFoP+7uSjTzKqiPgASMgA7J0OqqHVGlAXZ3mXH/VpmDjojAiTg7I/yjUFjTv6W
DuYf2lMwFWpyR7oIIIldb0tamPY1bYFR2QHBP2WzGzy9Crf5vFuF96l4MV2ggg/+MVTrlfZtkGyU
Rp1ge58c/zSgHvs+iIqo7CnEUf4o4vfDJDAh+5QOytpqH9MKVOffnFDrOu2yhyCpgzIF+laybh5X
pzQeo1ZLUW3t2a0yyVuwDZ0/dyZne7NfKYBsh5h2eDt6py3jNnAf/UHIFn6et8NOdlso4t7s+MVJ
CBUcxosJ2Ps5o2V7OYkJGS5PpGPrtPS9P9jfwE/wPZZD0MuGaisHp840As9tnD+1BUg+0wrxNCYX
eImjw+GgftUhtzS9LbngFHfJADZIsCyUAefbXp69X1I866IM6FVTsQttO15CehhN4zATP/jwlQ8t
tMmrITLaNdzEZaTxdlLMoLfU5qIP/bsqouXvkZ6ntr8iJSDFZH1VlhMpdT4dZtRhSpmIMNR6GuXv
P4wUCg6os9H9wjFpVhqEG6fNxq/68FQsatVBiGxR6RDGRk34mqE0Tr2BjLmUa8UNoU2Em1zwPfs6
hRAGykZPmbygPu1eylgB7apIQ4I2dTYeZgsik0xorGgGheuvNGQ+5xLh6NbOmIqITsp5oBhekaZK
x3FbRrbFqg/1wEBbm7sM9Bq37XlSjRCtRveyagsI5DREb2ydycrrX9SPNvXFq6QAr6sE5SEW99kV
Pn766a7JwCXQ6dj46NEw7O/Ox6x4ucT/i+d+1MC2Azsq8dD7OsUMCh/zfokkqooknVkCpK5VCyQl
N2asJwXUrPr8g3SGx9IWBjSOEKv+TS/jR5hfwlYdo94XMh2hJ/+WuuC6nwE7BknCPF8xQNdEVCTK
LI3C1zgHhLKhKQZrRgVlHeofs9IDN6lQPCGmaASPTcTfrRd+bePbixhWg8Yds63Xl655kzsnDWLT
D+OQpBsDiqfLCN+MlP7xArLUxqT1noYDTgUHkKP/QJtrL8CSjEObsWyOA3J7rVpu+qEvklHosf9b
aM3gOFho8HHA82ByR9FZkwU5hrvilnJQV19CJka77im8kIN1umn+3vIcBZ2gaaSjTUGEvi5UvKbN
kZK0usNl81Ma80ghiI6ukwJlEQyYCZ1oj5YcCsVUo0Fy6Kb0htiTwZ5/6Vk5URumOnuoEc8Z7lAy
UqmFqyIpFBZfvPeT85hwiV1G8n3QrA8OioRCJssmxIOMyo3snBhfVbiXq928NXPhZuG+jref8Ji0
FUuVD5Eu3VfGN1zgOz2/EmIZkLkUMfwUdjJA3uVBY+l9sV1maou2p/IkFZNPbSJ7xCvXyAirYI4q
Fk1u2iitDuNvvKWV1x9ODeUH4+rmAXQMevbUjWfFq6GGuIyYUVeot7V+GB+bNovCEA+2ae9xR3Eu
QsxcEvNALaAEYzsxRD3tVO85ICsKUTF5qemHU5Aq1eMlutrloFi3SWxxsf4MsG+0TVp6OcG0Mf/s
CyRz7QkQGU4PkNQ6+63eoIIb2Lo9tmdqqJ26XXmoEucREkn+sJ6EZJNvp+ERtghO1/WgEQojOpBG
ZZadGiGSqwprxJLgvUMXLdVzYDwL0QyXRJ1npFugzxNmke8y+vQ8FqcqL6TV+ECYPUpxayW/cmb8
l+NlzEdzBYZqga2rwUMfUmzYmaGQwOrodGeZbL8HEBzwCwP9Pv6S6s/PqjHbqJXhU9syw4mw4MnL
4QVfbrTha3+F/shTDAPPPXQCTOzabzhckpVezdmsWGnmtMPVXdGf4Wz3BikHuDGDO4sn1tZmCcKw
C1PM5MocVOgYlh4FDdZCiI1Dan8/kF5kfNLmmJUzjpmbj3JWwIVAaFmEs4gAPKLVy4+B/bW+NwT9
NYPd0Bft/c249Uy+Kl4O9Jf+VS9Xcx+axsBwwsBiOFA2wNEKSMTKIvIo+hO+MmE7VdKge3tta0LU
J6KoqXcGKVd564Fkrv1aUBeCZSxUohhnE0MC6bZ0Sf16AOpmojpEieEBTonz9AKXqIMSYqUiOyYu
Mye5WVeZP7JZYaMts1ucnRQNi/qWsqqZ7ySY+udbZDMy0VIZ7ULuA3rKjtuk0iR7qryZjokCnbug
QHU7Gw/SALIrNQcf9wOrcx4X6SHt9FvhljTK2ntD0UJVe5z5wwWdREdUhlkLcFBJyzLnRZdyN4XP
JDzIXkJbGQNcml+wIKzkI9nHo+5I9JMAayU/evfNjAALjJ7+WWm6UtzoJoHiQKSfLBdslNYA+Xyy
mr+XDVaJ/xcZMGPK7jI62EHrUMbmSezP2BnCLIHQYSgyKp/L9g4ioQoks5OTiCBRt0d0bw8SWjEv
+/WdXnwkuTWTGHo/Ph2p47NYB2KthUxp6xuVfu1CEoXUahsVldJi3SWSvK+d198ty1+8mYuxdWDu
S223LH7pecWh6eup20lvKNICEdDey1Uq71vRn1Wko+M0Zg3XFMFgF1DPxWftiHjABc5gYz3SFBJQ
T4Zx5TsZrJifbQsrHvNvsFaLF1nqj23ojYR9jAkdne9f9UPx8QPRakQGdzPtmYeeQ/KyUhh8xfvL
uLttRrWtoNXJlt1jMX//YwOfaNkxaKfSNV+t1+JBM1WBjANjjTcdJHVABLVmtvCjJARqY1t9A0FU
/K8PMmKKVam8pup/F73o/l3tsbW0EFzDk9eViHBzZ+Fvu7ap0sbaxzSe49/hjklPyfToCK8RvOe6
GYK4Z1wNe1ZKhype8ZtAw5nDgLcuX7cc1tdDbc9cnHQA+/7lBvVdF5yWo2jLUprtxzHp7zWvpHxu
a7g8aCsI7j3tIPp3aKO6dDZeL0W1f2ooy9bURcnapfWUSICLUz1KIU9xQ45gcMfOxvlUCC3Qnyzx
8Ts7Q3Y5+FzCRhXw9rvnXh1EFVR/tmoB6jP/iqM5BkeSpLDpF4bRiWmzFiu+rkavMk67I2xFUX9K
ZfGzYsG9aN3b8hpGVDcvQiGjat6vKfYmvofZ3orqgwTx/zukYwOeOTVwYSFpypV/6cAx/f9XhMtP
GaUB9mgt6xNhpc2R/vGjc9kobReLnSb5pBC5JSU1sM4h4Uk1nBB4p7GQubaqQmYtIZLOvFxWobgx
ZL2OdB46G2Vk1i4KQzUbo4ZuKtal4GL6qsKlOQICRRoLsnhIWXG8FQyDDmZ9LjAfXwr+4CFkbnJa
ziN3xh49PCaRfLyIbG4UE56RWRB/nZZBs3bnCP+BRdTbbU+pg1XE1v5XaBJRdB28kYfr6Sbicb1j
qIYRs5waJt2buCwZm+yd/Co7mEqWCZoEouG42qrHUGyV1CpnCXp6Lx6stMr8Br2k4qoWftCKnVsc
h3y+CYeDUAHl1V0e/pMPLd9KNGz5xndJRlpEQCLepd4BiGsNpcwBk/r/g35ts6DkKdEBfvUpKIwY
RaeBFrK1NA79Hw5X90SdN6IAX7Vbk03b2d3Dm5BMHRZzcfSkmIQDZtv7u/Uc1hRz/q9zQtEemxZc
0jdq0WW9cszQYU5SkntzJSiys7Lr0DHWaXBA81qO5dQggsI2FV7QrWFG9xfWIntVm90wpL+cJdTh
GvW/TkIRm8/8d579pyX0PpLbw/Jw4jxbJYEzWHoJJEHuiV5DtsREL1y9ha9ShzdcyivjZtVvOt4v
KX93L7h0K+Nd6RHQhyb3M06IMaJG8hO354TaloLOEONeBJlGu//teUh8nPW0cJzAqMestPVCp9KA
FPFP2Zmm93fLmKvSyo9qlc54RjoLm7/mcQ0XMsyw6HxG8VOzfBq3vflSMVEm3Ddlycw9r4opcFdy
SYa7Ef2KUNts5st9CBz7rAgCCpLVCNUg7US2xOoTrml4LKrsvj6R+mfZCVEJc7y/ZJB7r8P51XKZ
YQuBeHJLuC6d2gIlg0MRqQOaN+JI8Ya8n+J07Y0g3uBKOuskPrEeY8HSay4yTnYqvWp7bt9SjvE8
cwMLbqMsZ69UmVAK61mQQNqC+BL88CGwmRqxkG+Trgyq3LmDqpzdDEKMQDt6WrwOYFwu/H9i8lih
ek4XmHNxxVOHer7VS+yqWWFYJJFVmUwXJLQf8XBICJzIq8k50Wa4uKKImpzFWe59CxsSdoxx5J3+
EFmR+Hgk6bj+vlLtQUxLdwYyBbbfR7pPCmi7shqneOmzBSjJostQ6Chh2nGsGs1yI834arRisAMc
z8uUFkXOdWmn2l5Qhq50WyoGqiGQH8GZMmz2dZEX2bXtZpiwjtz3wO4ydIy9K2IkDgW8FvqE7pPo
+H5BIaVUfA5s46F3+UxrAf85xdA/A3G9w8BJlC7uV3c70VEwl4p+KP4rb1xHWShaK4WcEM7CXnf9
4/IW84J/YgXHQmJ7z3Su9FA1J74HzVoXR+zIxgPpqW0QYnAh2uYI3SfpU+z7iSyUfJmczEYi3q6g
KPhUZ6IPAr+SBHpTfzxPF0SbKW9ghxE6wVRFwLam2uOGfanK6Q884E1HavCmzM/xtjOp/FuCosNx
yVKcOS5IVwHQwXw3qOeAv8ukKO00ALPzaSLt6NLFf1vN2/eqkGnIAz9SS1QheZv3AzNaLAYk2qAb
WjarbfWB+QS9cpTwSx0aZo4FYhvthfooNiltE+1TUJoIti4xpHz9pMylVKOIbjpfjWiEr6TqtuFU
1F1DVQoglg/55Riav+dlSdvWcDR8fhkzt31z+zm5tyXLM2C3tz4eucDXW0WFQM8ybdFZiZZBnaGG
aYUZNm0/b6lesFu4Xl0irmRbqKoEKJ/DRmtPQuVQZIbEAL9bxvaiWnVf3HUX0FodaNGBW9bP+GaN
cA1GxG2k4gHFQkJvGjnD41Z45OtyugitapRNSSzhzgqx1Ust0RJ4+S591aBh+Wb4txRmRHHWZLl6
UWOJZC7hiCiCaaJbYewuIHb8BqwWgm+TqK2DLBSym0GmUN55L8Zb1XRwgQmM52m/armSGsEJvWRt
wKCV8y+NNWwrfUofrr6RsFMD5DA4yhP7k99uL7qXk9TjtSAtTXzIxKtVzHsXEPjnugt2hnAIVgJQ
rUHan2GZuEhJ73u1sQW2NyGRNsuIwiqV0Mk54t+WIbJX6prn8rkGXFZevRCNSMnP7qYMCHTL9i88
v8Mgz+PfEgMnCq86YX9rYAOf15UOFX53AQP+xByV8QQr64CQPufnFg4+Q7CfsIQEFcfGr4cy8POm
ApFiCxFmPvTJKi6Ni+Wd55RbMGnL5D7It1VUZewS0f5LMJsQF7UzKPp+X+DZ9uSpEr6ODu4IYlzo
5WtnBKD4NEAjdTkm4ToRUneGkfP8l3oEpHOaMYBvjfrODNm90SNAmmSZBHuOGTMuoP2R+IL2eCQN
/Zl28zZc96bSrJlRIx1kqRxwstQnoDeei9s+AwOySdKuI2g3EODgA/0XT/hAoZOkKGECqvmzVyyK
xIdEipUn6A7R+mumt+wTNvSgM66YzYcvs68WP5OxmjME3yX4r704akXnixuWQy5+q6rmwaQVqB54
V/VWRqdbJZ+GMaFsLkpqy8cVf3rkucc3Rih09gNM3abRsNvzrXDJw9rgSlD4S1rr+8MWe3QFNrG0
DwpJXT6gzo7IULr1goZHXh2EbtCc63KXbYSncDaRjGi96KOxXjr+M3SAHzrGofUtEd43n9RQalmE
aQH55VdIHq+kMXQm9SfFSMJ3eKyCq9dbGXNvD+OlOzTCXlUkG8Rvw+HXBG2vnq4P/pn/JbLOD+sx
W7lUEZfkXO452y0Ascku7KKPbbrXbDRY24ZEUzc24yHBGgc6y+U1JmJ9s2MbUrGL0rGMT0juAd4f
qyyEF9HaWV5wtabx4p5XOZ1H+Bw1lvei5UCGx+HKYTHdjGLFNZ9HQ69RMDK1y+Yk0OExNbv9c8CF
XlN9G1agKWxZqB+j+bncD3aqB88Uvar8XVJ/hAly3MyDKgiVJ/N8AYU2VabPkAGPDoAdU6EAdMVO
HveOZLI5WW1gZRT/2Wq+GsFTShqEFMREr3+czWs/htaFy19WhqKDoGgPLYwXg5bYqY4JExnzBhJM
SNtADDKYpGjmS2MfCRihrsN9wBTmvQWknA9QaMmr/y/PNucahFr/DZAI2UYrfIZAsR5eiaG7Zpwv
X5S7v4onfjL0y74yTMXW0CdfZ196IKA+QJ0K732+gFR9tYf7juQIYXJffT2+8RzxW/SMBL+rt05/
CFPBJPxwJmzugZ6hd160wyizXjYk7lJ9JBEKz2Y2qcHebosNN+cjZLpgGPWstL3ilcplLBLvGXiv
qdy/1cu0/L9mKkW683WSHehhmnOVtXkwIN+J/zUh99wUK5dRY6AD4VF5a0W+dnANv8oq5HY6BohI
c+s1qt1ZWo/Pze5L95rk+xGLUk+Rkmj5G8mko4gKr0yBab3LYa3hqM48q42GcIzdlszUDOlEz9P/
VTZZV9yeIBZaH9JQLNDXm/ZFJCwDD/J032ySULMSE4jOELO0aqkQoycTqXNgeO1EbekOi69tkCr0
ThUr/lt2+a2bBjjIwP72Nua3YcSFG5K7ss/06pJk9rWUjpZoAjsMS+0+686RG+a8rDjSrxeEfwgV
ZRGRudZixavRwryzCSb5h9EZ9fL5Xxe5Mfga+kyKC0Vfi6Go8scnuZWq6hMYvZEcMgkqifPNeQFD
7JLeUIHWvYs8soc696pMiAAXUb6ELdAzyE3q846lzNUqwo1qRWKiPwW9HW/ITfht03dVVKQEHqsO
8huWB61m3PDFs6vm/FPatZw2gaYYkl5Y9O0++GIZ3CTH2OTavCsykh4LUCarneP30JqBVGn8s1EL
iSq6jKpsS/D5SqmapBa3xxYKUJRCtbXMhwv5CuGB5mhIEW/fJB08QrB+siQ5xzuMOoIw3ZvdXig1
oPdn4GCLvbbHZaDI9qK9A89cTNTjXlTcXV67L2zjgf028YSrrdiK1qdQhIe1NyZpGwdcI+JUl1Yr
fJdh0ci9s1Lx2TBedm2kFnDMniH/bDPsNfSjwImBK/d97GSR1Ve3Aiux+G8NBjhoclEmvQBUQnp2
fbyHTnNrxfX9cvhgPGOAKykyQuqiuRTrQVXZxhYf5qQCZfJWCgqNgqa2NqlLvTOQdeOqO9OCCOSi
zyZSDrT/xbabOh3K0JpNaGka3wGwrt2QRFUzG5l/vSdm/EUMqA3mA2wS6Ty96Ft+8kTm1mi4j8JH
Z4r5umGOiHBSLuEInZ3CyuWyE7/5CjSCn6/BgFb6TJlAMyX7eUdy/sFRhilBB2tKF9kHu9Fd2+eu
4CkoPu+zeE2i54XTN8uA/LQEcGP62LuJnwNVVHWEqpFxD4HrM5ou7TJSHuGURDeKFMXPAILlIlv+
xJrjrpNxo2qgNECSv+o7w2f6RjKXM+b3ZezQ93QwDcdQR0AMCIqi1APHRjIUcwDIVuur5gisFf5b
+wfIRmEN2vyPYn5zRWssFiBQCi1zRJVTPljyj1nUuDvlpqzDS8BS+oZyc5Nixt9sH41rALdcisRQ
LhEBF0NhkbKhWKiOp0BEMSLzvxh0p+l75zR6aWK0LKs4E55HQVdBhsOccUHm4PgE3ZiclENXnwGV
ePTgCQK+tlUHEfSpa0Cpy6pw79qeXG6sGnqyCpUCAwObrRudnbnID8BI/kDMMbVU1mYtWFj+CwBh
w1fQCxNBWg8db4O6oewndC41rNVmAq5rlsKnJLl1WgufHcXLtveYN8Y4GfKzkS54qzuDfrz1IhMK
hccPcw3j976p26mbOAiq3rSSgxkgV61+FGqVEVQKAyAsaxV3jWX1KLdzb3Lji5txUxshlF66DG7h
GXsyh9oZ/NL/R8Q3SE5sPrTfTNE71M8Y4r2s5G+DTjPpql2lnQHIMnDboZ4DJ7nzAEUsVM8qs1gh
GXBeQJCwQa8rJooezo+jIS66aC7kxLRjuDJodHE0bu++i+iZCI1IJ+FtXA8iiHqFpX2Pd7YQmcHy
C5AnybKyDpbJEkdBUxTtN1dNgSo9nCbSOfQkIl83EwPgGLmYTTiDzTqGNqi6NHISFR8AXUcjnafY
jxU3fSZQsuEI/syLmGbF3vFZus58XXn3WQPsRzoPPqmw+cy4njUI9Gk41tS2aSHby6Hv+wnCpS3V
Cl5a5Bpu/vpXTYUXYtVNvlN/huXFRSuY4JG6SRCL7A3+xXvdo3h65efh4p0g+XmM2Cdp8Co71i/S
e9tLb6jHrq8G/grUmSnvw39VMRmgR1z70He0ItRGFkzacC0vFkkVixZav/SdSjH6j1RZFJAQr18a
xYAcntxvCq0xbWaKR/qT08EGNDabnE6R0IXu9cZhe0xaNSp1L2/YEVAmjLzQB75H4C7nTBikRArM
XtvcuMibysfJUkestDuGeDxj2MHXU03OmN6LciMomLd95Occa4ntVRpCfE4HvrvAOMVRIrDokVse
DsTApumrRJkG4MXcLibRCqBjIJhd/xt/NSKHAX10rv9OJir1j7rkAs8JU5exbSuKLXEJgJNWKDQ6
aaUehIh+34x4GbDEs2L+gsYhOIBXfqwtqss7aLAuXQDRQBrqk956jgm9UWIABpFm33x9FiiQMx8y
9HLw+8QJdgn5y6WcE/k6Y/xA8VTNEYzRZLpNT5vlH0Vx/1b3QKKBVAn0dKN+EBbau6yTJJp10Kd6
+lgzIz0i8J6r8MVKQscEJ0G/6LcMeUNVWFai0lVzVXnrSqeUhoRT2PkpUHWZvZN0fbDu2/tklk/C
ALJOxSu3SojSY3cB/3hkEQqVqx6yrNdr6cBrnDqKRRY0/rp0fWBHVabaMB7XWu9eiI6rqvq04VWk
bKUt5mwS0bA9G2YP9J5XHwNdFBuRvUYQVnYJk0WWFdY6HauuYIv8hfEZtsQwv42CXf8ZCDi2fPKU
w5KpYpQn5RF5mCrw31/OXWJlmJgbHU8IRk5jinCoW36Zc16pxqV3vIHjsJfCCbPOOGEdWlS1++BE
1JJ0RcPUZ3zjBpGSEWeLeUuhBFdGcXk9apL+YJl5b5dVDNkUe+ej/0pGc8romZ8Hd28+MiPfjeOG
+1FUY4wEYg+rSlPoa14o/TEzAVMSwdua2A+6A6MW/93SJdznWRjrO2XXl0tv63f73g2S9EaxL5EF
KgJ0dHEo4Ia0ol4/8IcZDzZhCko3wx71IYH2qyuT4YZ3MCFO2i8qguYQhzb/dc3CmlEf1x7m4EUM
jTNKMnleU9dupHWsPxWa19PQBzD1uapcfjTNzNEbspznvjUpeTHI4UqzJX/klPu9pqPQmyhlIinq
GNj6Mhn3Vn1bwuKrUwUdDwE1y4gYVVwELHnD6xueembz3rWR4X+crqfS0KUnjMjVwANG8nCKcefj
RN6LZzDfB3Qn8199gktCAa0e0e7fGCnGlF8xze814eq+Dc8UswukaIOD1Q7rNRIE4V5bNur8pp9B
BDQr+Rv0FyWgsKUPySeNoKXO8dachR9HjwN3nTC+9mV0HVs0InRZPgQUgPdLJ40AA0s5xQxof37g
0RvvWvq5deyg85EL/0Q5B9sGllQjGkcR3O6JpLNvbigQDbPqIKlOCt0qEJRt5WNzt6JJJAWMrLML
WfLzWyTq1ktoT3F9aCw96eyO2Wj9jNV5Hy8vyUQOCySq+XSmjXKX6P+cgrlp1MaIiz2x/O8vg7HF
5MG9LUQwxAWu4Z9zkvFnKd4jmSdi4se8pUzn7zHBmONhjUaMSds706oIjCbISbGJmc3jYzDIVKIF
RDI2t1aAB5exMu1kKKgskm68p42Xb+oeAqQCui5CsUWkA9rn3aKIsbpm4bMPqq3OTYlHLd5drXZj
Qyux8idZr1+S0VYQIFRCiJIJjaBogPeWUZlGnV5a5egEdqbZ8qNWzK7pQDP+C5kadSrCaDuRx1oz
8WG7NQtSQhi90R7Eml4J1FiPHy2f2izWwDYnfX+UzM7aeZ1xruWIihAtM++2bFWd8/XfzafftLMS
aAWyVZcUeGjYYoMazc6luosauVk+JrAEshN949AkoXMw8QX7kBpdSkQO4Q1DA3gaQJ5FjcclMelk
99C8ZR6S6Oy5PVs+y/VNlJuG42PfHtBu+tbArOC9vrvF+xsFB7Mj+Gc42RvfJFHR563jBcLxFBoI
GJOXgONCRaliY4g9FFWj4b7UzpBomig04oln6njhwfRs/FGZjTcX90f0oaBofEFpwgc4uV5YN8X5
I1BZ4MeFsuMfY2L2/UYCVYlrP6FXlIeL9946pL6rx8zEOtcTcGldnSVf8xXQ7+qZaWJe5gmqUIrx
ba5vBc1oZlQ874NFEQN4Jw/X6ip02jypQBUQBjHA9n0lDQxcGA1mQlDLObnZRAnbQe1EmZGVk1rV
g2LjLt5ratzA0d/I6gyfgghLxE3On/671lMDJsNolcqzBba/h7nuJfMtpiaIBPyEiTScjwDMDtnv
Va++fIPDRpIDxzCDKuqPm8Czj+05JdPB/qjLob5PxIDZAqIt+w7Zh3rRN7dB3Tq8Qt5EbbR7chOe
wH0D/sUyOTazkZyRDqEM9+DUq6Pj9r6c9Iu4ln84Zx9kZcdQ5e3oefFBoyaC864X4I+TIDL+Uf4u
Q2nnZOAV6UblazdA5BpLYg6lMthAGgkIVOb7HcO7yWHOwduTLydpb1hAHZ72DLWsTcD35kbPUYWU
qXGQMQmpt+W7A2vZ5sjA6z3yLWZ08aYMNU2W5z4rVlJu75x2kX73WLd/UNTTt3EJ0HW9ecF6cpFP
UJhcLebfr4IkxgmqxicpYusobVgHXouSzc4QT6gVnAHpgKkt00apeFGxN812twIfLjxLmkv5YQ2l
Y0p0IVkH+YT9PL9A3YpAIz0fXz0O/qHNgUgNcuVya84X7s4ArZM7q207wheS0p/Wa0stDLXzfEeb
a/L7/rD+sbNXCgO0pgYeBjIWZTFElY2vudIrsST2Vvo600F0V4bDwYN/nhb+ohk1D212bxqbVR4h
Weii6XPzuYqB/JliAVm+j0u43IEfv3KkkF0LYLubH0zb7iDy1sgirGZKCCbPhFKfI0wlTOzyXkaP
yVqmoVjwrLHplQmPjhrh0WNRrLenstDiWm+ZGUIWZkfXvlpJcA4cJNDN4cDS2+SDwUkODMePG+FB
yHhbIQinPgsZSyA/X07E3YkJpD+CLNz9of9Y6RwnHAXzdu/ISBozRPYCnVAgvSNh80jebFAiFFhd
VNoJ6UlFpzUjiFdyEkx4nthzMZ32xo8zWYNOacaNMqsZ69H58JmGdZ4/09Xo8WVPVIGuH37/ApbG
giir6gcxAyzW6Hegc22kp3WuVL4PsdLCo5tkXTBoKnxu96+IZxVZ1l+lSBlU5sY8YamPXKCHdwJg
9w6k8WO0lvJpwOuXWIfXemp+MHgAFtGZatRBPjjuUKznNVgun3oRJjwkypAyw6a1KtPoex7q5HH1
E1PjX+RoDxILukRoRLDUKTEoK5o2Y/+8Sm7MWch0aHBl9BFC8WuRGJ3IWCNKVDc5lb+BAwZgPz38
D/462NxQke9uKPqKrD5BDS3+AVlpeZNcU4pdcQfFv/7IcM6vQG+nwE8kr0uYZU+5k0UJqnw142KW
4g/k6N1altOm76uoQ57x9iepRR7W52ZSLObjYfytrA2lwj6s/nVqNDi7aC+5GlCwYLR+Zmjhihfp
/bgo2aNgXi2Pk76onMbEDD8kV7kAsw4jhQ4gV6VCGTqlDbwW36ESLDDIQlqIwJXEH0O1GsdyZ7hD
3bf2+i/kMJuC9fTUKQpgOlX8KIUBv7v/auvIUF/ccPQiK8h1xMOukuLH2JsluA2+talGF1aDDHCW
LCG/OJhu3zaxQK2E+BLvwWilPPr5BWGhLGhBPrG31ePSroICjaVguqdrlIX/+2QUGG24n2Jpy6Js
LN8jd7gCDMCAyLLTCbzEQzVCREKlQsCOif9hxeUjGG8SGvRHoXmTErNG3uVTnYD06uWuB+pTILek
h2u8RxpdDEqaPIyjCEUGjOXhjosXS6LvqXniGNSM+GET83Lpf+hIIeEK/6R/7/LgTP/150h0y1LC
l7lbjRRknTx4FzIhMM7ViFhw9N5PM26PQzb7lGc5YAo38Ip77RQloPaFRy2UnT/nDBcTrOGr4Ck9
r11yZISMsrS67l6lczG1hW9um+018Ww4Hc1eqLIoq8P2jFvzehS1RBz0teD1GuM2QzByQS5jNhNG
mNHU9t2AB5+NkQz2QVC3I5eRoaUbHevJ/9IcZtFH+2jiOdpw7mYfeTw8uj2aY4qscCuaeQaThUg9
w5cYyac788xUpOQVExFt5u1MaBJO0qgV5DAuzpCgA3/gF/z5V0MoGda1VBWTf29cEeZQAy/YQ2rG
v1eaLcFo6FrjF7KUnBuHWkJ3oVsShP827bbATW32UALs29b7nHOBPuWurIJoYuizi0fyNop3l7xz
yA/S6ggVEYI3PIppckEl8UhOB8fXu930MqNVxZulW5dgCQoHT5qGbwR9sEatHZFjm2CZ/65ymeFg
oPX8Ko4uXLlUgJh/Z6P5/uJHyC2xEgUp+9Bpx6P9gLSBlY1N+CjQ/Ic1nuQhlHWsnv0fbER4ggn9
fYNN19HgN2pkZqFGbfJRUkafmueo4ZPn3M8HMdR0Fe73DdkSiQBTbkZq3vxLwMv0BHBwyiJuOlbu
hu+qwLwrrDsi3vvUXGBy7uWIWZ6FDtWGfulEpxVYVeETdgHFWbvaUa6asHuOt0DZ13zpozmTZEz9
Zf2csfaPbI1Am3cbBOeJkIPM+J5tgyGVGZfYecWP68osE0Jj2MAB9+pQK2xmTVAwAq9Z074XqJUC
NoZpXyVXHyQiwSCyNaWsANpdbjRLLKmfkA0pkqLibYNaE+9327jzJOgESUCT1ucdepja4+jr/tKy
ukabfs+dbbBX4fYp0KGZnUREbuqlExH4uPqaQ/E0PjarfvbAmbMqRu2ykuO0NB0gLLKHesn691RO
Zfc98iNtEEa/iPbEZeUtNXWWGWupqHO6l7oOT5Xd+Ic1dE4YJ/tkFp3d15DYXoVb/aVWlbyRA0nX
/mFcs99tcbqtvg8YOmqc79WDuh6qE/ZtOEUVWiWrestgcUONBV6ubQOm/bDaC2vjLQmqsOmlQuZE
FQUhfEN20ezhxAlHipAne8aneBy7YhUkjUzWe3fL4FbO7lT9UWbNxs+runKTZYAt1c3GhoxE1aLY
BzOicGfFTGvHhTyuSjT0l1TsYdCv5wfJMLRRRw4PhctjqnIKClZBNoXo2DDAsY36irFoRXKPizDK
6LUkd4KB1BSHiDfHoXbslw9QVP+QT5th32QHo3SGSLHE1OwKRu5DxRBLy4E++HKxpBJBLQkovH1H
0qBuyU1UXdcTQELxhVRHDk0Gf6CRryd7FVMZkKp7Vl4Lzgyo6MoiQ+aBfgDm1Snr9EtW0GMvNqQZ
7zD7cDUPwC0JMOKiDOOWA/zhiheh44usqs3PKF/3xPmtT2QdVyZ3vPG0lxJsUErO3ZnrMaAuKyW4
ko/EeQmYLhg2Bs1QqEFyCRmqBsl5ybIxrI3rCkp63x/H/Om6zZ2BVfgRcEuCQPZMRfoy9g5r2aIm
ozr0X0PI6Io6zBnCLn0w45i9I1ydqA92+5u4O5PilMLEDyimm1labHxR6sVUK6CnzzLbvNZk9IsQ
n9Imi3kpoN6sVq0kcyTvkveSdp2833uWKMY3LcT6t6kkwpijRxu6SeyOWsoZ0+zdwohMB3+f9TSK
QiTgWT20g/G5/s2WB5SzOJYoMUDTWLtScvY8QwjP5TIEZXJosbJj4OjQI4rpikEBBxu7yJxNfNFz
so9LlfN3LcPwycprtikBraQCRof2JDe+PQuUy5/rmCSREowQ+E9FJuv5f0yAwdcPQVL7J+rAsvFK
mO7gMhCbToSkOHWqF4w9TGhFI3TG19Pvc3zOhq7PEz+SbV+82nv/8XYOO5qQKxnroNhbPP4dJ5C7
y0tqNXXP3E9LWKG1KtHBLXG4OkH3vuaMjZU2PRTLlopZLxiWTJPU0nAxIbxn4Oxz3Qw2S8TINZxW
kX7XFTeypBV69GZvNTHy6AGm6tEeLpv02f1w7Iml23GgihiuA0RrIF1ftQdspc2lTPGtsWBKW8rt
Wa/f36sKB2c/I/t8EMjz9CcYXwAnZweCvGkMtDtntGx4rQx+nPkL1NgUYwe5CdBhHOSrW1KkouYY
kIp9PI/+BkJudWZiDfhZCdL26HRqQwWTVgyRrLJiR9hyQANCTGVuo1khbpCkrZesDwZfCJ9nEhJ1
ML+blkd0xo8neLlFIIgR0KFTmNhoBexz3sYSyltR0isd0D/0AsgQjyeGMkFpXW5R4ixBRsSpn1zh
qtfS5KxB0eeC25MqT7k5Ei0veAazy9pZFbILvOCY3aXgm97r2Xv6lh9J6RJezqh5rNGqtdSZnZYq
u4bMF8yJteeFrQJuvNiBmiuF7UO6x5F8/M47bkgyzMFoz/zK6v4dhBWe2PydVJYm9NL2OhWDzS2a
UawTW7jisa6hPNSjV6cPCh+wZxJ5OLiifXU8thlyQX2/Iapt5GgMvD9q7NxD5LMPOQ37xYprDnB9
IqVcfc6nFuVwqMSqGmxxbjpSw4oTSo1rsETZ4dMWkOqcZgdWqt6UsKysOuwiseqkR4YW++ohqiry
OXRmO95ACraimPUJaXtkeyjeLIERSn5M2iCxz7ZY+oW5JDaOY5QEIjNP6ugWAtX7/NwLP86dMOQh
/xZm3OEcYRnkRfiXzEWMf+akQlHDLlNzhxrvNekegH8B1YSQGocWFrexBUZ8fbzrHD+uhOblJdRG
GE00GweBmG81k/jvSjh9p3GCpXjULghd9jieTi0v3ovC6NmULE50Ut7LG+J9JOYrOFW4PnJGiTk5
uQalRgucYc/mbMqP/PV1m7mKrMTtR+MXWEXcOWeyNc9M/nN3jkYxzTbGAoTO9+n+1hddUK4MsXZ4
HIppp4qdzIVmT5JelMVLhEx53lRn5xcLfdXD79/oCFZ125hgC40eyC/+qSbfOWAZRfrN7adbQCOx
62P7dkD9RRmoJdVYD3UqvXdMawkpNLcBDTSGHboIU3A1DCmqAkT9TpSPjVQ84OigJ5pMHtLRSuMN
p9DZ/cT4WB5af6iDvEqw0Axt/QKZbH18MeyPILeVfiks7HB1x1VriU8ZfAtOmILXZkb2rcQh3viL
ZmhgUJjD3uJ3f1CjnCUUcC+qMbw5/3nBnVjO2cfsuIFScWxMsDTJC2eHoC4tiuz85vL7rZPCl6do
bc+stN9i5jYC6gsaw5Lk8ReIm8utZN3ptKwZO5IY98pVqxp1qc469kTpD5GJmiClW8EtglLBApjx
wVAbqSTbWghpfs++sOMSncQXoQjbIhGtQqoSA0r1IjfwIGu4Z3wu6d7L86+9YM1Mizmx57ZbaDXB
tNeV4S2rQP5UyvH0Bj9KBas1UfDmF5DNflP9Y8tGgCtEfXUl77YwEo/WzuOZO3PfAlEsl2H/CNXz
8PqrDKzEYpNNhCL/E8lODg0bK0FmpHjAHO+BVwUE+m+Y3/rAKUbOCOpIKOTunWZW+TWdq/KBFR1I
VMMIwtVh8jTsKMXXadoB0l13zP2pd8aQs1/rEqyZl8Lq3Bjnt2He2AHx9hNDirRkIQcbqGkwcjVr
GAj+X984pmKyE6VUyXrIUk0iNvNdP7YDOR8NlZz3qL6qgsyZPzisRTnhUosKfoIH3bC0IDsE5v6e
j0xePvUb6FSzH1x8uNCKYQouQmQ7L2LyUQtZ04IonwEMuc7KGgmPhbIvCmJza/HtTuBMLATZWcAw
xH1X8z1O0NI3RiH9PMMgt7QDvOEoXU/1gA3/V/fO4fQJ+39PhYowaS3RZ1+jSJewib+nNr+ya/pa
KL91ayFZnNecxtYwyC3SjNjSYT4Ffz/GI6tf1OhOB29+Ej/iUXf7HfNjTH5GlxqhaROXmX7/kxlr
lTyRH1caq6oz1mqEZtVoPU5tk/QTVGW559+ewi25cRax+3LxC0l1oKjOGyQJQE/vXhStCx4P1WzJ
ORrlbCOorgeKLo1y96KgxTZFsv9c2dp4JsQBVy5A2YUqaztBjvOv8sfI+4/ysQziTAkzz7wPihlo
N/PIuedpv5UmMNwWX3Nr++enJnGeMiGjcoutsyGGtNJnWDdsIxnncN/0wQU5PRHy3wJyreTurL/9
e4sxk/8c7JpSPlilRhdG8rk+T5n0bhr9wY5/DXPHYvxcN8aXOlr91HqdesQPF5i3zsArd22IbGwS
bEEsMCP+bYBfk9QxBJmYGPumvqulqcWT7znuYW8QfvUCbgcGFEMr/s+PGRbdqHIb4fgBVzZHt23y
h561aLyu6hbhW3HQXdcxnVKMvRgfIJ7ys/ibOz5w7jBJhQ8zccVYJIOPorn4Uf+AYa7aHvlfrX26
9RPJYN60pxH0nphM7Pegn+zEPibsbhBc9H7xpKhpkAff7RuzhLSsEt4Vtj6YGQRMUd1VpR94N248
+B0yTUf3QknLLK7EXrTEsMZukOyTxRqyUWbAEIeQJCtIH65/xpl1Xcm5SGlh46DOYWtJaIexcwdM
bw958CoN/QMR4N8ap7zaUOoD0lufb8nsQWidQbAOI+HImPemnZzbTbUzLW6CSnP8gnxLAUp5SAw6
p1yKrX1PNuK0joQmLy8lHapPnk/mvNV/w9323avcudwpXW6rUPKhC5qPUt2W6qyukNZpheHDrDNY
P+N4LoZmtSpeWBAPQLS9vY+OlquHEP0ID3UnTaWMfO8/ddNe1YuxvSY3i7hTD1LVVjSz0Ytugv0u
ONr6+FX0+W8cEOZSv0heI2Irlj/4tqjZ28BJYCdotsFXeX9LHzdOoTM0aLNYDL7NpMvicuwoaMDA
6BTh4B8oCwVY93cnd+A51GjEMfhtVHsjgQ17lSNA65Zc0W0aVNor67whSjFfCaxV8oiaqn5VCV6t
DCzDvxQdvXL+GqJVL3EYl71eiCZr/6BETaAu4UoPWXYOxP4cRJVQexuCddlthtKvU05R2m5bNRn/
g8QK8jTQwEVzFK6tUnzZwsyFyT+YBxZKThwR6c6DZmyZ4U5lvPHGO42bq6547boWBcXcaVS3LNDZ
bbVTEqOH/UnWee7S5LL3eJ5nlg05JvKO/pn5forXqVoVd9ECmvlMbsBAOj/qht+bxAyr22CzfjdG
twyEWjNcNrJ5Rq/SL69N9YPwXJ3lxLi1BbzMQ1ameSledkcUx8R5qQfrqho1lJuYRpjNcBcsI9Nx
9I2ns3mtXpcCf9sxyn1dTTC8s9BRkRam2xsPaQMfBMhFOwB9U/WshbRSWOrRQtORjn6Pld9q0qLF
m8V+SA4XeTY96y09pgKNgPsvtt0u05UwZMS3B1tl6e0vjihT0kV8XGqXWOPAgHfiYIxhukLT0Mxk
Cfm+Jb3/LRNuEoVkATLcqQXZMh0427FkIhYkCbo/prbyBhWnOwtsxQpU01BuFguXU/jggH6cmiM6
UMwUGRk49DEiwRP+yiH2pEb0LYqRjHm12F7WwTgvbvajkrHI6MRPvk+Oys898lhWUmqB5JBSN+o3
t5RlKFy+vxJlXfOkUBMhnFBVgQa+rSpVy7frsJaWdNUemgRaYbsIDF9+G4HYWVDMlVm24WVn6DhJ
bwDogcIivDPMsoag61NgxiD525W8MGPSgDKStlYSlMjB5RKhjh3OX+rwDN/ZJJVDuiL9Rc17HEnB
az1AGEkNLrzyeld0gYt0LRT/iBAGfHj82qv46ikPvBP82euyIxRLzs3n+C7nVAQgK3XTUcWk8tfO
fJvW3nKTh+2/upwmO+Xf7MtBa7baTyiFkzrxJ+XIdlNQeS+lO5jQvVtGmu7mLFQ2ChkioCXG1Z8K
OU/XSABjALlk7DpmQmlGvU1Uk9xk3YvMjw0jpdTOZjkYUDdjhl8wl5T5tAUF44/2ifNCjq31aspm
akxREU8lQYXopHzXgsQwN3ENcS3/9Wa0RbCQBOthuJLrgrbdsJ2P9l0k0LCAdg/JKMSryGNotv9D
a836y/OoX4L4tbPtEPnor3BYOKY2MnssSK31oEpsgkvnxPijrbPKcx3Xia1QtoqzdY6WsktwhRNh
l9mJVComznOKgNKtnGr6N+s3WhxXtpwktcCWw0IzgMtA9p+dN/M5eUyP+NzyQ6nj4fsa8M1gHWne
YKiS2u16o+x3bHL8bSNlRfjugyxXtUvx1kfQ3MRca5X3RyIsV0oCR2uxN99UhtoTqXxY+kuOFXkk
OOQf/Bs2KuVbSZgh6eeaimp25zfk27EWEdovia1o5fmmh/RbTmAD16uq2+LV/llnxQhK5I3noBJS
FQEGJslMsFS3OxgPtKj/8xUFjRmedU75EsFfiQ0CBjCy/d/1BVOAH9mFQx192d89ZUD14oqt+vQI
W30aDlCbET34cdLsr2D0aW1NdOOmXTVvixA5OJtc9eYFpdbez+h4wKqW3yO9Nmgyr6ZTB4JrHSVM
9mQnOcSPS7emkNqBZzsSFybA7fkcRANxE9+zQe9FPDv6SkHtdSrIqfO66CUgfZcX8m5MicA2DNZ6
guZayUsb3V+ajmHpiRXbCq7ICiqw4cXoo8R24Q3Z28g826eI6rkBZGElYpLZsMm0uBO00BE0jgq8
OuvVxYPzre2gOeZs8XF94NJMSdREi56VLKlIq3Dy22IZWznuYXU5D3geXpVIZxZ6n2m7giGbrjmV
yvMaYynwcPTqx7AuDfBAfSG+9U8NdsNcrIfgVu7fM/JdZw9zzEsIk8uB1Iiov0dHeC9X1mucPZLj
3z+ZscQ3tObI34JxK2DdtF0P8zH/FagO6wbFW+VcIt2VxZLS+VzPeS2bbsXYwmzvDUNCNtaV/yP6
tKnbITRvbvebYAMJkvgxluiOyMFVw5XPvyybkRwMZF7j4PzKtleq4BAGuXzWz/VSNHC555f4jj8p
de/feSWgBmp5lLjDwIQ58Go7rBFLfc9X6HBGfb6DS7SWuJnPUOIu75iiN1H3Z2WD9vZ7rn81XTMd
jwsQBoslpoKWHjQ4YTANqKDxRueJBFTZ3PYUWDJ5bPau/jBfj/SBizf9BuFo/lqOFWwlQ/ouVOm1
ZRL+nmlcSKY8K5Jg1Dh9ZeseNv5VfThEIAEaO/81QkS7Py6649idVaHWyW+fx8nFlXEvomRJegLn
zNTIHWjqJbs88V2yKhai29y31r+dWVyMBPICyuAWN7a3TWKBHgJU4VlOyeC1Kq1jEbTC1iqgwfmn
fPzRR7OvuHF10DTYRA+DhZY5c59pfarZCfjjggOhJThftkV3X+GsbhwFtovAfB9MMJuJcBTNSXr1
VMRr7YU+LDpva2t8QO/dn7l3DPlKQRmjYrdeq1mYAoDZiplrl6BbK2y9qb1+CHb9aOfkauZ738Mg
zSRC9/RXC9SQiIi6bMt/kjONPgH3rGx6xH0quX0wfzdnP0Jf6/AoQo0c+jq8VW5FE/82bOKr+Xby
OEMBkOKTYGvRLrr7GSQjtQWuS5OO1wIn/58dNMzkRd8M7JT5B+thKsaudvxgstCfSlufyhIBcG4f
Qt5PVFuIqtRTVoyPRKcgXCk/ZtAIq+FFDnSKaWwdgmZONmbKn2RIxPVLX7wmJjtjyFibQ15JeRst
VPD3/Du29x+yvux/HsK6dKYZbjfoGza9KuFgFIxrr+Hw8F6shVz/lMGmFe7T9/z3aEaoRoK1y3A0
0Bzpx/E6qUcSd5r42qzWh8ztOBCRPKs1cghe5bdyAWbtxDTYLl3P89/1I4L3OTQmuaj31ikZXPKy
6d89uvT145J5ZWEuO8S38yqACpjosCC9/xQGBEny1Buw5B82J84yYhI27EEhUAQmwRAPFT2sP+la
saI9ds6o4una578xzOqcsL8CnQUHpkfYDVV+D64wJMr2KdWwF8IPWiq2Avn0mKJCEONFY9hqRpYU
ZsQjTjdZbQKQmbVrCThgpoNFw/g6fAdOz5DApvlvCxQrXcI3FlG8Hf0WSepnqMtDXsISl3jv5hi/
UgDkhdfiBTnkcElC2P/vHdPzBgwomrYfdIGUX39q7D47m53G8ngGrG4/h/96gTM6dVl2q+mKB8TB
EbqnwV9Z6UugwRLJx56GaWS4YPsC82tI3Ij1wiweFW0eB/loQULJpY5pDKu2eO7lEGt+kppMxjLK
wzUo8YZfOC9jIXFo0eR8mdGiC7Pg2/IwzE84YSmjOFvSKBW5LziWnGrx2kzJlVPWC61qZti6kYC1
vtzQ1E0J+tK6OIKKStbCf3AwcXytfFLlBxN15+lDeohgkCW+A4NGQ5w7uMH3EET+3hPejT0B3Ep1
wbdBO13E1PeDpIobdX8aSoHYWjcBbyz2J+YzCvYbcxz+iMqtgGo31njyszsiPcgvfqAds6e8ZN3N
D9vE9ZV9PrERJBnnOoecbWNgtjT5lDF/LBaF7OS5Zu1J/meM1bu8xnIcbtt0a1jFsPTUAM792d8+
qdH5QFeuw28ZSGkyQSNJSNoC0pdUAeb2pViILIyPZs1ksDxGCrhlQ/CHOT5BYB0XvfLADjx4Vinm
FRveNCQKQudSn3zKn+Xp/BNpuRICn/0MjWVR/4oS09sShGjQPJ8JtpuX3olbbO+ANe4wGEj8s3Vc
Gu2/cHGDt6FnDI6AMRQoQRDqZ/K1G2hDXOqcuoi/jP2xmY/ZSAAuBNVkIb6sr3IBELYtZ91qYpUA
ZRNBuAnxvNyXJOIhFQdxZVLdog2jiMtHreQxQMBaRq/ty1lA4pyb1Nnx983an8wJvBY8XwDACJ1F
tkZ8w6bqeUKFxubNogixES+xiY09fXsvp3o3kDm5s1Hg7bJjfesbySlgGFXmF1Xhjd15PZDy5ZBD
zs2HQaHJZC+PIvd3Li9Hz0QO5/vyb6GbkpB5+eObw5l8HSqinC9CEjbGOffTVeUBeTXfuL1Mo6uW
f/iCCWnk1S7huoyFMMe7wdtVGJuBv3YJCmJbP4A3GHL8kv73qoGdZp6/anEtZa8cDe2B9kaPnMoE
WirYNvAlJysKuXF6dFHU2Ng7b6QIh5gXuLTPX1PcDvlPW6RCbOQsz22n4964k1TqudUnmx56jlVs
baw1K4fDV06vbXvaxquxmdTA7jrX6qfUBd8EMl8nx0bl7nsj1+YoEGySZgbOO0nRSl3yd1aVA7Fo
RuO9XQUy3Vz5WSyG+Uaam/oEQbvlR/oS77z/4ZMjky0hgTjHlli8MR7HDm6JW1zORoso+V+37/YX
NOSjNxaGryaaN7jLYhWBuB4tuti9GAm/WJTw0R3CuKfCdIx1kbjhE4zd2qJiAA24PJzPDiwigjvx
JTzHRAGuy2wVSfyHGvn1auiwUhgqIsSxK2V1Azkj0Xp2ZKD/v83ZF5j3HXrQlaa3fyA6yzN2PMqy
AwNPnUOUBLN1PUyEKOfoAnE2bFJjDpSW2PgAWjlC9p+mJnUIYw5gCl7JuRaXG+3JJJCyqogwbqoQ
hlcMvO2OzCtRU4dh4ccr593M8JywgyKhA98Tzq/rE441xeouF5rYcmINmseBQpUn30rVo6PEG2Al
Z1nDdUUuE0uKhYPMqg2FGS0GAYLFrpxJFFIPZAjv10hP+TUROPHFrUoiW4SbxszBYeqFwXY2GTgR
wBTV6Pzg2l3bj9bD4O4Y0TCkUFUFqWRpTlIZWcq3I0aOnjEZ53kim1tAtMtiBN2YmpIhcx/VwFLh
3mKUXaW6vsWHLaiwWeD2NWA6aoVsG52loH6oYVEdxVW9Y/YUg800lc7UA0AjyOCJjCG0rCyw99jS
TpGPJ+ZhkPwCqAfARRkYLHxEEUDN69OjC53iAJjYGCh1PejdB2jzIOD2t3V+KpNbCQ5OXUhdFoJd
le3CEzwjXwu+FBh+NLNH4stiUO5O8KZPphcYVbtSKV8oRaNRV5YDNhAnbyUMso8pMxpaqG9WMVQa
ouhMJnEJVTpPxiJCliTERoRH3f2egMOuI2IuhQsNodcaAC2CoZFQx6whpnqSdC8Q2cnOIq8/to+V
sVfCafT+46auIeXreJlh+ZEYQT2LIMVLg07RPcylCzcjmJruU2gCHFICkGwJldaFUB67qyCZxSkx
QA4i75+R7+BCoNTrc8hKeAsqpQ2P8XBcrqR1Y2re+ECz8YKYMMU7QENiXqa4Vm8KKKYc6R9e3OXC
hIS6QstXbpEPi+X9gv3TyWFOtTT/EPJlmbY6ScQBbueaVPyyGU+RkekGLZIgpjPRciaAZHabV9Ww
Za8Wog0dqVa8R9YaPgKsjzI1brOTRcQMDG0lscZAyMokaaN/2BNXWYVnCCbqjRRoe+6IlxLazVS8
CUj1r8ZDq4RwLfcD2sOSHsFlpJ3ISrbz/ARixoEtCKRN+SrfraZ+rY7qKr93t9AyQkFXYElYHthF
dYWoGA6u0L4pLuTQFo2Jts9CwGk5M5lpR24dAPTnd8tmWeg1+61pSslaghV1k8jr1pxu6b8492N7
9ZHtoJgzVdc+mgG1XjLqEXLB2miu/2X3enVAdospZgSzKeLj67zJpm5NiTBWJ8vf++JEDzunpmoD
PE4KrqGK468+tAwdLg8i0Es1/0lUCaNH/kJdCzDDf19ZgZmnEXTqcXAVhFQMPv8FDXt0KDoWhyyE
mru/4q/zuuFcJBi+m1k4tzKWGOrwdVP2egzp3PfBrkF5R6aCfLxaM8+5FgbtKejvBuK0KLytWoH2
IBgwMGB3nmGl5E2/jNvzqCHe/7bCSpwUeujymJEqCxIBuEoWxSdsag11LjHwTS8XlP1TIedOXDPP
7I6+Npy58vuVFVnI8bjwKBTFMa2AnBxBUn/tG+GDrq5g9O3rlPtyS23UhMTEwuo95K3zqJdw5KXK
pYNQtQmYnrTO3YCT3heEpThRFYmYZIE+JiCIMZuLpx7g3O5inBxDKJO0A4bEkCh6bztbcCNz7dU7
puSoBmSoOskA2fOV4ibA/x8hN+gM5n7aToKe3ufF4yIFCxFmRKekNDPAhgXdu+RWkFGs27N26KPg
sOCOxZJCyESwbMU4XyBnUDIs4GZWektEwTieP9yrja0hhXuH/34HWdJgMvvAPPLjsi05d1BfbUGw
jh8UMt2aITXVHJE1XuJvMTFkodHrY0Cw5xh9BKiwyPSHaLwCZd8qyKpu/kms8cp0DZwX/pwvj1F9
mr7j4yAvV0ysFo18IMlLI6UyjR35A8wdEKFfn19lFjmkqeAUU3xYaJVwKQWNdZ6yyLo35k16wWMM
y91xA1CNo/1MUxexplzJFh4LNo85IaqprOe9XsbRll3cPPmPEAdY4TQp9qO1rsk75ZV4KG9vhPLD
7d02HBku0N9BOBxGo3U3aguJucmqDelJWM1/ALwCo88+A1jf/91sW91f6zjyOB1ZSQJH+jMmMQEo
sMly0hZHaDJoSKdLMUUOpMJvVxwV3EnvzGHKGbR8xrFeeRzZt4vP721mn/rrx+zjdgdwLY8fTl67
RIVfO6TYeRT6woq+UMSvCutwBh6T7rUeEtEuS2LRDQn9g438DGk1QBv+RhcUYzzvYCLWifvY5jjj
SWh8L9UW5z6jZaojdLiKz9ufZCiiVYm1ocwVIntCK162u2Ewlda3XWJ1ID0yqsSpQAPhpKNset1l
xWU6XGMJI3Da4aIn09ta7ZSafckbKut2d5DDoLAUgWN7wKrCNpM02mQ8Y8i5IfDC1DUfLeeS6EnL
7spVFZIwHn2JpCHClfFYpVypIqyYkeJnR/ST1q+CqRQ9aX1Ue9uayYyvOHXqTzyVKDcqsJ716UJ+
W4BlK0QOtoWVfzDGpzHwcgwXvwBoIqlt6dtlBBdihQEPzXCVkM9dGifXm3FZlWdT2mYuN3rFE8TI
WILWIJum48GR6WKamJeTIB5bCO9h4B2/ZRm9NCLvEK145t6MLQSzTq7GIzyYmmi00jBVyg7I5HL2
N5A73yo9RDc01nsWx5EhbmKaZlWFEKOfPAiI8m77Br33Pr+W1ABCplgDa6q/RR7y91t4MPmi0/yx
N/4d80bQUw6e61/lr5j/70xH2qTy0orpP0i/cW/aW0cGxKOSoYTPjaJuYK5PSF7Al9mfMlRSQUUl
QenRuLyHTNW3mg4/XGnIZJRhQN1D23HUsVRTB+NVLrx+ul6mhXVpquB4EVbLLH2zOS0j2VZUqcQK
mjYZscGbMJhUkz28KP5f1LuMvzGNlQCK1EPaVFN8ZA/nGmZGxZFSqH0vE87uWrUfSIsB3ykkzBm1
Tow72hbi47cbaeIUZnIcGxqoGO6d8/BGxwLCYzrueTYnqHtTIL6irQ1G6/IIqBF4N3iws8dVcd9W
L8fpL/ysqxtjNdRtw97P+95bF94/g2PkF7TzglsG2OKBEygwUtrnpXY2F9WGCdp8X+Pzkc+65UX4
81s2UNO9t8UJ21wIbY4gU5o6Pu0VjgOPLLzZcfcp2ZnVRUYF7Wy1+4CT/lx0DYvc6gaVC7aibfFT
FyOzQkhvOPX7NHIUgIuTrlJSzIbzvk2DEEh2EHe0FIdceHWbP30NyvE+hHTSbM9D4dZ3euTTkRM8
jsqPnhrws+QMSfD0ucuMCeqMDrQ2mtEXM5KeepPUdjmtSK7zS53ZOvy9z6qKe85Yk2BNtlIFvUKw
iHrEjkkykUyV4zqYnaDLmp0WLLFsoHMprJKAuAEKfJYfKc2gLJSw2sxIMZaMmTtCCTl8FkAPIL5A
WMBxvhc8RJlWSkkHIXcKiQ2j1ajk99jJdSmTlozaNvOziC/RW0COvu4/xr2j0NxfoJeWR0Qd/960
aMb+H7RUVeSqFHBRH7Yy+IMxk7uz810ztMcXQKnZnpmUTywj5Rf7K4q0zRlGkrahBydbf3MJkZz/
l3KylFi6r/FdMarIWEeRSsx+vLcyY2R1Gvj9aFHoRPSYb23dq7nvF8z5h3Z/xmrwVRsE6pyERntU
ZpC3Gpm18fVmt6Ccrc6iPN/DLzigHaNZr2hhIarTVuTrddjuvFeRWBbU0FT8U719PWNQGIhyjinC
uTRwfp1FzKPrq8u5cugog4BTYgpiGD5HW4ljil81rJTEgkABD7u6ty9gu5h0w2vk75YjIHCpvRp8
R9/lTfUd39TDCYctg+mrFhA13rPde2q2ovTwwyI4GnpMjdd9rZs0nnKBQt1mJxpvpZsUqzPgxRYT
D5yrKE9Mzhzg/jNZLeZEP89gOcLLxcqSzo/S5lBtiUVaFeX8ihzAGLrsenj0hLAyrOKFUn03PjvE
tH65nVXh9+ulAiQ7MthRo7baRPa19fBUXG4yIgUrTg1ca4bZpbbKMXSeirack8j20Ko/FMlQqpzL
Lzw9rgIUfapQNMaP88jFS8PM/Mk0vUORqXZJ/j7dF3cB+xoku7oL+YwOAaL+eZrE+551BBxkIteI
v/PNq4YnsGQLidVrduywxrEL7Ot+cYhXuyaYNl8S9ZndFaL8sjachZLOulNi77KEL6gX3J/qPcYW
yR5n+6SiewMZb9IAy+Ur4WDF4Uyy4DQcD6Ee8ue8JSlZkKype+U+VHdYocMX0CKVT/dF+qV0Y6v0
JA8lv9kwYkUylLrlJoCWo1nv11uKHcDivCBK2TUBLRO7WOlkpnbdaf3do/GKrOFOG1h0PZGYUZDP
oBPOFonTGGjDvC7Ttd2li7hLgocw4vDdbhJNt1kri4QUBtuv+zhv95AN52MGJpZ4WouVmCB8opoR
uXXcRBN/GaURQToKBGEh2tRxTgec6jnVou8amm7cpHdfUvRPevhjmGEqWkEE4/OULJcgZLGZM0Dw
QFloXJeUZg495SjZy0BOlxn2sGgToS/NCoQ7v8241WeeKYEZi/ixcPo6h/uCpwezMlbJDDvJtMr6
oMUISKPsKPLlIM4O3oufCYwvoPJlLcst65ScZsHyptS/PvLjHKJ3A90n6YfW6J1j3G5kvZSmsSe8
cQzTXpN9dJUqggvFDAliDdHAoIxCvOLQSXpfexl720Awjb3LV4O5Men6Q8fu/5PQpuXZ0JGCyGDL
1cPDARocHlZr8LOYmzkwN0W/Mo5zT8fjuY4uSX3okvKMjHr7HCCTRkOCO+hWwNBDl5MqmOZ5+tiS
UUy8ESqWtqLtcK7BIUaHZqKyU19AY9fGQJVYdxCd5VGhacrVr2c7oE2i4DQtQE+pfgXWGOEI0jPx
la0fY9peO7L6V/z+dCXiTz/laeg/cmRFnPPf9jdvPvxq0dgU64OaOmF9mGMCIeHL02+SDI17oS6C
SNfKl2iHLNjF7lvxMiq1Gf99IHMNI8yYCx4qyHDhIlxIWAy9XEg+Io3Cg8pq/HSi2i2LyINmMJY8
7EE6VnuS6nZO3APQl2dvyZHtAt+7qf/JFrWwWb1FysIcxIj10iyE5NUEqZPXz9WREPS/gxEMD2Vl
tJn4PFPZ0ADEgfic5LS5LO12zAZUVwO0tJhChQ1W1mCAyAdKpdxJBAgBrpNA/hiIGYMVwbVPUydh
/jYI3Bv3tmoOva1N9mdhFQuu7iHYXrnk5RTfabfkwj0f5Ej2J8iCDOgIiukWSYBDa612zA2sib1M
VL44CeSsJGdJk64ZJbj96j4MirL97ivj65JQSGHWC1KtYaVSPV+dsdHb91GZdl7Ppq9l8LKF1S83
I1LcZoEvhKE6a+vlTuZJOlvRh4wMqBaQLNYK3J0YyAfY35n7TqXdHvMOqTYCyt3tXNv77RLaHdAk
tgfI7TZLLdkVF96RjRgrKd6mwVI7rCsgewiZ/I31FXncsYJqu2BPYLAFIqBr2MM4e45LfazeVwTp
oROAFVWuyGgZ99ZdAmmbtuozxfvCM3uovFdV+xQNh/0rfp57uFEa8gIPBqz01ZWz1boNA6/ERXH7
pNJ5wwgptQ16R8Ue2mp2QyfjD9OQYYj5R0DzXjU3ccZ05A38UCawZ+CCp67ojmxVb69StRHVtY5A
HSQ1aPbFpr+s3WgkmvKzuRYV12BeMAIgdv5+BhVTM0/5IIOaPaPF9wCBhuKBXUjyJ3lckymZS2cf
XVTMdd+1aAH1qG4VrlOHUYrUiRP78IcDkLIFcmOXlTb2ji6RCd8B2PZSnaF6PTECz3aCqjfVZAuz
W20pOzEEzttAlomOu1kcvTVECRV5fZran305WhED34sVXlrJEM/3/LGrJvBicVGL1aXlqjv8Vp0d
WPPnuZJ5eJKyXFDDskRWEy4pXD7aBVBoqZZgyxRR7O5lxesHQSvYw6TBMDzZdUah5ER6E+Sp7o5B
/693bqSWL0nPiYhkfPdqI80wR5naEfmEPtKDZbSXyWuTElcfqoZWk3qaGFn23fTBRpAQANzw5L8e
+0wKDAkctTw3o4ka0kk2onv6GIALM35j8NrSm+Lf6fSd4zQbGML0pJwMrvxw1fCSOjwuo3r4Yz8b
n961OR3s9RSWTZV1U+IR4zho3kYZ0rYsR7EuamPhl02nfgzo3AhjQKJstFfBQ4gMd25MJoWab/Nq
KMhj0MChATTUqXwYqVCvvAdZMq0TtB0ccf55kat9eKu7E/ctxgfy7IPh4A2wBUkW6TnwmdWYo1L5
kECAxkI4rfKShRXfIbuef6LOMnKnk9Wzron8vusccYv6N1ozhPy6U9wrGNwAi18HtjVwLM9/5XK8
QHplzKjY+LhJcyXQLvG3GpHhSW12tKG89zfXsENoWyLsFTfLFCF/jQlw6IlyUlir+XcfDJYb044p
X9gO33kUhw+u9kLa0WetsVmVlCPi88b7c7g/jadF7pFRpanGjWV3FvKF5tT3WMDoRBiSOq3jW2cz
2OKQT8vGCgjTIJk6ldcWrEDK+/MrKyFAeF3AOyO5IN9bexfxr669t10sF6uVwomZ2oQCvflCeuIu
QAmrH/+pX/1/mc2Mim3goqDvCXGUdjlFrhpJbRPUgcheWN/sd+Epzn1vNHmCPms6ZaVWWuaiSMGS
wWYk09vzG9ssawAQ/b1CDMro2Xb1s6brG+jEcOddRQzGvIAODSLvjCeFzkJTc9LGMeeJNdf2htTj
PvVmnULgL5ZlzB57eB0HIaH8QVNVDvOK2ZQvayBp/EDF1I2uO9CQtx0B5mX+r9UMmttSgqdviyo/
wrwBYuJVnlr/ReC4VjUPcumv9vdDc1bNI+mjEDdUc0m/te0cXB+wziLuX4MxernqGhb8iF+OF3pS
jiF2Wejjjomu7MsOD6C1hL7Y3GKroMDf3VNglRWzWNV4ACkHGACGLpx3CyySDrGrfFendyN+I1RQ
sksoVBQi7lxr7wDgMpUnv7VzjAZGwNeL3OMfLivZnvVMRuHGiTnb+3tscuI6ldaBmf0yiJTnFcu1
+H1inuijs4sZ39OD08PFkDgoHF9SkJYfr5/bqYo+gvXwWvYtKIxR/EmJgWHX7wKrtnadF8nUcpNb
awGwZc2lkVjz8F3Y0pa264Q20Hxf7zJpESwjViUVXHxG+EweqEcuW5Y93OvuWqhRXmZ7tJGBe4/S
v7l+0F83lxUYcrVIVuC2HYdHSEaREjrtUt0sriW467CEE8uFmxHwUGvAN6bBXqUwezins91oAeYo
3xixI2I8Oto4Asmk5VSyDB81AupNEm7HzAi0Hwk8wEM9lrZUr+GXV9HONywdl+dN8gyNHARjQm+K
llw2u3VC6HnBDs+jMjNUdkJMayz81I1aO6udEJIFCxKO3WgPH8TtDyP4KBpNR5DbQYjArL1VVekI
6BiIAKM4pRelGvBBHegkjCD44Y4ze0LVS9LTaGJEQmku3sg+ZmTbJZicjDN/U8kiW1vJmpRWysVS
VzKkGVw+bvo3PAUixL1GFr+d/0FPLs9JU76xz7tB+wWE6tF7aaZu96fg4cNYt9uqM5xV26+Mn9sp
//YpqCTRDaKXroPkQsYEXyeXByBeW1Lh+76ULss7DSbmRmZxZ9K1ys4CXgktFjtmRdmhSJROvI2l
fY/bcH+gDaMB1tHuaGvlf1dlDsjTrm1v6I68+tl4BqITT8COTl1v1Acl8au9JKOyJlrwfPBwL07R
jKOB5XY14A0hs2fLUP81FXxAt3UrFx9WnnpnnCilfPHvMq0F0Pm90P9azENovoAMLtjIrXk0mOSx
DmJWrsiEkJ2LOgOKTmskuaqgVeCW9MrALcbVcHf3rqFVYx+xK/ooiPSXm5GhJ+9O54tmDvmpZgC7
1CSG9nRnplcrX8bLN1UTvMooKfydAEfFyTDcLxdB7vg4S3DNEpLNmzY9SkSP1pVlTVlaq+v8zUMm
6A8meEX5Toj5YBnHH4OQySZ+y3yQKHQYIIGs7iFbL/5HJWO2x846JcDHh+fmp0Diks0s/WNgebsv
54KLeQwOK3PWHEAC0okRXVrloL7QidEKFPnu1vAvRe1CwCqp55K3UsJHH57xkJrorzX5KCt/yl65
HwJuVmMOYw/fSDmKCdO7jCZf9pDPmAk/YPD+vFjZt0nxkBjdDCiwNiC3rm+qE51GWzbcV3CTmV/s
oFmgJPoUPDbILR99g5jVLNI+PTFwgxfP2JsYD6dzBZJj11XTlpfziNCoEbj/TJn2DhjAkhuK9t8U
eTot3NF2YGnY+11TuJyOOiyERS2uxltHO47aQsRHVxszjQYYDytoupsFI1B5f4OQfzKGaJVAQ8VW
m6jYA/Jn4ixCT2r12L67e0XVVZOmjLyt0+8PaDFi04hCo2oluRYxmo7T6hdIC2Hbd64K6HSKDZeA
i/emgZTahBz8mIg7j2hUE0qbv2ojxRRnVvMIuf2fXvS5aEzac8TCetPVXHdunW7SwQsxwXOTrX94
runaf6TgyVZi//4IinyqNv5mm1a58yTXLr/GqMQ3mPRVWSgS8sQj9BZBMWw4F1bLDmMomLIcp+xJ
TLAtJOfIQ1wGnwHUQcRci9Jg8X17WCl2tkCw8FUO+mzGQApSeIw9voAxQD6GqzrpOnyDLMGabHw0
EMF5vdMYsO1vy4A79Z6fo9imHpHOynDnxg5QOKd518IZFhJ9xS+mF7IfKOy76O6eseCexPYDpKrT
xAoiB+X8QEqTttIIYaM+Pwh1e1ZLWD6Wua7voVdGH8V/lf7rQzT8X+fcoVh5erJK6De5aM7Zj5St
9kinaoFIiLZqe4K6XXJggopt0uWVc4dSR1yDoSUb8ilJ6qKwtRTjlLRVLpg1PPBeZp0u1GdO88XX
1f8mB+qozWodsnguywRE9HaxfJ0WDPzIgA6VT+Q/KPEiY82IOGebAf4UTe5j6AG6h74oKGFCJR89
R43u+HX8Ee/om+mF8mbkaqeIHPNH7MCzf37lxcNofNBSh+Grkkpq6eBmItddh4b4/eOftREqeT8B
mtscq3skF7LcNyOw07X/E+9cYH1+1RU3HsRtIuh2sGBBzvwfpfZrNrlBpmO/T6lLUnSwW69leUWQ
Y0lql4tNhrXXhHukAnP0mKocisMwLillRf6pEr6cR8SNp508a0oVzEXHSLpJ3LCJPPpD2fQJsRPk
yG1LiJru6qj8SivonlFlW3pkZ700sBjgF4QCFI5Xd8JsbUnpq0R+fkDsV1diQhpOUvIGPqq44sFu
6HKhR6Z9YRCbmQBm/wqUiT6PI7S0eZVz/LWTt33hs98a15cnb9HYH2tgMktYfo2jR+XKjCi8FxtE
HiZRHXbHGyRpFKOTF0JJAdbHQv/CrQXxr1ri3v0hOZ/ZSn0nhLCj03s5wZJe8HJiINeHnUgeqLiz
xs6w1s2q8m9QD2+fadSDg+3zB6Uqrnm5xrHbDftzIHgSW6Zm3i0MnWCbMg4EcFWh2ljZcK/+YLmS
rflR8yJD+17/xe36Qt7esRMnLBsrKYpt2YS/+xxJhpyTO4Cp9ZTiJlJdRFPICFcBKCLyTjD7fNe1
G/HIKGTAvwzztqxnpPU1y7j/27YM/QgTLPto9txw5jffX13jbznkSVvX9Fa7Yxz/iuOQsavTMcgA
Q+oUHMuwVdvOSvwZ2EbVsfFGqov9+6rGOmi+YB0uR/b7Ze2vkxWJN6RNWoLqmrLSpsv7UG1XCDHJ
YdwcjgciPiCj2isbiZBSWIFb6b0Xn2ofWgWsj40zW6eWGJSLQqEz/jfWHVn6dks7j7VtZ+BWXeOy
1q2JPC8cgK1+aKboPPaWwkmpd5AjZ53kkAf5Cd3c9e7XPyBGQZzo31uGTPWqV8IknPR9cISKZX8i
s+iPTqWChIYW+7ObxDK+Q8PZVy8Bf5EDfoVwWWZK8Myf4aHs9q8OCZ0KsaxgJcIBEc44Mf+FDRN5
9d0FYxXwqEhrAsVD1Wfee2LhjUWgo1Gr63BLlqtIew2nGY7vw4VXR1FU3KU81EIsmrBizmNE9Fqp
7Xo+f+7HJY5W/maXkXlLuEcO1Nys5od451Ee7S8HlenUOSPfI3d0jt6S0ryEJ6Gh/gJ2LtWb2Pns
+ViXB5Lo80i4dqFT0INzLGqr6+A2M8e2onJN5u1V+9dn91xZTOzmp1mWmVBHmmGR9KmJnTqP+928
hrblXnBuMxda/a6jzjprdz3GNuxPmkl3IQQv24R5KNIUcOY7seNzhZM4eXhIzhK9n4PJCn62/pc5
cideTFBUqxNPzkq+WOq64spWbOlvpxDlEaWj9ehg2VR1G+FXjSxcQsk8V9F0LNqGz0FsuKbLhj7x
/qOlTNfougXKNmurpcCajqWBf5SV7czFnaU7C3SfksOVdA2AnqRh/zFS4R1gbLwfcRBowb+7kQNT
uGdwFcHgWE3PdyCl89Gwmx0HUhNTMfTfBJLxsra7k6TaiGPVprhmqISonopU9i4qL843Jfe1ZmUI
kLHrIhL99aXEsN4iRg8yYate70sx8qrn/XT4k/BIARJXLuOlNZ34eC8zb0nYy856aflgtdiY4OKe
HJShCvD76lfR/GInMseFZQsL2OChA5/KC8kloQsBbqM0LqusJv9o4TgKHYYmQCz+yXSYUrMxmIe7
sQQSgtDgb3ifOoDrBnM1uXh9f/xmVMMuVw1WqhV4/TT4bI7RmVfpkjZGPeaj/JZTnC4AXBFWtP9H
szg530xPhWTpRSKQFi5LWf1j5LG2KD/ZHCNrpplqE+ZZnpKoCiSW262YyBecf4P1OrTB5IGK8SoT
ly6jJQtget25RzHboWOjZH6p297UTM/X4qTbNtMDi/Q2862gLaxqTl/oRW/fCvwKiDUQ+jm/f0Xz
5u8LPR6ZgU2QR+TjL14T9FmagmuviwdRGc2NihJ0ZXHbkJ4ZaceOfuAhVSUd5ovRCXIlw7m6H8fg
L0FwOT70MVhchN2Ft3hPdp6EfERT1DEkKJmUN+DM6lqBQBfs5ZiexpYZGbOG2OmpceTETadtIuZn
hJwRQyVGaifstAE4i5djbtvXfM67HYUpNjCtQY/D2gLvVvcgT8Vcbwptvg5kO2vC+KKlf2xjt7LX
FaTqOmU1ePEndQMnW43EIRMaEODZpV5pXohiRyKDsYSmAW2RyEhfBkNo2Gw1AZ/DcWuiNykKt1FB
fJUQOGiZkr1rU9YnXtiD68kzE34169UxFpL7GTEQYTjEmesI28SqwmyPY9oqdmsAhMaisuCrEvxL
Up1l8KFx0Uck9ea330mGpUr0i8KzuhpcEVd6Zmac/Gj2qhafV7Ge8ZkCTAyenaUqP8NRRiVU8h2I
0DwX4vQPCHGZ8ZsBk8wH8//rbcPm7CktMMvpxCEZV0PNeMMzXuv3UvfzDhcPCIVvi6RwBtjzPamU
cWumlrT2swmU2oezX/WeGFyXEGYPvsuyzxi9FmEY0oLa3e3laDlhasolUw8XziEUB4fyWIV8g1v8
GCKQNIS72eBcsLBMPU31DtRHz+J2YqXA0XRuMImqykLJyWqrAXrcouV/D10Gic3wr3Y85vFeG8S7
TgQqUlaCn8jGUSYsNSaH6GE3dPs4QGXmmVJOX/IRY9QmGs5M7tSbjVQmJzWYBFBNL8WmQCggy+ol
tCUBj2216RZc7tDsPUcXroWYerl7iBT7mEFSho4x6sExCJgo17/3CiE+XrSjcDSc8ZGV5wAtHvfG
4ZG0i8fF+5PcFzE26JIEtGi2baOAb44mFwlEj0ZAUl3Kzd5dCd0hqqVGcnD+pdkeeWiSlPjavCVG
y/rKmyE58e/NDlOZvXny4AbzRfhuend22bGOD98qHZHQpDYoTqurrHMxx+7xs1NKBLjFrLGlbxsT
WeuuIpNXv6LdLfrNJS3IY4qqvcJ1wgpfPd2rwidlYrala6tQPyViF3iy/CJn7iDx+aORAkIUl1VX
qcqf+y79+83bJIIFGNT77ZIkC1w/1P/n0BxEz/vGo4/pAHdwOuDQfDfktkf3gJUJ8shjKm4Cpnc/
qP0ZsZ1CgWt2ic/hggnqFbxmiv0rHMtlz5NSkNPiIWwF9MWQbN0gT6sGE836ri6XvQTq1nSR8sot
W7UydPlK6K71BLCr7sq75dpH90rCrAOf5R8kylIRFOZVMJMfGh8oGNoKVZ9vOFyJzT5tmq67MT1g
4l/mobs+0cQFI0OODmcUTBqgA3AfYPFXSC+7K8FYSoKESqm8nonJbdom50oGzKb9SKSOhqfYUBGl
Iifawsv57nEfYiO22b7YkeqCnDGHHOhwFnVaIJDmK64C27PnVd0VbyAp7/1gHDs2F7xNRmnBLUm5
CkXRerEfO9S4HVhgA8uUeu0TjOjzev3VDkVoo6mWlPSUSWGVm8L/a/wMy2UVIYXE383FNo2OIu5k
BJNH4iwf4ToCXfBotJIc7gnlia/azBAqD5en5+plCbz1w41CLuR2GTXyu1lpSyBmj+KBd4Fce5NZ
vTlQPFav+4HpJxfLAPLUbBmox/57CzDqogxgw+hHigVFy3puRnaTtuzS8NX+wWYdOL4FVVGKq4Ci
ZJzX+VYaI2MuBiSm72GHY7NUutRXjV2hgq7fcJ1tBQTZn0Bmt08rya1+GwO3TFPpNfQHQ1LHJ5Pj
BsGL5zRJOdjpHMNu9LRzk7MnDPaNIizPezr2l5Ci82FfMmmYHCqoEVup8z7MIS+SwAGkLhJLytCs
obOPckOF7tblyBC3f2JEnCj4P4nv6+MGJ32xss3zkqKaX95Zsac5XE6PwM/Y2Uz6laHV+/11igSQ
1eOTHFtde7czLdwqX84+yNHmxR8ZxNfd/INxsmgmm7TtnaWMkRfxDFiui/A2vFyUPGfblQwWZU+R
B2v3Ip1nkaxIxGVoa7VjC+IfZASJHa/TZBw/8T0jYYlOWC6os1/zPDkyqZjRli+ovGhx7f7yXFaY
drSGl9TWMU+q1DXqefQonYdSDWQ2bFcGTTTI/kHdaxweIe0zbQGToB6XUl9u6iNIemvPAOjwY7df
8bXdkuYE9EMXS6Ojnkq5jb/qKjj5HBPFRLUPdubOUvVlmtr1dLfxy3Tk75jmW00rYSNvbLg6ZLET
sYhYKO0oyh69aw+6W+ONskRTpqUTwtegFs+CsFpwPfDBh8zz+ZR3gcybJTZB1dA7spdV8fDK4eSc
D23q6FaZXvggulBkJgJFLeCXaLO3TvxdYMd/84HofGqJS5s29+NJI5fGMMGJPsBSU76+oHFtNFrv
ZQJuzqRPatyHDpS4eFOO5IZBb97ZzdsyyZ/7myMaawXgYbsK3Xg9qs3oKW33WnOv23O9+lntUEhk
TwOvmdrvPHi7niat9ZtIasgkZ67dT9ehY2cGS9LMVAbVTOcIxfaY4j17hmpgk2abCGBJUt0076lg
r9AQnqeo/POaO6/ahB/bkiVB8QLKxRoHhb8E5PTJYTQLhpS3/lTrKH6+R33RIKEiJ1KEcLXhg+Ov
dweMAeYaeYEE5/nZjigtzv2G4TZmdJxEnkTaxmKQArmTf+oxqY1UEyhd+bILrz7HaZW5QoNUmhMz
kpYoUzolmM9fB/EJZTDJqhA1qaDslf4Pi679gLR6xGoXnJ1wqS/gEdRtDx2fn8FeCNLvOafrnDuW
nv277WapvbQaovEypw6KvOTVGIT2xhZTEqvb1K8uTLK2uQe3fN4hRvvWCqH2oofCyHBDj98dgIAQ
rwzrRGB92YTf5MKhAsKnGB4wtvVqaKExR98gBVsRlyb6FLWVQq3hO1Msqcbma6zKlFAflJJypeN7
RaX4q/N2wQK9j7VraBPtfwTgMbPG0a305dU9pF4W+mw7pe1t2O6BCxJdeIxrewinZg+aMV06uDL6
eAWlHqlv6FqX21ofO5PPefR3EaKOljsqUeE8rh1OloMJ1Vl4pkQvc3pk8rdoVQ4RUqW3qiuq2QA5
NQIH/iJjEIf5FlmOg9w+uS0PAbfDg/mK1T7Pa86RnoMk5tzKU7SgbfH/jy2SC+vnNOxrBT8+eOJS
7Ye2P4Miy0j1wSHvXIT+o/g0AMGzwLOgnLKenwSWIZ7G9iIh08dSuMtU6dKCeZwRcD7H6lgoVXEc
j3MBrutGtsH6VqlzMzh/0bQDieDlzX7fuJZGF04J3138toA8EKT2tBPG+BzWCAa9viKO5NPdMKtd
QNGxpgB2emwclsiNJ21HRnjEQiEBoXp/a76o5WgAbD4dyYS5AUHJc7kjkmCPnyF+bG3LkyGmIFFL
1T5GlMdrEgH22/NuXdIclBZoGg/nGL+9HgV5M0Qn5QvPHOg/Wn7jIDh7e0M2/UMB90Um6XVKjtHA
Cj+aGzjWVdMUDZ/4zqiTxzPoHYG+tkWrbxg9qYmpPN+6Xo3/DqdFSLEPdANNC6zSwOJHqPXo2/t6
toEIQNAlJ2E8CBPU8O7HTjGmjbOwggmrIlyiahJAV/91QmzMJeg/sp8NwKAG3hKR0w8b38JqtOY7
JZ/TXJQFkxEpOUFi0S3EQeysG0iiMQBRpx1k8OiWL4CddRVnObUOX3J5CYzUKAXbaSdIGuAERFg3
fsR4aB4IJxKGlMxbLwfFuI08kb7q7XV1/dpXkiiZ0rwHSXhVeaDDmFmr5iaRT2hKy4ALZLLwUuiG
CuwLA0spchqtttqJEw10fh4huGKFBYEkISLT/1+Gq7q90osp1Ag/FXOqMAktVQ40MPgw1qcSwH0y
oHMDWboxtEcjz7Hqf8rMYAMpEC5f9/By5DS9KP1UcbIIb1Kd+i4paszD2W2ib6sgXMhrEpBFAt+f
/hODhwckC6sXF1x6da8KyO45kBP/+JO3/TMxcapTXMNnp/gPIMhWj4ePWS6W+ctZxob9FSOwoPp5
6elTSPQD/ZbVLxXFP3USPy21Tw65HVOGe0TH0580LzNgmdTUC0EFCSlOvKSzzY2azvk/IR11VpY2
q1v5o6apMiIJF234sBNN89iMO8NCXuKZyzDi0PdXohDoEB7GxoY2IOjCtPEqDc5otbKthuz3ludw
Z4tT2dxGVKUda0VStWYxX6fhAgInPQdPLgxV4q/OMLZ+oUwytWNWZqY9G61JG5sE7l4+/I8XfV/p
G68w0U9nqPU3R8H1jDFVPj+4vZ89vxjGAdAjMVD+kOQpkCSiMrrpZZl9PJVg3S3KaoFKuyNqVZKw
+VivCbASasVxFQ/n3nFxhD86vR/2HpMvn+zwMPx8QynlOdcU9fnswfU+QrzEdNaUPGu1Ro1o1p7N
kgM66RHewhCM7TIPJTn03GC0u0XoBJ32iNSEYNvBqmB2NLXI5++ydfGxHvmubgvArSeQuhYOJ28D
Vw7z7nSWeVSrTnwPehnjuWm21nJ8g7Cbk6Ff/Kiur1DLx1uaCPZ3y5Fb7VVStycVBuSPLk0glncG
OuHFunqR2LtjrU9BK56RKq2zFIb47qmNzk/Jt5/qMG8l+ULuUyFe9cw5a0Hi8OpXIgCIIk7LMbiq
/u+Qr6Sw6VXu2DlTmrJIq+ePt6ySoqwSZKRv1jGWzvpvonJFZAWCujE/foCqVp6VV1OodrBE7U+5
m3tEiKOedQSc43m/rwmevIG36/YI5bbwr/W4XBgb/XYhY476qiYdefj9ZmLHAPm7rp+IFRfS7Fa9
VlHhzVhlIuUzDr1CacMuD6vj3G0e7nKLiCkIfOohhup/g7RR8io+pG0AqYfLWpADiK1nP6toOWx6
9mz2DPvRkzemknJMViUWpu7qb7eoJnYmdPMR9KuMNIyuD9em6N9OFRf++WDp85v+YIviUG8el9W/
8+9R0ycVGLclFrlc7KX8ooXL32km8S0fXhCj7NBd/ZF74J4IvTtQgSYpRlCFg49nR+k/TYSxg1hI
DYJh9Xuti6zbwDWmiaj9jSu5anlFBOKuBX/Ekx++C5/TV5L42Ae0af54BAkxbcTnIWWbzOCWlMSN
HdNcRqc4ip2BGD9siN7sUQzOlsj3CGyvxtkmfWFmhSMT5goQDOxmUl4o4Pmu3QlelHmQOQeAmfqX
KDZPEvJofXDuPsR7WjvYlKdTy96e1SUnUzYUOsFQ+S5tY5d3EAaJoVzLmumi1PM70skMTHgp7BkU
lssU6jvaJFHhtxMXVlW36LrpuAlrSTx1GqH/38GjKNhWgz+nTp3ofY9CoL7zC/7U5NFB/K3PPIWW
hR3sPuigNV+OwoECPNzNfN9I/V3Gqz93yRbR8pFPdsmxii4uC/DEFvUxPntrcMg3krNFEkDeEa6U
PSHg5JnXgJJgjGGQNnvsYIVUtVVgmycj+8w+ijzvZsaeWSwM/KIzoH+4FDYGFpUd8tVvYT07Dzde
olqSLBFRysQBnS5dgFEYWmAqQDdM6DeSXa0U6zJufk0Q3y5soOY+AG5I3xFpUq/TJjJlTkGtqBic
GjKyYcG1U059Hx6fjiMDw7ULWBU5LUKNaCKMsZ1iqTHCNTScdrEoUDotnWcuiawp8TWt0fYUKKER
wxa+t2GP3v2n82NKt+FeTlxAbigIz/8eagL2CD79M9/y61vTSn5AnutXlBEdRkCfVOKPrOx9VF8T
9mgmUECCrChXLlB6zzD9rR282aprXX0stpKVUA6GYBin9Fy/9IdoiuqpLQogV0XsLiP9KXSnyi4K
qRL11351V2Uh+8UM3PumV7WeiLn2srVUJ/mLI2xL8BN3n4MYw6G244xaPTUVa69KR3/QIpXQcvbB
FJ9MSlvvEN2Rc4UgqVZTGu3PizPSOvTTpd9flp1u8ngzAfcR2mDpFA7DomLuGa3jTE55BWKV8SVi
LwHqhjVSk9/N4WQheLZinq3l5ygyLhb13JZ88KG7KA+C1lFkyEpydtD33XoFUCwv/6wNAD1K3wjX
TiLZ3GdLAKztWE8A7O7vN/7LUwsEu3a16HTYlelrgsMX+0p9Y1FIhH7nEe4HW39Is+8TGTnRnaJi
nQAt5Cp0tBaASQ0uLSLCDDKQYcKQctvq+72lq+U2kK3oQEA1LkCEala/xxMRU103VhTU12VFyBh1
1HhChz7x1pzsLw1fkjddr5cH1t5N8CLWdhcuRCYAh+gFvG1snonPJpnUcgNe0XW05il5FuO6okNG
p5gVAQ1laAHox4mb72GrfjuFXpRQNMdTzeCVH4FNmxrArDo4JsJEHfd9yLPP+1MW1LR7YwgtCIRK
RhOiQJUq4PlfNcT43YKMezuSwXOE+ExfTKIHfI5/njPXLjaPKm3/vjIaXxp6riIcS8bc4WCGO9z6
F667/3MyWoyBgRVG4D3qKepYab/9i0xtmgnBA2ytsdIRzWq19gl5+5M1mxvSjXL02sciakYgc4SL
tQCNyCr6B2n085ilUKziLI4MssF03TeetfNXgolVBly/GeA6znBQ6eLgeFujaq+Q3ZdRVJmxHmfL
LUCunhD8HA8BFf36troF5bPGausxfWJuU9ZeAlFr1ddEo/y2Do5cFgnA+lePippJ8nF+nHmRjTkR
b7rs65feqvlksFYZ1K9HUUt7e19hwrkbNxc9sSLsuS6vWgMMYjhdCXij95bTEAhDsq4YrCIQlrxs
eUffG+vr5e28R8al4Ke/APn4I+6SERDS8FJN84NSKX8X1uOxTIn3Jp93pGD14AoaD5LnT5cg4ZVd
kLyBBztBpLyEnTQGwbR5SeZ9Li15U123xjsgUST63biDtSGh+8hkOF4eOAsXlNWUpyvlRJriUMAw
y0LSjxbBT+p6MZe7OoWqT6Ay5YvxwgL8X/aYPCJ9BVtMqTz0FEySJinZjQN2sk7VLqxKCjq9Osc1
Tw3MPYh4mo8RC0XNIo+p1um/dKUj72PueFKqOKctkXRtiJug7ZxhdrQOTN1lIxjjbL58fQ6JD34v
gzZbMsRvFWWlcCjynV6KQjFB/u+HCl87vMpNcDhLgE3mzqmBb9qHoBBaB+urImGJz/DLrMvDfuww
/lU3CiK2Hbraee+2ZBc1xVPnBRpn2uThMBmrGzGZthHcT8M695PPi4Td3EKKcDO1aGjfGLlaEid+
UlrAx1SGvade984c8WfCE94ubH9+Srtn10lq8dlVDpftymr22/lPTq0QPwiUQMuX81UXz8VOwLpL
YIJbRQ9ua1OhtEE+wbs8B8qTTxVM/IgUFVcnPKcG2JcWkiVbUtAYpdqL9/udVgN9XOV/MWu5LqKL
trBxKNGyTU/txauTVP3Jm3gt/a+WlQm3y6H095XMsY/SKeOlyONuIqZ2kiMnSTGEoxyRByObK/0+
vj1q5AU3yzgaHpDxnxL9Yno0fVRPNT06ISzch1COFmPD/TWquzeocOkq8nujSnPEI2Tb81Hu1j2a
7nG+u3j6PVrhCR35pFaAzhOE0nEoKy/bknFs+frAkMOWt5q6SMCgjzqAd7a93AbUOpBkhazjAv3G
+jbGS1G35DyfJDg9f3m7w1N6nosvpqza7gLCB75l3F/c9r4hXPlyLOrSsHhNOBNCb8vy/q0GNQtj
cB0EW6veyIgwOdehPKLio7GwbvBcl0DC5/+dl3pP3Zs1TogSbaoD17xVzXqrf1tMG8OjTG49QCsH
af5PMWOvr9XwWKxrRS1qSUWjjaG2Q2xhoy/6jVcQWnQS62nd0pKfgX5Dkuf89RShpg6ihIoKhIys
3q4H2MThbtKwVx+MF7LVcc2i6TyJ+vsj3d7pcniwkEKEXtgTWGEqkyLFXq3Y4iP+PcgMQpmTeEDh
LI2fPGtzgGFz41FNZR3Mf928f/ljbUpM6wZiiQkJ4avRorKwR4aYKjHp740K7kyEzgVIAm2CboKA
ISldV+qny6Dh2cogDpko93EvMEGevzTAkyOLPWMGvKvuwho2Y+ty/wn3VkTpdQUyAaLJJ+dRxEA+
R4mxqVIz1voBdkN3eVwZWgUEVb2isS9gGO7VOYVvKJK2RHwNOHDy+gIbvuc9JqUeQKA2i2B3/7PA
boTuvJbm0zjhbQhdBDgjP6o03+Rc/IUJtVfGeNHT4nCGU/XGQMV7030sgCwLI1wj+O4fy4G8OqxT
8ElnHzZNAIlNuVQuYZtZ3Wvz24RIYZxSLMvfAI8h2pXMoyom2lfMvPeH9Ix+WPWXZiQxJzceK60o
OEeDgCu1JBY6GPp8p37oQ+f5bLyxKNt9+IiRMVkMvPI6gcMprQdzKFtvKgFTPIG2/sga3+fAJyLZ
WZGFDp/s0tFQMAEQRbA6jDt0EAy2hoOWkN0HuuI1ntXql6RhjZP0do5KppjyPn5BdUhYW3Ap6wHM
0RekOFAG9m1YdjyGTjG/lHNsurj2eHtqrBSxwpocUn/EFcnqbe1bnJSxJKFrLRHUlPRh18zpIl84
NOxoC02etrGUwjnRrcGpP5HkaAIcvvWbbb7HAzZEfRdemLCnAVz5dgrzZ7YKl3SGrfO69iYlXWmE
tOMOKeE3wZL9k6sW+ouZb+KT1MswR90o2s5p4xUdDfFKtEGgJdm9vZFU1DEArZEE8lTIZt5Nio5a
hMgIjJNsf/qloAkvcHFqCF+eGclis3NSyBoObVkNMQma9CqVF5hPeprxvCVUsGqv96LKHLGZm03s
NPjS8j/dIjj2Gt5h/KpfBcXGKZ7TldNTfbVvzDhB0ub8u515XudtAsH2r1c0xU95hxYI/XGbLz8I
UAAYDQuedaI26OnBMZ0Y6YoztssxmG+dzezmeAKgQK2Qd73v1izrsCY2nlmZ5D6C9HkEvh4v38lU
be7Q165FDUCrsu0qnp/zE5BUrUQa6g3d8Nlqk8JiGbJ0nrsh8nxJzY7ByZyxaMlrRnvntvVToe+b
Wd/vQCbWjb5PUiTpC+xIYhgkhc5mp/c/QRKpA1qgfx4x9iZaEic9ZnH/YuMmVFVE8EPTvL5fPCyX
AfiWDZYTrk2tju05o0FwCeYZbNLCpP8MVILudcyT0p/z/d4llj7LNpcSa2p4iAZdy8YSFecDp3Rf
LBF38BI+hXQHizTaghvyjj+NXpgulfyUW/Neznoya6c4wfbyvPVft8+iZxY0YKJ7Z1bnD56khETZ
NsxMrfFl8EwEvBrfot9XNwqjRnXhqLE5LMPltBGq8c1oGa8HdAjeBEFUcXObNVIAU1h3JayibEAz
IarCumvx5AcZNHSpIjmnD8ALJjWdm1JNTZcepIayLOv+piQhAXBIsCBqiPE0Rxl0DSlVje64i+X1
K2XIVRnJvyCXNK1Y7klZO3YesqfmRzF9tH9sCV4TWrNdTTNEjk98xY62vSSktavCtzSvtwcfC9cm
rDCLGdHEncjphBZsQ9h5CMYODT9Ik8a5MKKgaW5z+ZDMJqG3+RA8aKiv/iHVd6yDDcvTcTkbUqlJ
U2AThsc4btIKF/MTOD01jm8IvorpEnDev8qWjle/EYBX3VG97olB46F5VMKdP3qQUKeU8PGaC90h
dHjpmlOO1lA8i/w6GxPfMo8/Msi8QQaGTY7cYyeNasrmAf3zb6VCVOTdlFqZuLxzF+8KNbF7RPqJ
96rvHW+Dbu3kO83g6GRwcWnCkfTXtitQpc8ZA2uZGDeiFdun0vuPL/1i1UqUFjK5vJXBKIxvHkBE
YE2VPUatZGhD66fIT+aXNr2f1FRMmP6g0rheZvs6ws1DPC4URB2f/qdN4ev4Xt+DlN93TEAKOLRW
JDPbM1dcnBzofUH/2k+5EUnDkO7jLdyZ04Li8uCxYoI+Xv9WAiTJY1cgmD9kOpAIcbtJPSTAAkSy
3Rtuq4A/3SKUQsip3eUOEw6sTrfs8vVa13jC2h74B3/xXdTdtznY7Ap7UC/TiYKV2ycfsFR1teqL
FS3r4cefI210hVFW0R149w90Gs7Ssxhq3P5MQH1LKJGmb8cyG/MI5LPUAGcMQbU9C4oRMY8HoQ5G
jmHFpaKl6vFIrA1Avnbg3kLUn97k8Ug0NvS53pg0xVuHiAVP4QJ9tKFd+4Rx5El5a4HzMRNKax2U
p7CzC4E6C8sywdzrhCQbF45M+sFVkmczbBJZAvVFwtAx+9tsPr0iIFGnftqA6mTTkbBv1fM+fjqi
E4nkT2YeWYO0lj4wkrk342qSc2DVORZt2Nji8WOtiJxxpJFQvNYsPUUQy4G+eGg8L/YNmqF+Ph+6
f3nfWoFDOAwaW7c2T1SpxJrUtM+NYy4OSY3BJnTehweFsUXfgKSLEnwIzUUxGcwXl+sqKoS9Xb9p
R+T7CY5RPSft2vIiBlbu+GWdsSyLbibcT7eXTCdQvfo9+nlSUgw4Gq+t32/gOPO4mzh1gN83kInL
1fgO1luSfNOIuunSV6vknqAEq2Kyh2AVschBGZj9/ONFd28cVXdl7NbW2lEMYwPqpst9kien6m1X
IdiSneHxLflMy05jycgKSHbzELkRNBNDW1LGD+/w1Uft/dohpFwJL+4tS0eYRsXLPI4Ii+mqNGXI
ZyOkRdmwv16rJwY8UBovA2S6s1NzrdbIrIWhc1++JDLzQbyRA0Ty/EoINqRjqX0oYDMeAGhHGaef
GeqL/LCcB2wJ0hD/BR9RN7JgsdJXZF9u40OxtWmbqQqdKDM3VK7JY83DEWgXSlIvCD15o1ByE8Pc
Y8ykkRSF3axJGuJnyjcXBb51ioqk9uPuBdn515tID4md43caEA3k/aqvBCOK8YyZUBj2m5Szs7Ra
6Uxdr8ur9VW4vD1YDmJPqymqHVmxHpIsIRjnZkbg6YehriKL5ytiHT/N/rwjdxAwgMljj8Zqr+Jb
zSLLxFpUPoyKsVT59Aw1KLNEDNUjq7n0pB0YrVBHYOY3T8+6tKqkkJtNAWWrlzy9EfIaaymlGtFJ
M7CDCDFqNUh8DB0le/7tQZsw/kkT0XGukV6MAyC2fYdpsUA2+hWwVOPO0q7fFENOp5DMTYUM49Ao
evOKlRRXguTQbCAVE6S+ZKI9PVR4U2W7z7OLOan8wUseFHTccwuM/O0mCBRJEJa4sJOFj99Qi9bn
L/Zn8lhBTUCbBRZOeJqIdwb7mpDQplIzTt5kgsuiSd09s/y+MT9kPrc0TkKgx9CinlGB3h4MmKBz
AofgfHDAFf6fiUhZa3RT2v2ldnBHMLxlXvaate4C+TEAbvHNDDv0mm1AaMz6lTJKmgD36BA8Us24
W2XtYv7Vxpvr6zsmkdDfTxkox67jIH+wk0VUKmzUrqt7pA/lJ3ihH9+7sobIFncGVV+iXt+FUOcd
FnblRwQV7+jAIEjdNeeuPvCRx5b5FGM7BOOG89T9drVxoFlMYzX1VHQKxIMoEVDo/PKWLrVW05tA
heOCNzANVZvrT8aAW2cGmUCaGp3axX7G04+/BrLZbNxDze4rqkkgjJ5WrtaEIXRbWO2GOPwU8sy2
pdg8LwiXlyKL/OvUieG1w+NE4R5uPOg7IvMR7yjWKbsA7EY6AzU2s+Qt4njdr+O0dM5obLcLbKc9
pJlTVdtDDmPqWbNFqCm54qg0hYllz2ix/ODQW9jWtXaIOXOdVstzfBX4au+UJXestAkKYwA0uCGZ
lVX4hX0UM3gDIbNmMbw/opB4kXWINxWVG2G5NtehifW/YZaWQw41BWvvCdHbVkF3D0dkNiss4V5X
WYbxLwN1sD1AYokDcsQ7R+WD5zErZB/Ftu10pbxWfy3uIgffT6I324BZJtKXeRBiazXWCwJT5YX9
eIkwanZulYlSL52rdjVDO0AADhgAAHArqR5cTcwgk1mwlgjuxcIxdNiBuOFYFIT/aXNWe22nmHx+
JXEmcw3deOcW+9ODEIdQFujqh8o4jqi1WhcZJNWrL767e2DNu8c3DjUu0NmxQdS6Q0yYFh0H+2Ms
XfsdiHfhCqW2TJCNgXEmzoN6reWWG9GXEzd4ILT9cx/Jl2LyO4vp5iLc14i/jyfBd1HUsx/Aiko+
2hpgBVeTrT5R8gdmYfMxH+QfEl2YiyzwDP72qvublFA6+Yu+EKCo3w2BOulr9ln9nr3+tl7PdzjR
EoZrssdrGmgJRuUtvJO5/PtFZhb038SPK5Msm4QEr8pXuqhZOMvRtN/BkjuIrn+ywhKG/CNq4t/x
AzZoQTZJPCusVAMpPDA8/EwZ85mG3azCeFcI9g/K/QoMAspaDz5jVzyVxqPsB7Iut5QekEUyseOB
D3m130jKB5i5Gp0Mo1Nk1QCJrgLjLOAvnBCHESHMg5kRpVHYb0sZqhjP5OtuqvwZIf6Ka6nAsGYY
W9HlR0k5Vm3ivi+KGSAjEzyrprE4cj6he1ZdcWAD+SunH525Ytj55ayt8NN6enchIffE0Lhe3fIT
x6bKl2c9dOY1LmqC8/58DxFPyk8kOHj++bqr0VPKlwUBp5f+VvcrhakfnRW4X9riTJ335Jyz/9St
Q0Hxmalm6bobGsDSgRO/9Rjm8T1HNB3RkCH3y0F+9WrJZgCLU0xsx2ViSVEwr86qmGXGCTAg8WkM
0tlWAnbPvyKX/2L2XxsKtFz2EYhHKvuHr4mgGeDGKN4OLhHfdjf+DNE4WNZS7sl9Mxh3e22+WuV0
P+0p3TTeSoc0/z4j6vQ+OTm/I7b8OsvqIIAGgRNI0++qRCPGLrjOHitnn24UWsxjOWc3P9sYuP3g
sykRrpH4Vdbso8m83O+AuO1WGkEu4zZxxst7/kAmyzUw7GWtOz6/XKGyp1+WJLU2mo997Rp+vcdc
h0/m9zlcendfbyOVf+7q8j0bnY+ft8fCKkDikz+obp57MmlLddUPOTFehkfjTYLoh28qX67Mf22B
vO17wG5YDlKgGqDEQHzmP4y7M1IONiak7mCY5Mh5LnTaK2xfoc0EwTJ6ALOWI5a+nCQMHBXPYCEd
24eds9k665DNFQLa7Wc6bbIZ5XM1wJRoLRcYj2KG8FBDLM7+ZrIGnFodJBVK5ah/c2UVsQEW/Y6B
GmNaOdZmZQHVkI2bMdIkOUWl7SHoqKJD8naYSjtVdgBNiuIZypgpuRhrfVAnA8JsFDoqIxyfgtfU
uzO2xi0dnhnFOR5LeclbVHqJvHoEMnVVXF1UVkHBHaHJL6+6CTQiTokpoVz9r/1r8a9zRlOXTYXf
s4j5u3iMDrrxwIzE+BDo7Qj5rf4AZ6UeDXm+DgdLQt/+59d21C1aqKB3xYjRrSjCsr1yo26K24EO
oclXhmQUgaXFTSJo3UbGTD5fHzAiTCGlIoUhXXebukZCW58roDx9d2FJbsvD/0sHnQxykwRity+B
Rvk8dM/LMCuaAHYkdFIyGXCVna+7Uhyx5NCi/1n8rzQXI+bPeIHU3E9CFb1dq/pmUcDUGM0cZTf+
rdabFHJYNQgws2aM42Q1VG/fXYljz+EmFuAMqS/Whi32FrGfIWFRwOrrDj2VHzoTV9gIsemari8U
+GhWxqyYwb/pkCG8+JigAj4p2b6CdDFmEV5CIbwXGQ346f6q3pew6u3WPXwMmTfuO8uekVA1ZPP0
r+MROmN7JR26x8/vdtlTC9gZJE6Y7kAhi9+I/uCOgoJhwiFSZ7Yu8+7qc/7zJMMM2+Q4LinvP4kv
vr15964Kvv0LLogLoRO9M4mSPdNiwTgKc4jC+N3gYWvTzrUUPwlH6Q0KYBP2SSSNhPozw714IusP
7doTG73asDc9pDRiXfS6BXJU069wet7RjHBdKRCz6vakmxuBhb/so9DgoLAdw8LaS4wHgPCQV6k0
gZTOOAXDLVVunTAF7j5AqNyVYvgKTWPN8nuc72Zr1fUFA+5OUa5HHvmKMr5DIPiLithaFlV+myGD
3kibSp/47x0mXk7MQ9sKDUOoH8j5cy6lr0FVfWkla/c9QO8AJmuRrVWjFAdz23RsdbCx9Npli+Gt
cJUGLGKMHArIpUQtlyhe58j3ILF2vMBIe/6hRmpTrFpO5pngGzchbNrH6RXVMShUnsMiXaCdVrSG
4Lp1K0kWhQeAwxF3GITXIxl8mEDKOD/RkDWKM1m8mZzyDGM8+rPs2I9fJEsoLdNnTh4dqCrXhaUE
vagKJbhG14u58EarIqfr0dZDGHuUvmP/hT3R9k09oSMkRe0DViO93lilBMC7hfS4cW/7lpqgsz90
IJM47Q1WlSBn/7ywpOWA70SwA/qXcFRNMQaVRxYEqUHGjAtEnY69gBGYFibYml7fh4LXRh5PBymZ
vJfjzd4uSRBXqFIEHoOkA2P0oJmbgVfX9cH4nM7JQHSStK7HKnsvjFIydDg8agJdRMlnQXwbC4CG
ojygOmNbZXKCeRLYRGg4X1kMpKOXxDC1ISO/CWW0jSDExpx95X/NASKzyusngMrCth42Is07U9GN
Al72yoiKLafG2cbp99XbXCzf314rz6vL0zfEJ7khWIYAxKHwZvhc6/aZOMqAOLo8czJGWUnMOMh8
nS+rHo+0g/jegLjmKTl/Wsx47aL465G7v3iB8mKCgVWJJLuP2REIWE5y2O2laOzWUZG3gM5mXZs7
FshOFEMyBb6D8aYqN5UKlV2D/gzK+qcwfSh64b5HFgxp89vUAL+ZR1Ns61PswHN72XRy3lOFdaG4
Jh+pXNs67tfKegB4n49xpP2hqyPz8v1TF8YlqA1UBtUTYuzZFjZwqeYSHVAMPN2O5kLtDkm1bzP1
QofhWsTJut46w6hGhJNBJPrl/h9vYtyW7XUUEbzrZBpTtla90IW0aTZKew4kWBmXttScX/hrom/g
YSakofFM0zAnfEkWcqHg7EM3tIWvGcjrGGZxKq77YyM/W91JOiMnWaEm4mo/qgmTb0h3b+VnPWwL
dLLGFXANI8aKKz0vVrzYQdb8wP8ccqEt/9FJo3H09fsAQSWEbd9RwqVgZR0s41IzO5xdGesuo31d
AqpctWuFGILA93wjg6JeiiT0ZoWcsfXVDEnqnz+MimWv4GW3knFMeIeycMSqFeYCePrBhvhk0vWT
tH98LuzPiiSJpy0jU8dtPPDacLyPmHgMHsQZRweg/UEwpIlnrSAq7fUpZ70rwlO+QkjrwcsWPhFi
Lfa7eRDL6EjkRXolqeISaoJ/Dm1Lo1IAptngYfCmlaw/s7MF1pRUl298QnasB2qFwFm+I9MxpliM
xmk4zajA01Y5F8b7MN4IOyA8Xcp0+OuhJh8/yCHxP7ZgG3xdPP3WUBykXgJwmBpkfjYXmMUjSY/l
c3mi3FTnQUkguzCUdSSEqq6aqt38p6t+SeHk4lx3DCHyq+A059V7HnEflfMD4Dpn8nr0inOwrIed
c51DOJj0RyZref2Fv81W1xKDmx5f2/kJb6yj/t8yVFDLfutIo5BM+ZPPxWc3IUj2xZ0tYrOnPjxL
v6zYoKwb6GhRmGDDSOFr5BkIVI5T+lTTa9KKq0HdjnMA+THjhvD7y7Hf3CykwuI1NyLSb0H7pVkV
nckdPNAJYRUnZlM0gzHytCR1ZFADZSuPlrjokUMBUPrICzG/p2u1sqR9cdLxHbtuED5gFHASQsWC
+9/xfSuKeSSvswacp1Yq8ve5yFv3NMOrkgDKWekjc8dISPS3K5M/RXU1deiNhSq+PEZJnaCHuIxw
cHam/Opv0B7AX3MiX2dYn1T+rvdnDauyfbGZ0lzs5t3Slz0yzEC18y3K5urAOKterDFItMhf8hM2
kvNKsj2TM7FSvZlF7UmJv6rRxgi29/TlScKU3+XJYYBZDFbwFBIhlJ+T4jStBgj36rLbwnvzraFL
DyJ4DKEFnZhjDOIr75T8CqUi5wURmPPhdBa0sWrYaWsJYGf1PqeoJoXbuLKV4Tv5yycBZVJNbJ0P
NyHmU4B2f/8GRqD/klv0IYCpxG0BicIwnUmDGkXbGcAvtrZzRbFYh/B6VNhYIzqr8tDDDXtvmSls
NIKErf8Rv80DV2OHJYpec1FOkfTRYkfYzZn9TwielhzHB1oAis7geSfCkbxBA9OixWG2PtVmQ0C+
3XJjlRHi6roz5Ew6gqi0jzc1ikUcXV7HDKekg/9IXmjJkVzLEBltyug00rfOVGpqbphdfHX8M6ws
/h2PWYr9xS22oDt4Auy5NXS97dKrJKCBA6u1hwyGrhOS4xxXMNvPuvz/lqumdKAURqa09g/LXrI2
D0wfYIqAXbpO/T6eorvO08MF6tyMcUqNJwz3skzrK4R39t+7OGEP7Ey8afhUSZ55gzK5sKoQ8ptp
goqEjTc2wtkNC9S1RU76BFrKvlXzvstDU5aiiJwrYf2M8++wfk+Ox0AYvtz/88C9r6qi+ODlszva
MuWbf1k6r+tw8BipYQaLd1W2UNdNDOkkoAVfeX4hAzOX3Zo4GI77psY5gk179G9YVDltQUFJh8Bj
SRu002+YHwQNhE5X7IQhPlQh2vR3q+M4x4q00fsvLSBEtYmGFQDbyK0EdysWHEY3S91/H3p07+Uy
aQDjTBvLBHZj/DfwVLN9ikGgxNLgRf4BU4GgGc6T/TvVdbifODBz8qpLssLXMixjrHvXxGBom6VA
Yr8dtRF3/OFd67FtRx6eQtw9jcyFemZdpTD9ux4YKsixl2m/5dSyMKQ0F1nOtSGK/6ZSvru5gUiE
21sbGAKJLf+OTEpHkNrpuwLfGYMD0gJYh4ZUOa7GBp06cbUfGKMD4CoNqYf3rR2uLMnGNxE7YEAM
AIEz8FFO/ej6pPliI7IvwA7DpNTfG8Z31IxCbrBOOFwTLKsjen7o/M5lg+mw4oDuUAlYK+mP+74E
qoMJ9rU3nMY/t5hmb86aX5L4d75qdx//59ZiLxhshTpvj8gA2q2yMmtPT26vG1gErnB48BoqxKSB
feJ5WJu2oqTQc5Ey8J0E8EAfstAbWlR2yGJMPABb1rFJZpA5zlOKOHMjfSOw/cnSm4Q6WZabJGja
GrnSz01ZE/qogUt4CsexA76nTPDXhwLVYBhGSsWknAd6hiU1csfndWiQ9QXR2ScV0aOtb2ktukS3
rWDWpHeXKiPIZuFvYqo1jHDnmRGn+iqamgQ6yYfz4X0A2eUd7rlQN6vA4FeYepf0xJBRa0AbFdmp
A/2Ad09rwiJNb8rkGg2PZSjns6nhz8eNylcmiEqpEPLV7zkeyU1jbLKzfQXjA51V9XgAySEUtIfn
mc3eo7nCtEMV1AWi3L7hU11I5TeDNFD2gnz6qWdbRgS/6fr1ci2yjdLCbQbCQOWM/bdDcDsR36Qo
7IIbDuFiBfpbBdn1CAfW05PGdjMDRlyThm2rct0nSeqVSY9y2/RnjrQsFcqp+T/YKluzYWmR8prh
1No3x6cYPoTfX0xBgPKDCTRXNTcwawTY4qOgH//riJCPuLWKXWuN+u14nSvuwtCY2yJnGzbFrwsg
qj6aL0+wWw77Wp4w1NsM1cuMT2IsAdOO+v9ovW+vwzYH+D/XK8q1ghgEfE8B/0iIXpzShcZfoIjR
G1kfNw1Whpq2UwlAdQJuvYNu7yEWTjpp+uwdGK5p/QoJFK9dyA51ZcYJzxc+LFi2tdZMN0A3TviK
qJen7TAtS0Bn9iltvvwvVLQmOAGYpgrfs3C6M3vwbyFhVu/NYGqIZs/Kn48xGM3ribYzNECu9Vsr
3i4SnevT4CMPbBCkSETAATmygMsf10bSoSHq5PpTf4mRoXqebR6H/uRqxfcB4vtULsD0RDr4DVhj
EHlCq/tEn3ZUgf/02ceFdtC6hSKBVWbRWsbVb5vbF39RR0tGu68o5+j6xi4sUu2JWbPs7rHawovo
LEoq/SpBMXvwrcWTrWwu2BuEssxMhqkVYZLeNSYVLQXFMe1Y6Uok+F5blKpf8ZR8OvoG8o4kGJ4t
AUdyBzaDudYekOBfZnqzEbuECGvGWR+HsvndcsLLSUWyZLsIwTL7a2ygciKiwEXY8irB2Vo1QdjX
WXMSUDGwSEXAsqwGqA7fxv8CqM1cSeFOPt78UAeX/Ul8Onl17+87oJRRCx/PkSDBAAwcRAT0xs92
7f7cYWC/SOWflLOOUaAYPK5UcSJkBL+6n1ihS4UnOtNRJ4YOuLj/AKuPd7tqkqXvQFiygGtQiVjl
jQBom7QR6+gCA9LgZrV7VrBDiL9PYxOCMC5oa5jaET0CrrJD59bWxKnT1LyEPusAJLE31N1ZvWeC
/lIX+0NJ9SdvIOq9LgZSmr7qZmAwqv43KwYdhR6xdLAIbtmCbi9NCDHUyCp3/XCvr1FPR2+VPdxd
jC8AUvARlr1WgJ36UF6cKhRQg6lyD2zZDxzC8JbwRgG31aoNZTz/DxXACefDgQAJiGnUBjcAxcuC
w2dnLY1PWSfo6llQwmHwqj73a3BIr6MSbuxxfq1HIhRv5b6gwhIHFBTBvSem39mWBd3hT9WUdOJP
9DhVADojWDZc4tYX4tlLlg37iV3iaL5RBksKxy2e0XDw+ngTbPAGEz0cbUzqDFjxb3iqNa4hOYYW
oZ3UxrZ2i369QpIDX3c+rj/u2Wc4HrHzC0SsTNr6R4kWjVmsWMwRLwy89VAnqRkZwv9J/UnJqvHU
XdvuOQxT3W3EAGlphTdunQCKC4K9omq+NYjrsB/HJey9+naqBoSnpdNVShMmbvpl7An8XgfTxtsv
8BwWWLjjau10y4dJR7WEHprIykZH8Sw0u0k4T/NQdGponC12Bk3DYm/h506keZ7DTH4iLXflWGWH
QAFOA1ru4AHATNFqbJPulb2UKZaz8z+HWrZ0osREjOGI2UlzH0RcpXNZTJL58ZS68fqGvGIDv0AO
HRXEDiBcNTY6fAOv7mTDB0DuFoGJIAjMCuEtq6X0tdsQ6r85s5nf+SDj2AX6w9Fhu6CQEIjVdIeV
JXFYXtfK4OCCvjYQruaS0h0xPZQYIM2NrTJRuj5Rj6wzB+07mHdjFwyU/KS3GBzWQnxT59cIwnOp
OpYzc1D+A+dry3D39UGBNQ30/ywXXSDBWsiE9icT6lG5tHAA02AGXQ2k/+bNAx/JnlcODFUL3UvU
4gcC8PZmNK4rQAat8rQDFfLldadwqa7CmgIB3Q/JjVQZgetZkOsrlSS3JvFMSYl3UCEtBowA3YMm
2+0whr07Dy8FWoQcGVWlLi4Px3Hh4q0lavO3TG/EAOT7770J+lvQrU6MRfp4/oaxpM+omYxUeErb
G1nUSUu0g4eOwMmargk2m2JgAwiDb4reBBlAA9qT8mfnSninAMIwZYBcHMn5+C5loEQ8JUvu1DnU
fA4VyvEH41EJ4Fdsko2Rc12JFLOLhOGbbe/Zg/IyD8egdwkm3OHRFQGRYgqsxNDV7UIvhTyiepWa
B6Yd1cC4iiSJY3um8wZWf6JJYv078nsbCat2pgy6CJgTfkg91nHkdpC/D9vbAkKe7w6IQMdAAlk6
1WgdZ9fxuTjV1OiMKDxqMRLvXsGJUdzXf69E9Mby38JCM+7OgsksRNonOA1ks0cs4Vc3iBEVlG3o
nP9gIMXluuj4vAggKOdt648TwAf1lsEERyAReWdEjo5i5FkK121SxmQgvRhbiUtDafdNpjmmGzS0
3KEDc8drSr0pn/o23G8Wkp+JWPTSmbIE74ZuCmljFwpaoTim+D43SqvE6n612X9XM14rSH1UcnsV
gIRbv/ZcUkLEhdhy4b0/nH0z3+2WPnkfEe2XEHeb47jyZNiw/UgGCE77UM1ek5BjGy6cK9fbJk3G
DMopMHsMqRLClIUe61869Dq+lRDaKuQ/rz2Uxh5uoEZMZfHNNFUcFhfMVeKLlffbnEYcfc1esj7i
Pf/KYBxMZwkCf9TUz3aRRsLLPCdhFOtFlRwo5DnKocoPXXj7tO6Gq4t3Z/p9hRIBZKSPyoi2rZTY
bEH+P0X8ZzJVBV4vuuzaDqJolpNk2ZABpDqQJxHF+try8OToFcKZPGOYU0A1+aKv5y0Y6nFk4XCm
M7Sb2GfZSntv8EQduMY5ZWQ+5cGyWOHNOwmY2KHoOsl0yaOm6pdOvywI/I9lWWueLLgMfVz7KGqV
vdvmTEC4WelVP2PXocnMeRjV35ULnPWjcoSLYcVgAWFSrzKTYJAEbSXAMq9QvXNYg7faa7L471Sk
NBHWvIedHmBsALu8h4HWawJZsnP5OqVuKIA5e40QjQOyawXQaZ6F4RfucjtpCDSUWiKCx8BiiCer
4MPWrtt+hgUBy+Wz1AxlKxR37LLtlFs92a90ngbaBwBxLNavWpiZaksWtpUW0vRi6CWYrHTxOUWY
0vt/QkYfCsJYC+OT8jVnlK0M8GCvv/vP9Xd4DpXXxnps6fiCfp/3gsF60/8Fxj5jOs650eQPLvzH
BinIADhJ8h7Qx5Ob++yMlc/ROnCR9CZOrOrh5WtD8yyA06BrK2lCibJ06+m3AQSVHfXRdaD727+g
Iv3P+6XAbGW2Pma+Nks6eP0Q/jhMJwU9BUAcw6Uch/ZSHV7xkRLGAQ/iVMSAJcQ1Mw1LKRHhgux4
uqPQ3GMGRwQ/frUc4M2lDS4nH2HtUWJXwAbIO0/WajIbjssNUfiCuWJXZxckHaZ6KeHt3CFfgUMN
n7QWXdfy3hztaFplCF1qd8qOgXaST/Ro9Z90a05AYYIbwL5hZ0plwtGL5ZoH4rFMcui6yaKYgxFq
k5/xYCzeug0WoMdYJp+aHB7ocfVT7dXD5QGAwA9CV44F6rEpSeZLBTS0wPIWQaJVyK9HAe8eiPC8
mHpe6ZNLL/falwnANGcr3kX6WeUxOmfFsDy+HkGGuYnUoSOeCeXIccXP3bCxkDySe9hC69kxfyAx
L3UzGxJwMkMlXEB2FQtMKBpialjfeUoDBNAR/kOCGMp4Cnuaq3WFdSvyDSpmcuuIXavGhfX8H9LR
/pbzaQ7Ax9GGMu1KWL63rcY2LkKa3n52Q4U0lPpB9ILqmN01aVZGNuFufJtiuOhdfpvVUPUOsZ03
4Fmbps3uzzowE47GKNv7DG7T7f9E5QrIE44tqrlhOwJ07K2XJV4WZFcalVqFvDsDfSZTc5VQlRnL
6YBGBW0hpPx/qAHi/7q5GEr+kYMgTZzRUsdLZXYqtdK27GpjSI840vmSeJu9DoAs2ySZcH02BfIG
rYr7l1M4wSfPsOZTsYIqAnmmxeQaNcGO5wFbQD3NkfiwvQmQ0xaW6fJeG1AbrroPWT+qk/rAyeyq
HZvrTdGgVt/ddK0Rtopqfv4ZJ8EDr2JIo3i88bwyk4pFgK057hZ5Eg2lyHHeE9KzFduE2e3GuT5y
VlLfkbB9j7FsTkZKsuJu8+J6TromzShs6Dq0jJ9bQeN1cu3yg9lM4t4pwt20R9PDszQnXJgPrPdR
FG2O9muv9fUKvjStk47XHczQJRGFbevaH+jYO3YsXnPLWyhBKUi4Rz1fax9Sy15N16XDz1D1xlkT
BEjZPOeynabFMvv+Bev7gxIZvdk1DX24OindS2ShkTfbQceqHIw4dTACdw8/F8Tp5UGuZq3q6IC5
9tS5UAffZLowWdsKlzmNImXip5QXbWcGUqKTFCElyNAkwQj9tDZnR5e0fZd6QCPK5CmX3PNr2XQw
phjtr2ad94efx+7/aNIImgJvzXFCkpu2TsjXK/ILJbUbfQNRQbirQrFlspjBsLBRhvGW8Kp1pa7F
2pawBVrlPcvR+A2Muy0Dh+tBqy+bKT/6Hk56CvfN5PyPvFLRmRbberHJAKtaPBHgkBwnsDxy+GxJ
gdmGGB55BQk1ueyRwntdzNNHs/Al+FLBH5mHKtX6805SqN3N9aGUqPU3JhPihv954WP//efTVZa2
Ms4WyFt4v/jSAIUPodCG66w7pjTjDsRis98UXfelhP20VaTiYO4Fv3JEC+taVElrbc9eMkZJ0eal
z+kAuevLoTfFamn7WtXZHxuCcjyn751KCgYliDc/kHtB39VSNkuc4cgf402oEvNAJly318M8Quxr
buUt4azSxuI9k0as8euGq8Nl5GKKCc9SaFVs2INheKPPeig9rQKRK61F6JM1nua8vdmDjcUcaQSs
NYtBgaxcLdznoZhxUQWg3ybEUHuQ3mljo+Ouhxl3X4NaKOI6d7tuu7so00zYN92dUmLCQ8IoknYA
W338wqNFYX4Vb7eReF2+xB/7R612uX9CpxcocWn2FZ4OgACKLLCzsFvHmyyLTk2DBNXfqjp7S6tP
VnB14iFWdMXIAki4YFoEoFtdaKfmlIs+sOOZzypi1YcRcr0LSaGLO4AEz+v5cCkEIWG4hMRA6A9T
Yafqan3a3allolgkib451enCZoO9YrTfxanlsjriwnxLeT/W2CYlOiaoGn97ecRM2Q9doI0knloD
aGZeyX4A4awMBjjMmUe0e9go0w1yt1BOYslOLfyoBA2k129N2Ju5cyRzQBUSiJvFOqWVROgan2MC
qF6fqzPlDDjyTfTC1GLeKl0+2EmhgjoDCA2yAspKwRdJPKFuFnt5Byh0FBqOTGsA1u7tIK1/QuY4
zn9NK0VL3O4YjBxNEB+Zl1LTiHlZfA7n5YlgBXBXmXQQ33pJo1arBSjGR4IPe2tRSSEmSDqcdlOG
MaWMR0GNntXZsJKAt2KODDCcrTSLWU9msyr4GVFUvXVvWsCTmU6MdS23fnVh7yg39uv5/AmLDTNl
IOn9qJ1lSsY/Ofvg6Qw7eOgfRMGLWnlFvsZXjMPGVAw2Y7YtS3ZKHZYmjSXFkisGIYR/41KVn27n
WOTY9x7oS97P+U1WRsftd94z4pvg0QF0GGE737w53l3WjLSco5Zm3uYXNmvqiSegJzNl6T7Oiuzg
jbFJA30yNWsy+3t31vP5KB6meQXfePiwLZvQ4GQKZATfW53NeL7X0Z5wU2+3jczAyVVZn5ZSMbXs
m/SzQ+uJ43s4OJohkk6egZDDtC3Ko9CTQsyH5ppwuMK23vpVOgQZ8nylCsEHIjRDBdMxlIO9t334
++3R3qH+7bd99A6apsGzyf6EoexsLY8MokJjnTNmyYlGjwfscxl+n0hDMY1vt9eHzOUaxK/BFvJg
0u3/angWIoPeLlJBgdvqY+FB/zu1gW8QGsQKOWRl0ljmSAON+oPpS1BQnYrzfebbVTTH0cYVIQGn
znu+XBi+JwFq7H6u7WwP8qX8TgwUyqMXgMHzqcSUsc6v1dMaSQm1hIX3DGHPtnePqaJthaUihDpn
Epd8dhK9Axl4v8t4L9gwcxf7O5kFDUUsOkJd0eagDYELQSv0wz4Q9fDvvVFIYHJzLoZFAARK373V
c/UsBtk4UGl4X6Xv6N1M7HrOW5FhhQ1PitmZGriSQL4Xn6c4xyYlCUUnt0MjLKAjezHEPrIB9d0i
9HW60bZM9pV1FxWe/J3Idnwq2cWWmLYZfVEWR2QrZ3EjCrodXBKRJGEIEaX+q1JStXQhYVL/OAR+
9YJdVL378rrq5xtncuD3MK2NRW+5aGAkX8p/LIqQSD6SCW1F/YHspyW+wQA7JlGINdGtNIFFiT+G
yCxe7Ag/enSeqkSPQ1Smz2jXTE/Snc7gQqcJY5vjrK3uKZsudmaoKMRxUbWOKb0OtbgvmnfMb6Yu
UO+FAQJJS4lD/QmPF0b6sVTlJmYHdGAfBwux02QFFjaZrjUAwSuv/Q37pso0qNaALg0BgNEEssB7
WOm0wveIP+57417lKAjhimJIzus2Bei7MkanC0c7ZvPxJtEGj/wBKajZc1ALKtmwB+rCzVltY2BQ
tNR0U4uzhhyoJ3Cr/ezerBmZgw5+pGrcQcKTS35kzl/lDjg6iiDGwnbfKybnUta9WSoCROiKJXTP
c+taiT+cqJIPbqWenDJvajAqDwRu7hd47H43QeT/5KTXh3F9r55KzSpC1e2GU0E7ksK+u7I2Vh0Y
xSLqkuKoFbZODUJG4K6O3QUfFSt/9PuR10GwCMo2Uo5I/cCU3bC05jYnDsZ+c8SFkBGhyMFPdxKp
WG9UTF1WXzlwxrKinc8UvQbcLQOAqhzcmGLDB+SgUXM1GfbmuZ6BZhVXqHjTHFRB+rUTRlfLaqUp
QIMvMmbyxPrBtt00VE8fL3xYMuncb92FiKcSYbXDqw5RkpMiaGo3Q+E7+7qFbly5JElcSekSUkSQ
J0pDT6JYg3mduocZGgF6qlZ3XPFuQIJc+MxtGKzmvbmOXAHRJyKAdFVQX/tVyNmOL+RlqObCJ6+s
7FiGlP9bi04aZSh2RpGrOzj1M/uORFb5mUcVx5FI7H/zJg0gw0aKRHR4l+mi1w8TsZd8SONIMYZR
xOTEs5ZoTgTzTl2WULeOQ/t0Tw+EneSS9SLcJ/QEA5FSemX/pRh5awFN+ndCwCruOwx3VfQPgbje
lncnvX7hw9x1DM0DNJW+1XxeMwwG32QQ1NOqmXpQZkrbxukBQzNcQJtXdk6vfltboonqcW4cfykk
CiN9CKKcuDtNWRQ5J2/Wc1osUdhPAktmNaYG+gD0MBAOnmAons/DXneDaQ1KxPfMVm9XkCKti/fB
j2N0DCF9VgrRbB4ywCCROsW4HY19kiccPCZIiwxzHZ000JrWHwYKcwAGkgxi6n8Ip4pnOnk6J62M
fWWMBWVr/g/e4fIlHGOb5+4S8GuFo/NMbnuRaMHYNbOtiGD5tmhq5ahIgHCbShXd0HzL1JxWcgf4
e2ncVNhhIRvX/tvEx/sbhtt+MlhLy4Dl8Hz9GGs7znXNddXJE07mQ+HxDhHS6k2ZI1owbbSRHe5Z
N9dXUBxc86nSZZ2x1iBLYCya6/BJ8IK+v4cUEtG5OWEfbcmcwTAY2iz9cG84kPc3fEvIspmAcDl7
1FDpUflxXzmP1fLeb9cMq8GFI6eSJas+tMRx/86DRMgz4J+0zVdgolLeyD8VP5s+zIuYhJoNNSTJ
JxEOmEziln5dJ2OnBvQ1GUTHAfpA+jOcYgjTwfKqI8j+dEEZXA5uhdvlrlZP+fqf3r6JAuncAwNS
wUqBhZu3zh3nmLWJmMckOTbetDON04jhvrXO1eqSv87YaIRDhI7L+R6pzbSHYR5MmJB2WB5AnkjS
Ra2CvxWfCrUlgVKJxFZRcGdz/i9clGBrz3mMSKQZ/fWFcte1xOjGSXI9ebmmE6ovfZD4oeiDE/hV
3oD6zoxskftMnRUrv0IRy5QcozC7GMIaS2Ybozplwq9uJxuA+cEKtgUKBgJgTrDvdYgbHK1iMxgi
7B4BPBHUCaz9nvRznJZtVSZLd5vRs3G8e8guj6RYopoHjEHcImlv6qOGrfbMSX4wWFYuPRck4t9h
d7yqYOF318ukruqw2Z9UUPFDRWUJz4IiUOnkjOZwHDdGSe8z+sk2hF6GJ7dGOAx5oMGfgdQw3DoM
4DlC8jTscn6eZKg/DNnj6DeMZIfygqRk3b/A2GD/+DAcQCyias6SlJYIHcISVvbibRgNVqOfCR2d
myxsHvhkZ9janmbsGvwIMt4A/kB9pSVtVCzfZ9ZnCRUdmS6AYYnQdteezZQgc6mNVfuKZZmMO81i
KF4/2sIZmXi3rVABk4DWm4A7oVcLVZnF8hzAXyMTXgxuuzR53QDJ8MgCl84AyaxFyEV1YgcFbRNf
7xa19eZNxsXuxShS7WGFFPRT1fs5OEIorbWxpQNW/RZu/D2RZoqdGqQxoKyUwS7S0B9c8taKeGlS
iw4QdtB8ckfBQMqawyoL8GpapXWUCrJtUeXb4cblUoeUo5kmhgPue0DCcci2hKRm7rRP2TpxmHk0
Hlbcnlu+4fFYK6fTszZJxmTu26lpYanzR6IuPz4PGDv+18dqA6NJZ4jUyTdlNBopbWaebC6lSRF0
tDMAiIUDrwMNgR1HZTniExPEAopvgw8jZZHghtM/zTDii8X/fq1cQM9N6vHlm/kaG7WEq2X+WesG
gMbGBLS8eeHbq7FdbnKgfc6cZSzCrpWyqaO5yeGCJRfI4O2oDUKFXasRHRFkGcfWa0+PIBppu4A7
6EwTcyO1qxRomJzR0sZEuvqjWuam2wuXC6Zl8e3u7A8wxse+z3jCoY6Xqo3iNHNBmb0zg8Sz3yx5
W9vEwm4KRPH3Ays5DrCqxvGzEJ3LZzGDOTD46GvznEc2pZ9r64IukcSvs9ahRcL1kFwTK+fmNK3X
KVVZ7vsGakzQGVftW8WJxEfm1wxZPgMECj6lirWJrtIUdEtjAKBlAVNQiPbMqPYITUP/dxpXcjL6
wFy9Efsws2ba+wjNgFXWnn4mlGDU0l3NEM+4x90Lauc1oz2QXwssGx9oC56l/TAtR4ZMg9+U67y6
KmtRDEMgjVN5tevZ7MBMu+UZip7z9UpJG7L7+ZVS+N+d1f4oDu0dRHCtIIOgXaCbFm/9PgFOhnoE
gFAiw6MHkKKDOpMA6ijWE4Uhrju6nn/dMRjbKULyucjjklyBEXSQweZdUHDnrKvYCcUT71plgjcS
TKRVSNG0hGJwIxz4imb9sfrLzzI9cu9v5uEg+trv7syGK5IHxxGR9zA4O5v3L1SdXcQJmWezFID/
urj/Smu0KnUwtNw6ojXptBMpy+zS9Q0EWPbSmDD8Lm5O1kpVqgXfeYLrrri+YYHzDQ2cgaJS/zZX
KjPUEVjUn2euT14Sk2ldfaExrWUE+fFW+bMCpLy6A4OmDbCD2HezLgd6wzjFeqzyeqGa2mZHqyUL
rmHOzulU5kt2wLDluBhBINQD+rHI6kSnBa8B8nOvMUWlygs3WauMuhHcz574Wymuw8qlh8TaBCX5
z62r0nPXq6ACHRgvix/cErkERhhhp73GGKsRIveBnu8A8R+sLznY2jRunaQI4NhaqvfceicrPnwZ
HyDcFzkzxXrbe0p+/N4zCD9t7fRFU92xfX542p1HJt9Efx23VUJvj/ak3f3xZv00dbYBYoY4jnaB
7XCx+QqxpkgFgWo49dzIYn9FGx4sV4sp2Z5CDRTI3evWxMoc6lVhMStLpaGfEC4FIXo8owWgF9jj
GBXxEBpRQO8zbmXVNdBcCIRAv/Dl40BSMestIbs9x90JunvFee6QK9OhB3Lb7sJpnP0dY7moZ9Ww
FOPMZCNCrG+QTnkLfUvkWKu71klpS2F0uwVLaJXWVTtNzbCex7Jor90sgyYqfBjyZh8hcIkTzOA6
MHj6UBddvMUbELTG/rSwOR78TAkNIWAnpamuNIeA31Rz+c4GqbgfYnckDpl/tcfA/eyACorIfn1m
zoqZH93vn+IuoWF8aI0sQDPJCAfOFwQFeExzLWjOfJLmR8R4fnm2cxjALIhEJgBCwrd/YX3x3/Pe
45VZl7UKu//R8zYtV3G1HedEBSGBrEKfjlRdWNqfexqpj2pUQkFtTkHDpAe31NdasHlyJlUxyaTZ
HIi56U7Xyb731uYHGDf6dGDZMkCREUARTKhHta/KnTkZikdL/6L9k8td2ws7lYJitNRMozg07z8n
M/g34siJkKNjbkQ4PttwuVll5Y923Kuc+98OCr4Ti/v68f/PRlajRCEEaWpCMCap+MVWqRcM/p5X
8Onb1p49eBbTRvAHoP1rQlYr5agkG/AIt3Mqfje6LqAKJSIqLrWQBXN2X7k50UUOglFKxoxm3lGT
8H2H/XW32pQWS0qhYFjR50mJ5sKWnwN8PWm6JrhkRThKmpa0i+cdKhB0d/kllSVIl4XEyJvcDWBz
KXJZzYsrXULu1LC1pnY/GRYSaxXL6ew/GdzE1Byw13pwWwoH/fO4oucSllwQqfzsbHoYvK7on0QU
AhmbXVGWWUigjbHJx7suGfHhuJQrvPDGH2N7Ogkvpuvure8CrR3LxD5hFqs7xK1z30lHBIZ2IWNK
3UnzcIeXZjuK1pLThcmM8XqvCwHi0pKsH1rlOSmqYcPYNfjFbXCRm9Q3rFPZvzTgIQZDFv6KTXy4
Buy2Yg28Mr1Ie+GsY9sP2+jyhvC3EzMqhCd5PdxiEquwmtPif/2OcoedIjTHgcpya3XhpXVjlr6z
qJTUtshniGcghDzdN2JeNQgrZqcR/LFM9sHRh3UwDdXKq/scbeqq/1XPpO2YzQiAGdE8Ts8mGz+Q
CP88EQ1t3jICBIUDAenuyMFy4ooH/iYc8ljgV5peL1JGO2dSlfbuJ4Un96VTc3QEoeArBBwAmwKE
HtuQAu0lmtIYBaaJ0D8c8YJWTQyaRFN1RKhtKLG44Le9oUVuKdktukBvp1GAZAEsyeXtZCJgf29a
lV5m7HhoywywJ0fde7bmvrjlLAXNdvGIy02/FeKq5Tl4igckjvZrtEtxQuRJftmI/X57sScuxe5+
GIqNfv9AsIH7dt9iN+QzkvhX6XJvI4KI19bz1IHrxsnTjQdhwKLke9p+Dir9mbarm/UIVBpcZPPB
d6Qz9UKz1wxfWlTrazliiqd6zVwkjVrqUeIZuJVj5FL46v4S6eIi/36SIBKG/p5ckBs+2RX2mtZC
SzxLTSWMd1VslKGVoHy2prwu/LJzfV5IIbPRyMEcolfJROPdT1vt6l2YCZbYd+tnV53UQl4gexWg
DqaUr4e3fozJxeu8jZ4h+S8bY0PnZ9NKRxI0mr3D85xJzO2a1gfJ/ZxPdSryJTUHsJYVkXat8kNE
EmOexTMwOtLzPrnfnlkOfbovprC3iIAIySvgaQzlU170F45PXEg5/Pll/qpFEKljxcAU4IboAWvA
hZlwVf1krZExLSut6cPWHL0I9pugtRUvBB9bc4VkkK9PmOJWoAVTgP0b43U84VsH7A93XfldERCS
f4TItGRuL9mIjN8cJH4uqwuGV613Dhm1i8XrWZKR2yvI+pKBdddnYoBKnO6lRSFl1lArKCBYyXTi
rWBs1Esdpt5mxCqeOFXXUWZXVtmGPR6okgvTg8oX1Or8raJugOPw/0vLe6CMcBSFfCXau/bRpdQn
wU/wtvLxMCea29EktJxZDs1JV0nVZJci6wj6KoSa4zFUTDS3qiyuvaW47XjK5VTmWq2CEAYtJVIE
aLFFaCUuXDqe/FlofZ26rIz497ncCIq6TLK8Hbgx0OITo1hBVXo0HsP+oa4MRAxCiNJAqEV7pPR2
JhJMfgpzTJBwlA4fG/7rZQkPi5Mao09UdbAWIy3zifZ3HOqNCZI2LzOYCjVMgPXx/x9ms1plnTo9
2OTSOsN572pCSa9g1hIO0rx2M7LoTVv007gcyCl3cqd/jVd7w6JvLeduz4okkHF6dHHD+PoDsBDO
J03HvFuY1U/qA1PCxijIiqExCzA44CNyiRuUqX+B69aqfNIbk439Z6Emu5MAEO8U9zNCpC3wL8v1
LxUT1crbHvtwwPwDF9tWfMq9gAOlMqSpdow+LY4je3ntRa3GFrPbu3i3Gn0wOTMP7AC3lrybcMCh
cL4b0Z1VgBG05nyoS+z3YNmZQ+DVbWkcEV+bi/x1ZaVmBpkIMcqL3bkO212+5LEMO1giAGehGMl+
+J8b7nP7m7n484tizaeeqpQZKm1YX7xMFClz/DdV2RhoUm5MoF0HEArPjXF84PgLKslbmz/fWYoC
A4tzRmapjQHX6e+N3UCOGH51Symyh9cqWh1TVZWG7CtPNQbBxpuW454TNCFmavwwrBCoMxuX9Dpn
gtypQ0OFGK4qEQuZ5xvXwPV2kiGczeMGszJyNBUGA89bmgw6H/KWacX0lG2QOHzR00qylRfD6pWp
xgr+NwdFkI0VPMJnfe8zLr8Z0l4IUPs3DwBizxLt/vabokWEb7iUBEX2M3BOwizps1HjFxBpf1HI
fMGbD0NUkknYW7uIjtBknkyAbwtzTSINW9yJp6sf52T6I9DdonbjrQXYv9L14ItNmimhvGxlMPHk
m98CprIqrLxqQnv278xOWDc7BHdtWjMH3/Yp8nKG2z/hjyGO180bXsEL2giBZb3ZypVdkTVvL1mh
2q8tlwuutthQXXpQgqVEP5SmoSVLLVUcTgzVSAy7jkppA9BjI5gQTJNBu/oFAQ9pDW/Cm2mA/DBH
WuoaSTvXrQd4WCPyP1cMj0EnUABY73IkZUQafu1Cuo8OQ0SmVcwmWHnoi3aDQqN01ZvrQlFBuhSn
Hee8EdDhsYn6JR8tDrkOzP6WbBmARaukLdgmPTO5PrFtWVX4ldk00/5IMCaTR35dCaMHcGaQkrjA
MaExZ6PHDqU9vTNxh4998JgQ66fzjhbRqCWyt8HM9xmTfkfRattSbwAGV87XtI/vvHYpTvWhiOw2
P/oaxIKAu4iP4ramxDFBDFJREXnml1D3kMn1xjszNaRJvFMbw31XjFEmzI3cyf2VGPPSn1ShKosc
JsBUrZD6izuls+kkzJWpEkdN9aAeoUMS1ptX1+MsWwdqG+bFocV/+k5Bu3TnQek5g0hhbXOqOzGz
DY7eMUgApaLmp7q4vDV7YrRH6ilyLn/t5gEpESCNEeJdGQL5vl26nqn9IdSyIXSllqOD3RF36PVZ
xPRk92jD3Rfdro/vsmi16zMG8Um6gNsjznpn/8+gCv6+wZv3v9g7CpK3JUbzdlaBESjzhsrPAI8T
CdouNBf/QdVgKq2UG6pk+hj4RHSwqCfWK2llSLHXMAP55J3ZdgrgyNFpumd6EbRXU+E8K1SMqVwq
sns/kmjZ32i6bD7wTlyjO2BvdiHqRdpg29CGx5TEKLbVd7qXvr0E3WY+Qt4gEoKxpCz+ZtWR8D7x
fm1v/UseukvWy0ufKzgh6ssWrMPAwALpqvlm/nKZxtWwq0zwPkfOeBc1qaB6oramGHym0upUXhp4
f/AoDKL6nMLl7TckC36cdijLi9PRoS2CSvZMh0A5SCUZv/7rEko1TaT5gqEcsaeLTpYcwWyGFhMD
x9yjnLC/5PmRgXRkaOUdR5UdzeFs1mL7cm2fWpLVmHJaVNdYhkPiB6b7kWanvXXJ0VyyI32mTXN0
RRdBfx7gteTLW3dYLgTGWfp39EYdhi/q5OXn9yEzwuCZYcynvqDvIvERdZj5gkCade3BsaaES8iG
n1tqYRRF0Angwu6yg+WxxthfZmpw3/H+hL/MCqd1g+GWcneJbgiijJV1IThR/N33yox0snFxE57B
SfTh2ZCUohQ6NTQ/bviar2X2eLVTFxXGW70Cc07sSwhN4ZcdoBEg5N3MmlJ4nLQWdhUG5IlLlfzJ
j2/E7VNVk5QSBLk03LRVRl99XMDkyAb2lNQw2fov8laU0mRLObnKvo5wWQgoPlvfmEUS5Vjq53l1
yYeQVGJVioSa5MeoUBeB69hquUpE9BRMHVvpOzQkKPXY1DGj4svWOEMRW685bR6KDx6ft/Vil6lx
fg2CrmeNLfjTO+FYjI//CxTZx80wHsjKLHMP7SDM2h3TZFCo2M0PBLfSRh4Gg4IcSMJAmx/Sh40f
MpHdKExXKg/hBgRSbIt9m6K/I1GvNqTjWnOWuH9DVbkF7RF7tP6s3VX57wfwewbKWTlFygJpWcKT
P7G6HajpEbzVXwvWvx8G36GSB0VCt1PN6ABYkI1JQzHY/tc7+ZlYPusumihI8OrZCBMs6y8EziUr
mgVnz0J1caqpV478BWDgpYVVmbjwGy0EHEm56XB10wB1byKvx+w/vrR9TK6ilAbq2Ss9CtpE8SZm
3+FqMI5+75de3P7TrIrgqxI4W9102wn2GMMnBqhjkqvjx+IF8dBVDPf35Y9jhhfYj2xsPQWXLXRP
JdYgJyqDZvvzDO41LjsB3diq3e5zXyrT0jucq5Vnhjtr/RPocnlRl9xKFpRabbkAlvsY9FsjIowW
Ubs0z9QYk6xd3a6rDKVsZkQuoB3f4UB4NgBkvAYggB3fk6CLoBfJQWhnwmgMlnXpLt121ERC3sWN
3T3sL5fm5pXfwjmnCliijSzdj/dUmuDhBf8BtuILZnK+Q4MNhWSXn3QzLDLGg5bJUAk1yZX8Gxt8
Q7IZQx34RCPu+RrdvoszYSoyhJG8Wm5cMui4K6Ibbesc6d4//emC8w2RWL+T2zxLSNOCHDPMJtXO
IvSnFi/64NSQGw09UjzlZf7vBfERn8xvinmzXnrRbZwW0KqI1GfLGRBASnQ50pw1jTvZkb1/mdNY
GhGFQyWo9sWjvng10ZT4M7RCQbQywpG3wOlRii5OCsHlsg3JAv/rhoqDpD67UqZJWoFXN1prF81v
OZVklAxVozJy3WvijUCntlbAWE0kY3Bw4Q5QFnsYjraHIegn9P2qRrCnT+fzUCTdWMcp8RL6YKjG
wMIbBdreyaNzckUw9Qf2IcjyrkvyJWSKBmsm8tODl1BOmbheyA6SaQiqUwekjd41LBd1dHSn+pOh
RROiXex8bOtWOlp8ok8EhCSSOgbbr23KYHZ+0UlSLaI/dKMcOxIlr3zzs6dg6tCf6fTEKolCB0G2
ouH2z4ahZuFt0UZVVMhcDNGadrD3Yi0q2XmgFpyo0OfAVzZgNRZeAAzHs4HdH0A8EItXBmf0dBXs
BL/gPGQdH8eZINYPtWmcRz+kbmC61j4XUlqVj++nrXVReeuWYBF9FYdgU6s7LF9xGuZcOmyVqNjz
a7Y77fJME3EXIGmIMlabQRy0j6uuI8Rj4ua/lMBqVssEnyhwqrYZTmb56WIOhiU7B8m5SxZ4RYRL
1Y/3t+p8oPyPj8o0GFQxJMDp1gpxD4vl5XHJbu5DrO886Zwbud5m3eY1/nCA2z8HDSuUOe8X+vrT
GrYpshMmy+e3R95ouPaMaFXdK61DmM2g8GhSoON9CO+/MR2/W5AR396xdrtEKupgisMfY7d388CI
n1dAaR++jgWDBrYfmxkLpEyGpg7Vk/iOnYDxOyS8VwxTeg+KWVDCRAPR3It2G0y/Ld7tN5ZCtnCO
7ZH5mJS31xv9nwpYu2Um6VmpPhNlGdALGkgfe482yNgqutJa5TXBeZkIT8WgWBBxHw5XqINtdjOJ
9B6e62ZyC7Fg6XxXrY23z3ziWaQ4iChPckASjo/bMeihfPf43j7UPsakMyRioBQORXH5m96zLqi5
XT3JdJ/rLa6wvRg+jfIhjhwwSJQTWXF4HT43TFIb9gBR7dBDruEloLeiVFzCzEtYhPNEdLmRyEb8
xaqls+zIqlfBEHR7lowm5jsKtRiuJ2+ZwtbRlRRxO8/GACuBM0Q7dcL3SfF7wvFgSrIqMpX9X9ij
rJpeLjZ7q1nMIm6/S6eT0gmbtJ2w2GLsTRKLw2CUm3YuxZIPuCC5vZMVdUh30VOjrlQKq8H0r++h
fA7/2HHshFMc3WIy1fm+I+r9eN62KFJf7KW4Nisu9+GxWklbbjHTAERjcmAlQeQr3+AzEIdy3Pye
rtLj79OI+2ARIBQZahUm7K+I151m9Fe59p/Dq+81nV61LAxkm8eFBp8GAcIG1oCCvxsnSFf1pRpv
sPQDB2Dl0orM2zohQPvD6zX5vA3DQVClarPSUYAL7ZKAa4DY/RbUahlsrOI2vDN/tZmxnoO2bDeq
ktoVvC/PUHOAVsHOipNDpWBdiCoLcDlSz4NmGRXCoG/mJE4bQwKT20fJORwQ3R41Q3peup5pzVXx
VHU9pH4RjhuNsCyz61otTXLKsk011liX4Eu7sZpPvmL7K5kjCE9XdaNKpfrU5aYZ0uf2xJmMq+YV
49f9GDg+FHMFen8ZA2yq7bzgC5gx/yumELAktfzKQ00z4OZIa2U6JxqmE+VN6nKiAnB0LSE7/61D
wfgLpKxOITAmsZXrpVRQwW0GxvcI9c2MGwWvrsuprUrPI06ua+1bn/hv2v9CSEE8jseYJ1bgeXKs
jjEi1Py1Y5/9s3TtHMt4Ko0k4a37GiZVVhSKGd/X6qcELkbk/np9iU0SjBFsKAlNVFiETBQXjCKL
G5Hpn24B8ZeJ5NjZpJi94wv7J1rkXpQfjbro5iMY8iFxsQKtI8bSkGaf8zthwvhkud42WYDKhQf1
4+7WwvU9lUbAYizxl/de7i8W3RF1H+qkG0XSTru6T0+ZsTBeYVHbFQw9/nnGOwz9UHWnnBx53oox
DMlneH7kpz949xeOjdRTjviixGHM7mvvxof4PhLzEEpWjRj33vtyzhuczXjxTUXtRirIftrU5eFw
t7Q1N3WhzLiTEThyYTvPUWhKiKP0IeWqD4AKJ3fVgY+6BjaANkHjBnnmi1r3DxNudZjnMndEH3g5
nL5e/6rRsERzs6cwjOAuik0scDVoiQe5KRshz9jjIR6hfQ6alx2x1jVh9gZwckoTixr/4m03g0PS
FEd4sI5aMhNlsbtuOz01/b6EjaJ7M73gmRzzQJMROVvOM+LPnuXxf0ubODmXSNOTxjxgGr/pGXRO
WLWcjS3eVFjDCLmVdpdMuioByc9iWGcZhs8B6mWKOSLMSFCQMhhHyCezlbA2+6HTcjWNGO+pkaOK
GRSgUFNEVR2tWBMTkMI/QIfk1mZ0kqH+7SvqMUedLUrn8KcnLvwd1gynJpXNKHS2hmZQ1ITFRbB9
cfkCnB7Vnot8ZKmrq5hspDSCOCYHvRqCznc4+0zdUpdNOyO4gKLSEulMNUoKVYpsz5SJWVK/YMey
dt1Y2H/jx5EMFjld3GNMxOSqzg50MwVr1BiD176OZeCjIUw1VIfuNgD45jNSXB3rB7oZ2RHMwXtR
GuZm0ypcF6Bz1fdIFFiYY3dRBd0qnC2uAKix7aMT9lgQIk8V+p/9m6igtYUktYVsHYctBqTyynwl
3fT0O+0sxIFOnRu+rDGfU4S+J4ggrISfDyhte3f/s+TGpof6UNjsMt+aaz+Mkge+3gb+6lN8TBO3
Cjo9/0aRdJ0PXbUugSTCGuFW4umdDnZLpyRDaXOnZv1wDVLaio1AqmOpFozvsi9RFse4A5IOa7Xc
dEoTCvcM9T4HdtUmmi4uqjfIcZ6qvt9diHCCl1R9UE43Tm/p9+v0P2Q2eFHOscgZxWG/PyTaQa16
W9D9yhUUxLQKjm+pHrzKrUaQn/5JgbOd2Z+iBGzqeNZCjE/TLQW52pvbQoBf/JOLY9QpzNMvyFWw
LTfATAajsMoqJyF66cVXn59QXnbNLic11OAljdr469p9FSXQb5jnK6psjjhU2koj31YeXBN2DqrS
1WStw8e8AgiMo65r9EpB44RMnIyzC88eMYOT8UE1VYEYhjWD0Hqa7NGiXs0LD0jH8WnEHKjiXnTM
zJBqLzONy06hyF1JkrKiMxyXhpvOwOKu5QSQoE/htDAPS1ThxGaiV5VqPkMKDzj5DECnzGE85ZvU
dTVMtbBXT8ZnOZvQ1Om8c3xorFrXFvbzNPfyTSaS9w7eVoS9shFMLBeszZeJgBLx5xe9AOMiMMXB
12sRpb82kXC5kkmz1q8trSF/GvWPvg6JjbAQlupErSrkJubMxI8YV/zLi1kDgor7OCRqLDfGFeDB
bYQypH+g1r4tMeE5yxBuZIIGCHGwV+aKPFgrcK9+LOs6G0iF2qPBtfKM3FpR31IhYhlWEEpmMqHx
JsrKGPmuO6/b6UjFE0aNT5fLHZGOAzvrAGU2sFjMddp0qrNB8ZEGK94LB0f+hCfyKhdRMo9USBLL
cfCLvlJMAdKIVyszZF4T1eS9YlZ/dC02rjL3qTWrS9bFjVgdvUyGZbfpFU3JIMGRnpR1XO3LkVlH
+U6FSs2Vhk+19KU/WzwB6iHORbQtGocK5bxMlGokP4Ceezn2aIIhAtOPID0M7CqgSBg2ro94yPWK
3fKmSOv9r8uhh3bgNJ3t2mtzU7q/aZ6IyQKDtZBDOLSedkSByELSwb0IOJn7aBwY2L402cCMUNJt
ILFhhfMufUuWBFMuatVZQenc7XP6DmnGjzXtqdvRIHN8s7KnQvK1biUkYNtsvflQw1NzOXAjI6sw
BHJtLDZc/qbcDO0BWrhoSsSIO+89SP03q1HZ51/uwnC+rnhc0r84Yp5+nNCYKKNYctr2GWKtWgxC
77GV08+RpvNZZyKc+I14xA8Yd/gAhwLAUqvY7XbXSvVB8jfKDw9jOYq+nxAOkqb6Myjax4Z99GTB
BYyac3oL4hSL5wQW3V9JqOpQ0A/ig4llKtEvyOcrAbEFXJQ+wxc1D+iRiGirmaRHoRycqTEXFIm1
QvYvUgtu62nOHe/6Z36F65INrChOQOMocxGsGMwouVdNUjTJ0h66DZeutrkvxQrHqDDzvegdUTkN
faHe5vRmHoaNyyGX8OY9G7Z5oYZg9WePNhM1mXRRmEO+5FHJ5VtFPGp/t9DAxEKxJW1wYFANLj8U
WLixIUBMDFmzocBWtK3EtQDU6AODUwgI4s9SUdqJOVRIYYhnUrcVK7dnklZPuQbdkYyu9fGaP2Rr
PtVL0voHcOiBuW3vbmoPrgL6zA+MdHDBDwA8RNtLKlGzujkXHooGhFV3fH7JnMmCZG4yvjQEDxEV
VBKYDqSkXHHCoC4n8viaXYWe0KdDttnIrdgIwh6rgjjc+XsyVvwh4EhMM7zj+J0auAhT2Y68MhUb
ClENmaX3ANKBwI2sGng+eyNobLFxaTx1+7a6+XS7GKZg4HHVd5yB8JQ5vnJNk0W0vI1hVtYLiv9c
MTSxdPPTX4oMZHhdc+acgulIIKfyi5mc4SIvlb7wz7Mhj0ex1nO7oWhvm6T8kFXQB6HbMV06+PQg
Kn0pjRoeSJ+jbtlrP3uitTjNPU1F0ioiUTHS+2jZ/9xtYVE+rluNO/dzzcsp6D5nXXwYOd5n7Arn
RG6dwUb6tnlDyPKJ9TZpYZyOk4eMNrkpiZ/gP05pgP2tzKGs51skF+BpbWbuCvuv3ub7n0izJELg
AqSEi1hnkM8Hj+u59JHXu9sVNbGgGGMbsjnrT0RYZlmThwDSfXYn9Xp4/sMJ5+fIwxHTyhS16weZ
ywvOIRBMOj56+Fy0CofwfymCsSVUMMzMr5M5n1LayB/PjRB1QX0me7zT0aaoxf6V5fsHA1e5F3jM
xIW/FaQoTlmptMjGL86Beixm2ZxmHBYuOHyZGmhdJY4Lssqw7f2TlmRDnyaP2rSstfMUompIwDRv
RfP5KOhNBWHOapOEIbNSJPbbgd87mnzSyYZr4B7O/y4EB7SWsp99TNVkrAY8ob88sA4iGMq+AxID
9SkmJZI2/LIFg6JWGmRJz0fOPaFBMXLD1Y8jEUPyZvsXqXZEcPyOUbyTfGU4Nc/BB/mPvMzYWnRB
li1vuynPCVK53oOWVjVDbWE1ugC/hM9Z+jAeY6RuYipC8408HoaKBAhjQvjYYXSZuITSMiVPYzdX
P9QDFjZkY+D5QNGB+ZiX4N2571u3ZNyXboCxvUrA8CacemjgHJHqxpiyjoI2P2vphO8m4avbtA3D
a/u3wcPnQym3ynQ/tGc4HsAF960fgPH2a12HkZ47qnNtEbrS7KzEV1fqUEuCQL3ag6qE9PbVr+rT
wReK8VCijiNBTJezxcnJdnZhBUHIPK0bM0b9HWSbq1u9dnNL1+pz0FgIxpQVAp9whaDcwqRfAFnv
Sbr0poHQbyGZa5FyO+FuymEC15MFSwtRqM/Qg3ozRAtk2uPIWmG6Fblq871E/yWrksqXbtN6rFRi
hpoKVbTKEpOJbfsFd8NafhHZn+Twjjk8NhLjbiRyHT/5UDHnUJAGXUgkyXC4gwYshJjPh/F+32HX
1jYxqdHUUKhWSzmUV8g5MEIx8y+p9wrS975am3TNDshmXiwFoXcftdd/Bv4zeRcvf6nXXU1bFT6n
NY3PII3tMkOmaL9kXZnTtF912RmVKduPsFp9R7auabsc8Dekb86SEyq196zsTfL+/Ew34gUYwqph
cYnKR3k7mZjKg8rjlzNkayhNv/CB97BvAyQmPkeGkWj8KGCayc+9mBiLrhEOeAJ9vIJWqryvQSQy
ssEX1qXv8ylBUJZtJfER+X6yPKCvfLmosSFqSKqJF1nXALjzlUXuy9O+z/AQDj1SPa/XuKa1x4Ge
sjLz6b7eQwngc5Dd7KdArtG/GxPScLjqrqG2KVBnr7OtX+g7MSq1459h2T6+mHlkkCEWmh8irGrQ
K8OeM9Gz9s9EpdhUm87ORU2CUFNJfKTppK4Rh9j8hOsU3NY+A2foSoYKPUBcU//h49GhQ0gFogXN
l9eCIVLKuCFXtmP2BQ3cIsfmf7g1s7rCvT6oZZUzqqjJAfG3vTOP0MKmmbgHe4y/bcdgUiTQjt47
tiSQLNWlBsYiIW+6x0wYjeorG8fooRJN6ft9qyTj2IZoKxnJ5WaJNdKtxqh02dQfTGNcKrcVVxXi
Azmd+N1MwTVaQxq32Ay0mwopKZ2+ZHHZFz3zhXnDYxu27W/nS9iGYolClyzGFVqtL4KKrlDbkhOd
W50VXCTXfRx2exz+1SCYXsoy/HODS8q/KI1umB9qhgjdJCAbkB+Z8o8FJUwawwT9iA1CuIYlM7ox
D/Y8FaEWmLCgC4Zp2HDglAOb9MT1Mmn+fpxgs4EuBqMBgbqbGgNwqhYc+TVZvkxEqeGLaD74Cfot
VALUDyxJfKG9VV6H1qzsMwIxOZxxHxY7sqfKPJUd2VsVELok5FdLldtl/ZwrjOnBeGJuTazn18bH
PhDqNCOGMZ9nSZUerJCtJDwNfnXBVoADzsD3JZ8mSW23GhLMKSO+kpbB52F0bX/HXDIcyh3K5uVs
X5wmdiAL3YL2m2PgZAoq805KXlvn1mAfg5zpqWzAC5shoRmup9EUVj7cKe1355HsdmgruyzAqSlr
R1Oi4GFl3fRcVHSiRvEEIROG1xVV4QEUYL5XZ5GMiq+8zKrdraokYSk8TZk0jZ8QLiVegUUF7W2R
msX/s7zYkmzrb/DtWbjVekYRQTp0WuuX8Sr650yEvShbkPXPmXeMtBpYHAcZ3OpD4VKNPu11KHbj
n+Kf0cYpL4pXxTmJ4/zlsRQ40fGTTkEHr8CTppDUNsYA4Pdc/PyfSvnBEY4UPIRdccBGtoYa7P5B
LMlDf8FUzKXJIQ4O2yECXqXRZN3MxVO0SgP9lVCT2ftykow7OFskPJV9SeP6MeWmP28kvqw9OA7u
APDGFbKeyPU/DjFOFCY/JnAQmssCP+nNnqE0hm4KWzzH5GN5fQcMzr3FdEmGVDNe3ETtsgmqB1xb
f6qm48QBCWv3bGhtOxBZkTV8MFpPkxz92bbFAqcdf+xtGEG9LXsd/PsXWBP3skeIolkNEalczTF0
Xd1CF61uiFaXiUvWMbIt4weFROQ0IrtJACGdo3u3s1AryQJC6qQE/J225NnsitDLBgmJufFi00Bh
fZ3bXkv4SdOB21eC2laCYAdebf6R7fAf40vdjiE0IGma72+w3uzcPuj6OtJu860uHYobKek5gICG
bwp3j9aTy/3ZAbl2jHZzXtCxxh4p2Rhk04J6SF+yEC9nJF88+3mwSA5LXMvHCL/Y3nOpkquQGC/E
R+36AZv5peK8NCYT5xCbAMpyX3U/jCpKZ4ycO8bB7Yi/WeyeT46cFBFq0KqfkIWtazTe78yMHGts
VlcRkrLL2Tx+hlKWsaKR96MY4zYxtU9s18n3UXlBuXg1/ruapgs+aMTCkj/jXoeqyAnC9LEqH35F
z+7xVzy5WRbQEem4t9keWxyPheekbof6WbO8uZpmz8No8wjrl7RFnLpa6pwB11CJ3xZjzn2RqgJ0
M45woUBqg1/ZO4CYG/nR7LBjHZkO96FilNzoujS1EP55gH9s0F1x+cOCi8nIJRtmGouks+LHn8Aq
oND/7b+Kz5EqEbD2XcfeZ0qWGpyGYW087jia03go0xjpAMBag9jlYeY1SwAznRRE26SXKEmqy9zS
pQbal9tau6zv4Z92LbrdkE9QiI5coEv/1tM0orZ+GRiUdJ5nUYXGw8twWzSp7H8Tc6CK8+5MaYxa
jLOuPENHr1zOt0eM/rnntgQDgiZkGmA75LNqLe9bIBDZA65FbbqmRL9r6SX8VcKxHJikqnyA2D4U
RQq6ilWSstuHnimi4/qa6JEVtBVHtCpTpDblj7DzD5JnPXrpbhL1yYe/q85LEI46Yy4o/sFSn6bH
VumWPu+lzC01z/5I5RvJW9AgTHnivRKmm6GPHNDn6xyTVbPck/N/uxboEL2XFIybzzdJMyD2k+dX
w60PVUtibPh32WnYkLsJZ96tjZu2cd3qCZQXdPoGHKPgfb1PefAIr7uWrJ8l+AtBMvdroHAm6f5I
vsnN5+RUqkh128EiNR7Iyv08wcFdnW0pP5jRB6woVSzOmHUZq1sc10AkXYMDRRw/1Ux/GpfDzDdJ
kGy4VAgDGliu58Z2p07SxV83jlm7WRp+wpK7ZHPfxf8go0U0/CT3f/SCj3R4wPNtZkOQS7Ss8UHh
CfTrC2UlWXxeVI1BB8GAMWsmrRD0vvykru7tUhoqcLNhD7LXil61cHKUA4BbVAV8g3kcSmG1HnXZ
HS8vUflwwiCGXOXY0+ySj6fb7i7z5Z0Sr2Gl0Pg7xdNsM+20meWNL2IT8K5Yi2p8m8K38JcAvYAX
msMA1zRXOubAyxBTCfDX1jlFyrPEzh9RF2ky6DdRtyi/qucMszzR3oCkj+IUIf0yYWd8/T1dE1OK
nLWtyOxTAa5NrYk2vya6nAdNx+hFmnrbVr2q9VJmcvxwNMWQY62IR6LKWD2gJtD7MFUFwT/1Um+F
jMMTa/COQpVIvNJSWWGNHZZchFgHsq40FkG6MmWJSv9b2yc6cTnwIPCF0B+gtKlCSoUOYCaYJfrU
/sH6n5vao6HPtwgGCOBb2vR00j7Are4K6GONRqVhMPxDptHoTQPhZUJhu7Gq8JWPOnRTwYbvya3s
iVy8PfKvuqykrx5fGJYasrdDKuEtK0QEB1snXQ3VY648QctvpesZkRQqrZFWPEhHQ6GhEGPekEMe
YrUvn5XYoNPmQVCtqXh9CGz5WtoRkbvyB6OFOb62/mauIgRpDO8wXyHd8/sSyctB9GSZ6mo0EwTJ
6dhygh3326wSDWX4WsYqAuoXi3cx336UnfhUan6VzLQpuczNdzGa7q2EWCY7SaA6XAyXPdtBunEE
BPlw9NVCtEC//zqoGyK/CIo0zkfqP4EVKYa15UcDbDMmzmszcipzd1xfFoyBB4eci9m47DDRRHky
P18EvfsuPIgcIrJJCpuUWM2JDyHp3JDwiL7Uq2l1k3BUswsdWSFiU/jApBXCoZO3kvWIxfbUv3iQ
I2QGt2A2Vk9RB0Qj1aVRk4JhZk9F3p8qdc82AaayotB3xk+2BbBlb9aaUe5tlfNHpU6AVQCXiiAf
JrS8c+MZWdp/Jzyzo5TaQUVt5yMiSxJIap+KLvFQ76v7FCOvk4KbgppfS2rovxdcXlZ3hRAWoe1i
icHjQ8MX/7R9vRv4+aVhlgvhLrLiCl6m2qEI0VEwSVFzivKepTFOkoeugGFIc+TI4HEmTW3C19W5
axlhXI+nDuy4vf6ldZsahei/OLBlCpwBKuZivVEiQh9bMQ1HlIttv52bvqBMpWHN8S4+MY5CKKiz
B+PK9yLXg06h9odisSVDQN0nc6OjwpHyxdWvscjcziXtz/a2AF4CtpimrtCRy7tHUnxoBG/fWfat
qXJ02DBkyqxw/EkDEFaFxx3UNZIPaekELnGQul0E4AMPLoZ2xZetwETdgsfIWFoTRVxMSWUSOvWU
1D0iJ3DPQJN0ioIfLprLTHNmk2k3wY98rbWJBjOAGrXYH2th2jTb84BxtA51lyYKmlWWSnvZLAFH
BMdSZQ7fOwlhdbHKPMpEjxIVEIoI6oVR0JIEEvksnjoVuxZT0Zp0tRC9bQgmfGBM2wt7Lj9CYHh3
+u1ZkS+EYna3+RtXUwmZmTSRjDd5wuYvdExlqPpakny0oNT8qm2BclSC/6OrNiE9ko0VRdUUSaez
RaxSo0JH5AjLWLfwUyoSadvt0DfeA1FSRw/1bLFIhny7CdVErLNmjazZLrvXMM2vpb7B66pVcbuY
rVdZh7bnUcqyX0Bm+6vpWYyIQy2cR94cDZUi/ZScK8tpcagNPR2hNTfh65DY81shUeGzFT/gTAMH
ritXQLzmHyBwD/WZzxs3GVRDCexN07HoBHcKPikfaZZ/YayAGFa6/7moV0hrTEPW8+Z2fjQW/87q
c677n1X1EC9wuLIUjXfD/owH2pwe2o5o6oI1+1giI4s4DBREYOVZzPSNiBNP/oPZmHJ3hsBUG6iO
Tk1565riy8jEIdekfe6AOPvpXgfh+ecgBHBtWOwqvyjbbc8xe8JZsQOFmUx9U0U0Dla0MthG441S
hb2QJ/Pzy2dqk9sN+wbcd/BFEArXwwceB6JlPazwO8V4SdZM26TQ8tlFuXbnjhiJCXgDDgV/KdzL
o582c/z6uDMoZcZMLLKjk8nHgWmpd5mbLD4yxQzgmXonZ7BAhKJogXh8dH33Fmx1OC3ewQ0EcN5M
ubz/s4EyBB0gOXf1UyH19sqol2y7VYE/AyrahSH1d4FfCu4CXSHDrnZQgH680XLhSehDFbfAT/jX
zNPaDq91b08hhoIHngBO4v1liQwjz/JPsiJkPPy4vEGAnopz3Fx+mY4bCEFB/ih7TIsJYR8sXSnw
TvXHZZ0qTZyhJTryN3NcyWA43pAxNHi3a/7cnEMSGXccxf2fQ1LosnJeBYx5s1A/BDs2VOB13uzL
I+xbT1Ak4enFVW/i0/Dr9lE057oaClwhpsOC+S9UUMcvitiTqysJNelwhQpq5bDbgJR5Iuc5px6L
soMwrXfh8ZvYJW07oFTfkRtrs4jMarKdWjE+Qph1q5tVsUyiGFOelyr/mljgfjDCkR4x7CNxkGmW
wJQCqWMtT1ZsNYeFINqz+wbjSETOeEPhPSNCgY1Kk8RNQgxBhWQix11tZAXbCL2VdVVh8Ullewf8
Y647Wk1y/50o7v8d6c40ZeZ2PeBkqGfm4d8tWdCKwBGAtxkjY1tinLvLXGS6CNNXhZbW+sGbFzbQ
q6OdRvVsa5A3UGB5L57O5MPK0NbKYEpZ3sFXECRS5xe2E9TuY0rlKnVzRmLx2JRRFqCFA0O15sy1
SBixmzG+TF3dReaMbKtsi5qVw5k/L5m4h32mapGmQqWgUJneZ6FQHEkcQfksHjvo4GF9cr8ZHPkL
YqosmFIMaUocBCn1b7WsVizw+PPe1nSh/H9V2UTseJHMDY3eYT4T4EMIiCZ2INtZnQp8Tkiejb9X
CInVCo+YtolkIIkF43mG3FtdaUAmdVShkmNlyHo5iq8lXX8qS7n7J8hgsNUHFyClj4o7Hit4mQHC
TNYzKDWmPKz2XaWl0QvX3I9N33wW7xZlVWKTUkmtO+dsNphg+SFcbfzo80nL0ETKD/+CksX9vyz3
G4M713P2url1xn/yYkejMWcHeuG0MLNmISB3sgA5I5wFgXRK9TI1uphng5buWUyPqbUyFPBEXkm5
i4lf5NI3Mvid8UvBHymLRg8j5pAmtxrwVwpT7DSm8aX9PhtRRwOzoJDxW+T9jhRzK1RA2cHtCu1c
TWhZM7ZdIRNvICnNK8ZElPmApP9KwXfqkH3UPBlq/wcjLqTFJGAheFJgOH/788B2K4vQ4zbMvYo5
8VPfa2K9dM5vnfbZNUqDLGCgUt71KCQj4hD+VXfeqiCkHuLDRXcWO1s9G+pvVPyfmfLzCBg9fldq
i3NRYbOWUrSF8GuwdJiDF9Z1Joj8P5oex4NiU0OSxC/Cgj79WKP5MUFu+tthlG+M4Rr9rq9ojOeK
XZ9dnPUiE5UhUHMKJsxu3LEVJ0nCZceX1Ed8DjFV96ad4JDeGLNvnov1lspNTufbXDjM78oUQUh8
Xs+ZuOaWCFEo4A8WCVGenOfQqvL187fETBC/zIBYm8/wzznFhFi3QBr7eOqgaQMD1YkXNPJGNLJm
jE8+M1RZnF8OCFFvHf3lIKjiftMFdu8eXsQfeKP2OEKzhKRhMi4iU04D2arDmX6tS0bimwXaQCHk
h4PkKEtGxxKp3Zo6q5UHGaRzH3neKovsXe1hn6YaPAo/uDklDAkw2uHRUMY2SKAPzGbv2JfzuJ3v
96wtSvio5PTelxdkdZ4uMiO2uAbuJO7GJkiLZhgNCa1n+ZGyoT8t/xgjMnZbRux38Dg0teHtHRBo
JkD4PNmPu4el55uJV3MBgfKZ/+uT6YOQuUf3G9ljlFdt1vgfqHqju+9/Iadwg4uplGxfgid96XXA
nVr4DD8X1bqZbQohu9OcT3nQ3tTN03m+BWoBeQ+UKpe3G939lhR0mg1rXuy88H5Q+ts6GomKWcku
r7bVU13GK65gHPIQD2xtPB8X1MDs9ZeYY2CFe2SW9YHfoAi3hvSnfwwiiphLXbYZ/dvHf16XcyZ9
SI1NyXjc5z8rtrwAAU7UwQF0Ru9+6b2or7Nnh7+4lgq/o5xwGTdv15vlHm1MBST8iML02v12C+kZ
hftceRIC1L/6XXM3mY+dtZjv4uufyBeeMurFe4oLzn3N47xvT9+88vH039ZLsU5BYxQrhCFjVSaK
aO9v9kxr7vH8Xe6xwGB1zct8z+8QEvdLCpSzu6b19tKpchqZ3IVoGhKNSdsA2Q0F42Wkv2h3ReTZ
V2T5oIOGf1bWr5p+hHBwMV8CEqFoPwR+pnsH/m+RKjAj7eCRZH07S07OyMuM5pxVZ0zeLsMnYR6k
AL26vLMIq5LaE8kQPUX8oGBjW/4twbUKGmbeTzL/Jj67c3IRqdvkUq6k4/XFdHtOYfwcYyoluzr7
OR/tgg1Xqf8OVakvEB7CD4DNM7xFuvl+k2J27HfPGPDs1ujVj8wbuo8bCaH/b/3/SOcz9+Vcri98
V731iCqPwVBw/bSxd+BLdBcsJ6TuK++gSxWO3Bvf4VvFWcoRfWskUBHFrnJDfzZzwiaywSyMgBwi
ibYUNFIsn3MCBQXzi/l+e+6A5myO2OScLxchPUQ3fFEp4pBZZAwQMNmvmSdQUXBLmFS4T3sJ682o
hi6jUkKHKB1+Xy6BIqz46wxP34kU/4CcVJvJcq7Jb+1Ex39agSaxoCuX8GAHwu8cEIfyQ60XvFfE
MRpwPaY5ZvGnbeBwPfFgh8hwH4W5rpxZBB0uLabBAtZuD2JMXTxLbQuiRIaqUaOC+mkZqb/GOEYj
1ToNmTtx7RDfbU1vQNVjn7zVMbYQQ3oE+bRYGc7mO0uum6Vrc1Fnh0Q4u0nT8B8NkWicAR12DYf9
NZXHw5Jz4NhKSX54pyrwIm3Y4gL3hBkEBVfQrB0rbkF4gRNcteUX3A+ViHlVsqo9Duy8yWMbWQnE
vKg1CQj5RB+rWQzozCmh3I0DAZPyLbJC607ULmpiUzWLKRFE8jw7ZlIuHaqPVJzqsrPAhw3L1drs
mfMoYyLJ45/QmOI4bHNMMvRxLIdi4GbdqE0CbgXb5KO+14jFkfJc/hyEBT+K4b3LHgCG96DYl2Ia
7l2k3XxrMACGrtliTEYHgupacGmtVYDmithGScjHzxiYjp9OAur7hJLKwXLSOO5X8Rx28iLEM9zS
iPt4Ku54O/z30qEQU14qypPOTwFQBlMNxtjJCRGV5pkqI5yEGyFlQr9QFVtC+HfMeSlNzJdjKHQQ
a4jr8T+NM2Us8iIPiW9QQG15enmSCAm5TaLRfhW9r9PVxzLCBMnHlVnvHgNoaUBnhIhEVSeeuI2n
yYKQJUDIZIpn3qLGa+GvjGbx/reE8F9473QR9gPU2lzXDIVdIp7PVRaJ6zPAfVgCqraBTwJ9VPhd
785ndLhO4WeJReWh7+YGQR5LJY189/zeJEW2JGJz4HiVCVs4J6js/8/m9aG0QfdVyHfdOA04FgLh
HZfe9yTGvozoGhxtTSzxw+PsKa6szQaPqMg7S9pN5rHshTGU0+SajJLUH46pLG8PTgY+OV8+7+2G
yyfhQYQ6Cw3AQjjk4tDAV/jzN0hCS3oUrcJT4qHZApS4+hqXmCoKsSCdFNZM2I3f+4IOP1cRUbb8
hpRim1x8JECLoTvXU/6VjqlUJDLUrphEBPdRMKGDPslMouADkBuVLjJQcEqacWgzmBkOry9H6WdD
2j5dJldRwsIP/zyNwWMl++2++zdjvMWUIcFcuyjr6hl5cjMnlA/eIPDz5tT9WBcsRzf/3ZAiL0LF
mZ+paFwt9IVBIL8Wm3qzz98iq4OWWJ6WukNGxfLKYdqv0xXZ4QL/3hHpj8GwLrPzZurc5FJp7pHn
TBd+JSJhTMepEvzC/q89F7uoaGuR+67qREpd7nhgGr6eJp7Oct2MTNjD7C82cqY2ykk0s1kf7Xg0
9uGVliC6gbw8fJ3ror+1ojHtuqg1dI2bIW40D+5j2uFeWATkzPAOOsdvz5LGBnE7z5TlKymOGdV/
dQndp17xVQLaW+ZeNbqR05CxGux2BIIJu602gWIhux85Q0fIXxLvVgOHj/B4vWtmuw4Y7au41dTV
NdxZikb0Mph8gWQjPk0AyjAR+1KucHJRUkF/oVdP22sgEdvRq3yOflLTq9oUIky5RUvJkKm/qawP
EXBGT4uY6ltplFEhYB3q8lTVnzZmsIRqiTlK90VPx8LJXVL6Ssjnoy1u8bQfjbuhx1LojcyVnBei
dDU4gFXmve6Eevcck0c0NQZ5YBBOykzI2Y/Yxi+Y9SXEWdA4rLFFmvj3NnCPEl2OFQeVUr3hYp/Y
t6oqq+MbpMbaiH6YAfy/chtypDDtwTjDGA3zGJ1rn6/IEKMHCiHGiAvmUR+mpmJgzsggI/WoLIwZ
xRY66ZC7W6J3vAxbe0+v9ZbEEm+uN89Ez6wc4YZh2VpTlc81G3NaODk3pkBc80b7phz/PWnzg7JP
CD/svxzdqNk/iD3+FaraMLAte1smK1zCvkEDDM13czRbtKEqW+TzRoJVdfgvuNeuhRS3XO0Krl92
MGW9qRSDMc0WSqp3BLpASxHj0HhguSrR2+S/weR69cSOaW6W0NGuDo6jyr2b+1NZvURKaDlraYxg
XEQtv71uCCPbUeSr6RAVP7SOyx82L0421hOHdNfC0w8/O/YuN4QW1p0hTeI4NOCgyRPbxGHlhI/w
d4y9AToxgKla8sUBLzuabhpFe3aIxuc7xjiLZXIv5ksAVyR7ravSPC4hSCGNar0jV+i8S8YW6oIp
qY720FHB9Veu6fLhxzuDstz7hRGRPeuU0XZUWmgr4R//9kavIwbemQZCteyJATvdqM7MyUaDJ1n7
DNIAB3EsyA4VCpVtiHN1b26ys045bhXeD8qtVFGr934iHWzmVmzYvtEsLUjOFAflzGrklCLEXzjt
Q+j69rueZIsdI4N10rlSJGU+Mnzc1EeV1Tweo8lfGte/DmeA6xrj6hgR51ERvDG1Dh6fSbbkAMGF
BouZJTJoTWW9KDqJDt1gd1dcOJ/rNfSHgg8o7IdMDBp2m/w6N6EFpf5md+/0epS/hiLF9w7WZ5Lp
iBaa6Ki6as8aSx8by3xxx1m/n1PPwGcQuD9uo+knI8/oL3lXvsgyQF3VQ26yrTQ1fLCiKTSnhRjr
RKgql9KzwdF9U7wFPxNQI1yq/FfWPAHLT8ZBsRiu2CXQ/1Y6X9JLwaiShV5p8OIpdDVltT2AL/zQ
eQ9/W7PouICiFwuGZxTyPfqO+NxwHTBlF1z9CBqtEa+k+WzP2qT6DvHK9tNgDJCsE2gAMTCpMHkQ
3NCpX7hUBwIPdkkzKHmKVNQ8hSj9VvId8V0Y91WFvyiXUgSxkZR8Ff571OrX1HSaQMgVH+0IP+ol
fHpHk9gZQML72VKU4+tr1PxFUDmLz4BxFMpLCj2A0bfhu+L64wYqN/jWeI2AhRCJhb5s7/aqT3i5
fBqJRhuJblrFQjym6OZ9d2TsRDi14v+2pB1gjeLAbDoEj4JQCvGzVAtVyIt3PYUtkDvKshKmenJN
wHR8KQZv++2IBQPj7ikndxU4FGQCWPksZR7uPrNHKV1GRGTGtZCo9eSTp0pqCK+FPsWbIuz5jmjK
QMxiZezmQDJOaNIPM4NSyg6mc+1Ut4xCx1OBTa1md9r+SkQReIA4TUfEUQ0S2gtGCWr9aieyjMXZ
p356njs5vqCsjAnB1uzVKJOzp2jpntMI3V8zxnQqsZNPL2EeYwlt7aYdJAAWmH6NHZVjrD5Hp2U3
9SqxiDD4KRFv8JPBzvwMCd8PX4PkQrCcfcITsPoAm9WWh6cFZMpySQvrDW6AdWgUmZY7H53YGKMY
q442VqArmFWsEP6sug6Mt0RfzoKZM3qtx0vCHqxcmTGLDl7fKGw0tiapRjxuTzioqpGnclP8GtB0
mQJPzhx0eMAL4SjdZKTtknqZbnYFNkG58nFAbu/HEXK3bFAG8Liy3AHLoWn8bZ9J+X74c82LBgck
k0vdMNtpg+96q9abwPoHC5JYmjpEOcfSI0H1LIUh5f1qaVsx/15kWyFzpDAtMekdGsWO1W6JAAE+
w+RfaqNzL5ei5UlrfeRE+tkp1GOtyUzQzIKtpWYBA5j13xNPdToB5nvRs0pG5NEAsKrtkiFHHYjS
DfJV7LC6HxDG3B2sCkUUH2ejJMjWW8caBIPJG/jJvUQRqp2iy7AUlVlpauB1WM8mQunDaIZ+DVqN
jDV7FH17c/qTLvA0t74Wxbwdr78YnMvB6jOu8xJKQu/7ShsRrpNPL5ayIceoB7rROkbHi802snf+
G9kAJstZLDG6IE0q9lL7KL7NDGsUOl0CTOcHZIDmJRHn9HmDMk7ti7I+h4c0RBhbo/R1NL04JNT9
qF2tuSXogARMb+a7KhMAzbvgEoDIeygi6glo1zNQG73he5NaFnyl9/796glBKcCTACbMBKz3AQny
Z1IzTUGq8+YYvRDGzRof4KKQxJvBYq9Ho4iXxDnZBZ6oJP47bQBcToPq09RXu8ogHZ9Lu8iQgRag
iJXcYRqn04kU9cgtz0Svt8bf/fYHZOvyBfLvCmozQUahL4vwmxQoRvkjOcNGZCyKJO7Z5J4fG7+6
UTkgCXqqxdgNmn1rsxrggJ/6HRQBKPjUuKRm2vqWCtpdMYoQ6DyXBOAYB3bRUrpRGzkRj3FIdCq2
/CBlMU+z6IRLLWgrmOdTYCVQPpf2A3dXh2iO4PpB4Qto5RAOuWhFbTCVVRXki3MPH+MHV8FG6hay
96BeqHmNjMfNvp8JHtr/5x9RkmPTwcRJmx7rpxRy7EYBvfw652RU8gUuLh4hZf6bvm//vfjAN5i0
AHG32Fi2twph12KGdmK0x4Ww0wcGL3fWFCFgLPu2goVSFjk+Ls73QMXmXNfeKu2hGASzRv6w30iF
MnHIT1flNNZX+xA7WE59m+1kC/VU4pQD2VTe4yQfpksnNvUb0g6O7WrfYtdwV4w86Nt9NLmj3iqq
Vz/RmYEQIn42LChFEqea9FdmP5vbJtjq4tWIIHBr5sKeg/Io7v7b2rZIyrmLxMZ49uva3UcSSbOu
VWCAJlyJkxewMSk6cfIeCb9+Lfb+DCn+b8uUAbyXi644W3foWcAcQqTv/DCahu2IQDi/MYGTuMZk
X3u6DfBCx6ikEjjNd/F4Xr3/VKsyJGgf8kv0gYuGViSzHv56niyVA6IA2TT95WYgDu8BMUPi+XdS
25eAjdtu3q3BJfuki5YtnuRUWVLKp4B8MMmnu79hJOCLhQBX3vlZAWo0+gGNMqi+WeiUFq7mnnS2
UWQrEuFKdMU5fYaHGfZS2CTsYEMEOSzSF5vhbEN+/+MYbPVNJHs1lBXhn/D3UIEtn9vrox/eLGJD
NZGlcpseyZn1VnisfmRAKMpvkfvmVsb9PiifDB08xahP0tMLOxkob3orfK8qI2q2TL/8bhPxysSb
WCXgEGqWKisJQy5ufss481zIlnpqr9AIAg+INERYZ/kyLvVtapgTlByc1c6Kd1GjDTYdLRo3JSrB
DKH099qNYwLg6HwiKuTQzJJny4OpkdL5JjmqRrsJ6FaEyzxAj/8aHYkutVvGRCaxrqYYEoozq3uq
N39bvX5MqWlbn7gIGSbkK2WrMUToZQSGjkSiXZYexf3G0//FhHD8Ec85YvQYPwN9Oust/ZLV/uTe
dF5aEC5vw1RsxnFdsKbNg8fXPEVpvUOedq7GswYlB2teI4LjPZe+/FocgQ2Hm44R1j7rmGbTUxnu
UTNY9nbtB43U+STGeLmuTC3upPUS6w0ISjN6oJCQOo0bGehKtT+imErngroEkmi0Cped92moH6ZZ
up8ZL4RIOWJNfDBEvU6n+HQ2URFVx/FFXxQLDZnD4XNWfAh+cyW1wP9mYaQQUZH8OfluhFsAjvw5
ePZzh/tMc+TVfpnWlnbT3LITkOG2490RU1uXtWdnWNFqgJPRRQN3mcMR05HpF9czM50X8JOR4NJT
iVGc8u9XabS5Ta0gP/f5N+T4rUNqnWZ7GzvNOU6KHSggkiJKBfx3eMNjzeIenIYPqFwI4wpCn3lC
T/ncVK0NyLGr/ta9hiIHbGG27tbXKisw0Yah3Q6IU0dnK9HZnWi8Hvfzs9aJtrho+a4d0NzOKSyr
rn2Y9Vyiuq4k7DZh/e2SxTY3R0i/XmNO8OiPoNTnWSoogVqAauSPzPLhyIt3vbQEJyHqLbWL5bs+
gCujrJNneODT9IWxk7xdGYFU2bCkpcTpPH2IXCBepBiJCHSqXbIRBncqyaDapV+WVBxx6DOKXKUZ
sA007dtgDsDAZ1qjiBzvtzIy2sJj7hN1nVcaRsr6wRhTykD41GHwoXR8fd/9CvTF+RNDlHDMN7o/
JtsMZPw7ToVHZHzwrIg1Lx5MtNV+V4b9Lymzt97CHOKmzRMv6f8zfjdyVp1Oin6nod/a1RiJqhcQ
JIw38/8019JGTwmf4TW4B2eq2Vja7vOL7mzbX0H2V8e69ePIJ8jevXmcb1J/fTzi9P3JmeHOeqhv
n5YdKJfLKfiitM4NVwYLK6TjVDOx83wsUBvcf1k5f808NBnB1uIyihLdMHiLAj9lEZ2aiMxGouWY
BdIP2603HNzHt6dNme0X39cctXD7a+8F80mUI3S/PacNkROA0yMUbC4eE+dluNDIPPM5xSQCks/J
dQjJGum+kGMtpLiv6etOhaEkQ9WKbrmZyYgV+RI1ynUHtFL8vDFeJi9lMtOqhIjE4H5JjB/qTL1Z
jQZcJOz2+KphsNsNx4s5j1SKybxZrDpl9gj9vXxky/ymMkYD8djZ6K7vQbBqEQ7Jq+p6/2G+IAk4
cEEAjtyrzZ8jzhXQhSbz6pZIpDggTL0prDEMjijQuIfa2QwaelHeblwk8jypVP48P4J0reDgrI1o
Ss/UkzT2mZ57zcqDYBP3EUF2I2s5Sjpuo1mZNjDZ3vAMIyTOFg+3mFe/63v1H9aPILMb0Hzi49yS
lobiQPxZkgdjwGQc5T94vvPR3UpvUGi+N1dbmO+oivrIOHxLLQUnzqQ92RQp7UYELD9CsmwVVoXT
qoR+L5J/0t5t+8wq4k/QA/y//Tzjyt5LTH6qAt319KmuD1lCRutMTWyRab7WvHMJReWcskPX99x4
Aho9TQXHA6BZA2FpiAVExODcwGm7M47t2cUazJAGKEYlF1jbe6k2FHJmzln5W/MG4xHVFD13iLiX
1iXnHCSfwRm01QRtUWq+0skNyjD5SZLOhXg1jdSFsYYPTXduZHDnfORXlvuRXW4ox2X55quCnvbj
8paqGAAgb903s+NEEKqL80wXkvOTbSMYIHFGVzMaNTQoc2YN4SZMD4ftKt1OaP6k5+vps4fq5qKi
eVzBGunkrqVzy0PQv4cpzn9CM+tXNmfA/TsWIEoNJHHW78frN+3b6b3SiYI2vWJVOwCE1cZe2VXq
xlmknEw7A6L9T1dS8OOLIDefRY/ZNlj7h2rF9tkqu8CLkjapIYdEXmq5IO+Tl8sRW5q0mKMdHYeV
yl78gRFpfWv0Qv7aTFL6ZpJVsDnNiHLwMa72Sg+cJ2Tq6nWiwvsU5/kBOObk8Kihxx0h3qyAygXc
/YLF0TiVehNo5Mt8OEQAXUmDdO18EsZW2scBoXmV4QpvVBtQCSD3vLtcjhJJBzvLcmvNM9aocv+K
08yisftr1z+Pna+pYuzlcMehmW2gAthEvwzH2crkZpJ78qrGgNGU38vCxVvlhr/vdy4Qhxn6v80L
gzGAJMLTvpWSjXthRTjRegzoHu5VTC1nwfRNIqUuHQHLBydWP7BMEnvdwjN3ApiS91QgwWCpXdRB
PkfOmd4QTA9h4dJbli2sNYyeDTv5m2LiXQf8LaKjm2RIfVXbuJYYf+o4e7cuVyUeWOAiCdUTT7oa
fnOehKXaWR40WkDFiUCMfCGJHFlLYMxaBUvkdNBzkm/cd9SMMFapqMtcdn8sdnH06SuurHFiaWaG
5GGtCKmNIhlrqSfP7ifvyWKc9lfDQmUz4voQfW0EXPJJ98XNzTgGOOlzZBScKW1cO3aanQ9O348r
eoDG+GDF/l2kh0WrjFCHBCmeB+t6B/jt3WiTOrfe/WiFwnRZQjJatuQ7ivJolsSEzr/xsXp3M5Sh
6mCmlQJnA5WxBXO7Ma9CEV76gFhkx5Yk5TTK4OALUm1Bo7mYyJgEUKKG40DnEvEd5f5IFjb9xyLO
2wL+JG27OPUIB2IVvHItNdeC88NBpuGob3DNIVuTT0Fn7tJq0TgjTbAwdytjzZNlQp0nSizpD12O
u6QSrWBLfVCti9hfJSP1MvrIJIXOjLVjtjAYSuygaYrMt+SDAi0A2XrEp/abqHrIFWV1dgRcyiAI
6iMxEdAbmgmIAVyk2ByxDiGPW0Uqbt1xC2XHGKdRebdAO7unnoyoWjWjeVqcwsp/26LrwOBarFzX
+i9GPtWBcrv0ASRAgd3CBw+zCYt6KpZ0szhSJgdj3hLGgXuLS1dZ2Y3jkdOEztfqTOXNgkoOGjK1
CChw1wcmkJV8xREZ4UIjJ6IfaPTGHcgcaHM47YoFjrg3Kz7/gfxdaeuEsUatgA78llxzGgUaOqjf
3Yoq4tRtl9beztRwCb+3KKk08aWjPKt3ivK42YISBnXCb2SCsHHJnFJESq6hdIqJllbS1/ERCkaj
KI3xJmNk8ju4oqb74ffttg+Ra8XVt5Uiu3IgiRxqHEmV2+VvwqndYmKkTjfbQCVyeK4PFtTw0GR/
iyefuUHVjYqsR1O71pLiMZvOgPq45orj0dHdyRiOs7RU9E8C5itsw07pwvmbqnKHumEX3HQeBWwu
EMV33ckE4R+IVjnzGidA32Rpa/xuVWTsajRBz7TVk3Lv1P+fq72CwZ69ZbPbmoxbQiYStz1Jf0GI
8WGp3QNXlnpclyVSqDHObF8yrmgVfECDjWAu+AhGvdXatEi58VUuLJk29gOzSqcjZ7uYtYpOwKge
mtlItMO5CMcnHsQUuyJGDsm8sJHD9B71t7nhZgfCVfMSNqVVbSjv7HXr+ZM0UXRB+yZmQWsLRweQ
PJ8Ft+drXUIS/JLn7K+wNboOBnAieIxKmiXSSahMUL8M7HD4WU+XDh8OZCreyW4JOJItXp3y4C79
xuQbaqsdHUZ6cRCLn9NyxkGc/AhkJBRcR//aZpHB7P6X2McpeANq1FDXJTTdT7K/YyKJfMEmsLAu
k9YOOv5Rw0QUADpXlyoILc+ti59cvwg/m8lj4xU5HWhApfCbdvm877W+802hh27o1znQNDpbvRps
ahZEwTuLPlPkOzFGtU8Alkq0PxaiMa2+W92EW+1FGg9A2W9mBMi70PfhjgLw0cCVlf+a14SxAhR4
am2ymptWhQc/2foe+z5Ob3lNQL9Dsf2wDsqYRNPkcD5tk8cbnaq1t+FLk2wXXGS0pKst8iIUnM9w
cDoS7ptc5WZcwlEEyR3MSLcX8nWMpKznnzeFQxqLUWm0MTu9KYcHX4YhJBBJ7j7EUBSCMe3MjokY
QYKkjl/tjDf273D+ToLp5Nwu6tTojfzl8djsrbvzhnCoBA9K8ofjTuQz3dZv2oOtyIUo/mokY/LR
cTevHcL2VI/taGgTJASLlsgMkBkzgCJ1fD/xWTzCsVVzwEdhCGSX33IxafxX7SWAEaBkJoLvv6S2
eRVrgxFDb/1Bnd8Jyf+Lj2izcoMXmSynZjw4CwpNwxwtM8e55cu/U1VQVpuR1CMq4OihAx0IgSYm
a69TDxpr/ZB0ndmViO1g/kHmRMwu5fe754hB7BYm4lqmpZwdA0qELEfsS98kr83T9obX58/mZ0zQ
ntamOA3TaTCTyXQasdbPUnusfMNqqHkCekfIOGf9Kb3S+qIOcxTefJHynZnhmEg/SLNSR+Ksey0Q
OmArFDx977NhieB1obKrlfrQzn+T91L56nvuD6qyjomA8psREkOLin/sPJXgOqnJ5agRT6gP5GEo
H1C8VQiGQc1DFNcPa2uR4hKKFk3xMwdq8BhcH3rUraejFDjEYv1X9zWXXCxCLhPNvLHCekD9FpiZ
fXEkhQKIwZ0+yguldi7i1xVKB49JxmGcfn5IeqtOigNL1RlzB4k+Lf99SLhHwnZFkEd5Ah8pO1vq
RTOpT4xrCDKvFU2wuuIRAdIKiDk+B0LZxCc+DjtB9Skfd6Gbip9/88uYUwHZghTHHHK3A5G9FYpY
XW4GlXGcjG/0zQhgiPzTxaF7NjNEJ71T3R0V0K5YxpHwLncUfkApJEC76rXc2EBJZFAgzwpbXZOl
4FEugg0970sECEMtA/sIABMrmOWYEP392NgQ/x8pw1YJB9F/gMs9tp1vx/bVUHWYpcF7Ry+z7GAK
1lmq3cATvtWeb1J2bVeUJVYf5JO80aHfwrMWRRtbxvkC1Mq/9YrtS9OWCAb/bQG3FUd1sof2z8Et
5tE2vZi4wK7iACkW0z+SSgznWYzJYIvft6SexqaRmxcus7LsGHFRZd1OI2YlDFPSDJlVg4PkITBK
+1VeXrNzWDUBKg0ceYPi+54IMZ36KqYBBR1IOBUaW/0glbKhwS3i6+G8kiGVQDQXoZxf9uoHH5e6
5n1oR/UtDKnYLBn9ji1IU0uabTyffJ7S4eMDEyG6qYGEHPhphnhM/NjdBOiqPf4Zpl+xvSzka499
CdYCnwo4yD64wLlHmMuTrWgV9rLhdQRAow0KHHCr+rFOBbSO+Poo7766GgJ8iPxhTxUVc/l9xrGE
H2Y9nC5QGWRFUQya28KuaiakYWxjpGG/WLobvJJscjf5uWcCtGgGXE2vvMUlK6chnGrKoUSL00RZ
VZbBR2TICK0vloD+bV88tVBaPC4MNbqXgcKPOHoAFwcvmeQPpHICjre9Sn3sTKpjEWzU9WkoMtZV
qjM8tRxSbHzHczFIB2MfC7SFud9o1xzSThAAXgdDte8wE4CscjE8cEGvMVFUiqC7NfhHe7l4rhVx
pJ4uOQS720HqbcgVqV22BjAmF9oPF8GzBCjMyFoEufMUoYuvr90l2xhUKnOrljNMwjT5/oUP1wpE
yLi5c5TjLCKEMc6C4Y8HRZoWBz8JEsKw5CJTXbUuwZEt72etmPDyHBy5g7g/NM50Z+NbicQtdORd
e8V5f1zn26uML+z3cAIdbKrkHLoIEMjt3GkC+bWM29CThvhngBz0ok7dWEnveAZ8y+GrRZYLfSk4
WmbQ5MbuDRWORvAB0SzI8zepAHFe6htpyO+m4nOcU3xncL14Hz5QcTU9TKqR0uQDTwhmbiJzMCk+
dB4usV2O3DdMwy91ct8sVGvHLvXxwsh6s58rWhXV1PwCVaZ7pMa54G9JtjDrZHGeIh7zs2OK+rdF
pBKaEE/859AjwQYnN/X/MHthJh99mt8eZ8upKfU4Mab+rbOM71wG3kKr0cn6LfAYugXC8j1uUwy4
vOmo9ktPpp8438+3za871Y8JTQN3nmkm5tlp9L0jP/6WOcdGAy6b2IVzuenQx1ZqUmSdYWnMTZxf
j5WAoRZY2Wmxn4r5a9N8ScUrnvXj9fMUd/khXhHwdTiJGKc5nwFbDmOq2QXugCAUSBl1/xvZrIPZ
jJ/AJqjeEnco8LvcbQgZNXclQZYehZ7sc4fyWUlgubcVyRgT/0fE0pr4YuSb2mN8trXqYHbeKybR
voZRFILZrLz8szPWlSM3GuwcpqrjkDlMhWg2uG6RBJhQHefp3eihGH/sljGZBGn9Xjuj+g8q6K0F
B8xBe97dBCSGjcuJ8thRH1b0UDJ9gclutG1wqnJ2Q6+UqOXzsn1B/vHSrFOeZIpumAIGmkJmYgxR
pBmJUY2UcxGWDBGU7MlPcqyWBYJOqqUzKP11Rd+VDjz2v7GYc3Qk10tVSMfuZQIQRdWU66l7G6NM
zccZfRDlO+TsFCWyhV6Fw/iRIMl3GEOhl4tL+s4TvnGG2nzs70AgEY+nFQzfdEO5p2at4yED/niQ
ZHy+iOmDpsimdo1Mud1hPtFAYa8FFB2Z2SIeO5z0Fu7y5n51l4SZSEB+Fzp3fp9cJ1QS4u8C3Net
JyeHtOxnqpAFl60kUBlw+rNDO1SShT4qzVJaWYItj7yTLHINyvGjO+or1+4bVqbSIo0zDwhh6gfc
0kivOghfVnm+T44bqFkV5Vku9yqCdBcKrO4J17tlzIY/pgpuCxUdwA+upCjFDotyHO5WxgfJMVn0
84BmC3OCgMpxugLYeObGcsKEdUPb9IvnOzexULUZJ16ATvDZ6Pef0LGHvXrDTro2zeWP1TbjMX0H
oxZLxzarmk9I6/cT9Ulet0KdFLqNU0RB/xWsFOUQgk8cUOHPz8aOW0P3p7SzxjvzWo0BllavUUcl
X57GuJYvPb3nmKlosgQAcW9c2ZhsviJEMfgrk7HdgIkLZaNC1GRgdy84Y89S9teA3xs2xnTWp3J2
An2BOA04gZcCURMYueOYFUTH+V3lbvojGitSQtH48PXWmGwoRm5xAAfyjjvUU3AcEQiuARDcpGdw
DITB6h0pImD7RBZ9sRK3wXWNWeCJEQZXVaZQ867h3L0gKVqtCEoOZOi/kRxx3rqdMrc9os29s2aE
VWiYthImWzmAX+G0ZbbTCvfL3lNdLvWnncNPeP3FRVsL5l5JcF3nIbZeTXMyWiuNd7nq2Awe+huv
A4yWeW2UNRRuB6zn7ZAR1g24eiJht2uj5U/FGFEogZnu5YsIXbBLXwv21ZFEJFGQ8EWt6uIEJ8Fn
eea8WwdDNb75Sl3WyskYTscisTvwTn3IxvVpBixx+yhBZG15RmWWsv06YROJ8Np2DUgHmgFLYq6i
8V8g4JoHFbht/7/yAHqmn7Mpfxq1sbem1m03gsKp/Twuh11PfxCqmFROH16Wb1ZA2ctRtYZ8tN9c
a1xZWnXOqpkSHgl9DmJV5j1bqvjXS8p8WRWptsPZq/ggy2+pTWRp6GrbpvVF3qab8uGstXQmfIVm
cDdKEyzvgK68Ic09if33U7Ftn7wnJ/l3CQvVCqB/83PEsAcLFxKJEfD+EK6i14O0Qc6PDacGTdp6
I3j6R1Mh7srwWd7tY2KLJJY2uhdOyOAUU4Z15R8z5Yw+6utZak9aLf5KTK1rwg2BnjGM+yy6qjCw
L5uzrbh+yLoc05iJYnQPtOccUtYlmkZNhFjMP9zRR4/WQ2ggBLvMMxfm1RTj+SmEnhSVrSQJPvI1
voTg6jWW6v4ekAL8HL3uJYM+5TKmj0sabxMK9CoS26X1tsBuX002zEUZfeS3jOHmeyaU+UlX1nLh
uKicEppM378hD7m7PvaKe9wnGz/iyiJfAAgTev+CMuFwcRSzIWKLZ5T/10CDUU4r2LmCvdVTSiEo
jNQEuqIwWhVWPehMfOU2rC8z2alrwFfqkmPSEb0xeHzJ1Kd4Gl2BdUse3aClSDTkyLRSmGad0lVK
6xoOCmVxw062rT2P22W9iVLZ5oG6vw28W63Z0LFPivUy9vyUNWLvkBkZ1Nxi3ATaxOCiZKKXqQ7q
DTovXptpY4k7MTFj/E0ZBccIzXyXdI+UCARqUwhj1LBCEHn6Wfqmd5fsryPlmsTsgT0QAXoRxPxY
YeZrhoT5aJqf/pzKyzh3z1PocKi75LxNjcYP3C87eVhMIAxKG3pI/Apc/inMw+vQn8Z8DBfbQ2Ot
ajKxM8K0IxATCfpQ6nL5/Si3F8Pe9gjqN1Nw+ErQSryf1ghsCsvaclkn+qwm9Z0mxaCa02EabX4h
ojkIFvWEwfRlKSaqJmyDDuocv4CbzHmjWj9FG0F0iCatFWWYTvhC/D2hBZA5PB2eAukkPt3Lvnvf
luZPnDhMLhyA4fLGOJqMWi1NAYVrF+BnxTrgJ9ScLlYIK3NhZtMdvTya8EKKq4W7pxxBKQAr4dwJ
DJHMpTdhVLJ+MQ/rBt41zp5jUUUUw3sVWAvl9qXAFFkqtQMpdhzGDXV2L0vyIoPg4hGupcJ+wTRn
ntLNOfCNnDaAokghah4eC9MMnXHa9VPSsIfJwvRdf65oAvWRf0ZCqQINijSea9BTYuVsgcpiexi0
5yEE3UG+NCQjBBcQzlQriP7NGaaa7ko5J4fIr7bHzTAI0p90HQ93DxmXpHgcJF56FMQldn/6TVwz
rdv91rM/F6FrKlb/omFJktM4BRb+L6e4k2mXNpTtC1hV7t5GJgAKeNyN1jVyhEUeMDTEzNFzdSlv
JjE73yd2nfP9eRAdGqAOJd4NvBcVxiuyj04mwR5qoi3Gi/rgBe/gpSNcj8QwrILXHSb5eDEGyk79
zhLxiuDvMRR8TdjC2T119vwd1epLgdRGO7KHQJNAdm+bD0JdzQQxaaqIu+kQ7vJl9e8vI+COR+L4
hAZPTRgZXHlDuSlel7lSIsEhXvwKefRzPiryPyFWQGjJt2zQ4lLzfePWjCaUXd+nxS3djLIQkmnO
hhNWufbRcUKBOU2LtFanI3oAQycmL2clNPStNxsrkEJE78HtPAGHz5hOrkmyqzjv0jAVBlA15g3e
lq55JHELyIzOYQhguAzki8KoJ4q86jM11FEQiEbo9hBxDkmxsw8/w2E3DJOyuy0MdMcoWrwCoQ78
8Eswj4+srEtQkRtRUQkVQuoyS26qBTiAvRDoBCBPJ0HWFt7LpUulU5sI0f5wYVtZLVg61f/l3rY/
hzPMroGreb7tyN1aGOuh8N0UHi+cwy+Yt0VTM9JEflnz48grShbkg9TmHCtotoa5HZjR9Gsk1Rk0
YNQjjag2FW/onsXWf1PZCDNPIqAfLFcR4EgMEnXk7HwbcY6XB3dOc2pIhMFdQ2vTslGtkCPb+1pL
bKbU0HUrH85AJp2s5tQCjqkxaR4iuWjqloctwAY/hIatys4p8tjJaGrDBcQumVnXoE+M5oG+wJwo
RHorU+d3Fx7rThOZ1E1kwLLgu78mugKePBoGEXSJypkmmhNndUcTEXoJfIzVqjlr/a1OFZODdiht
wMQbRL3CjF/0hNNgVfXrGtChabbw7NYTSkXNyArj7UhWtAh7MkHcC5V8FMoTcqN9b1NRJN0wd6u/
oMsqNh3XQL6ryrwt2rl2x+BqOjCfzN/KCZUFK4NyYxxp2NAHzymzg5XhujoOxtrXHCte1mSk1KCS
lpAfunH4yMyace5Fxtk5TDb4Uuhh2ccYoqEh8yQXV2FZeaetS2wcDmtBL+/Z6zRgc57I35Dm3rXG
q/qvKAe+NBVZZe/ick0VWdqvgZj0hP4mXJ59/IDJFMYVfmCnXT5T/a4t645MT+tT81c5M9QG7U7e
qN63KoU9M9EdggfUOsWEQIUTI+hNXPf85qKR32B8z1+DoqxrXn+/BVJWjrs8PGi6caC8xc4hhqf3
cWzfvsUZYInRmyjK1X0Ztuels0OHsQ2r9ZIft5osLX/8VIK+86bSpVzRGoiRyCITtkyMbHJC+gUX
WH9oXUkDoTX4lJtydhtJL2OkAQ6MlbsdssGG2/65XD4WqwA+cXePPd2vUyrX13cssS9x6NS8oz0e
wAF+SgpfVOc8gHn79ubwu0PZiC5lrnLGcHGxs/lSNdOws6Vk/tAhoLGHBuaR2610GGprE5zol5bS
vuAWzAE757guFeKX4RYMd7GwvRo8wpxfPVOpSzzO5Mnah3lwla/TOdsHCex9Cd9C6NhdB7f3+hO7
yDoVPQI/SQubv6crbnTeu5ESlsrx23P1ChXwOsbQlD3Q7qjB3zsUcpy76Cj9iiJR1Zmj3K8Ly5wS
RTM5IjlEZFuEeb4E8SGh4ZmW7HmNWNId6i4uCl89i18OpknBoaNIFokIVLWY4wu2gWzJ1yM8XyVR
YfJLy4QGEJVBgpQBIDK3gFBWhb+XTptjIIBJTswrjcq9huweBpS+dyKxnluNocKfWuyXCnK/1pX4
fY64pizrhBae97lFJR24oXWNYutQKej3pRze//6z86wFNVuPCxxP61SBUqa8awj24M2g5ZVhP7Lk
mbQ5s+fQW5D1XdUm8lEfxjrhsP1/uvWdeQvkitKp7Sq4kdiOqfNGVL1E2N3WCxbbGgGTGkG/d7pX
ZPOJ2fl0x+xnWz5EN3jD/rdWNN1zXJjV0ORS8ycRfjnUlyWHfd6wrNLubDDMIFB9e107VpWnGxBo
NBa6V1F9G7p+VfAqYn+KicZcug4QzlIobdOFlot+dcy3PKemQigI5qhxgrMV8SULxZvm9q6Ma0Cf
rMOz2F8tj8Pf7+s/NtClu4GwcVV/vybeb9i8fjVWoR6GY1G9venDV785CAFyLMnde0ckq7Q+AePS
XphToKBExFIYig1wXswfgn0HcztPnhvP67Pwqpq3ro45OFVBLLDTNsjdsnBuuOWp+mut/qWtFkrT
OjmYXhYJDkyc9hajF0HuokNeOPOEZc/ga5ZKJZeQHypW+rXI5J2caV4KcFSBIUHh4qT2eGQVo102
PTLWe3TrFfflZ5o7nUL+kU7e81+rVObE1qBV1arA7nXpLLvupALOtuJeK5fOznKACSHRnAHDIRVH
C0kL6edOt3Rb4XHyqtfeacQkwzCwXLl59U/vu/yQHWAj9qarGOXlHvJdjZltNi6ANq1btYvoX6vh
cakoOefiJJp5rKZqf8IQmys8m7NE/oj+bmjXsQbPCJiYDPnxR/9aR+DxytN9LaD7DwfMM/KkUtAc
ueKhRRNBzR+IIGnxeMD7AD3I6runDZUZzRrLoL7ed7I8MT0gxYyF0Ov6z/88n0QJbTc7BcDis3rF
LrD6ve1wFFZ/v1d1Zy0AK6zyaHq/fWSW4ToTZbBrp+rv8ka3Q217ES5Cwecq5dYjwP6Qv+iHMnCk
hYV7BfqJa6rTs67MYv2aR2U30DJfLTXdRyOBaJoq4GxQIEMYET0N5xaSCUFy+CMrB0khtDQ94Lye
DCepwcWGLyJU54J4s1+dIs9fkTZMZ2XdX/RVxru15DfPAI2SZjEhbM+sDWNxlpi9XZ5AIARPd0t/
B1gPnnHv18ZFamYuhKQbjg+8k6h5RXoa2f+/dZpFhsvDOHGkfRkCyz9bNJf/UK1Ze22UK6V3Fhl+
46JepPUb5beg6xR5Cwy6X4EIr10vRdvLMSDvs3/QLxBtlWxhw74aWG7KZSIVAXH9lxB7DzITaOi5
tMzyH7lAZ4OCVd0YW/l1bSZvWZpIsO8nMUspcd1iiw5WOqv5sgjAucaXDB98psbhkHsOom6ZZMSS
rFtfm6VzCp+LG+dmhww/701Uvf5jX2fje3pXfUAcHxH59F4FTrUdxCSq/L0Zbr9fOs99yofDKak0
UhCEZ1359vYrSZC9B4OjH7ljh4O2bwT8TwnDxpInm/LrtEFuvJkAJcely+fAw0mR3Yt8mHrXlyXP
Uc57yRn0cm0F3pxYgn91zPTfS/GnUOs3EJIsCAVmgsM34atI6GkSBdtLj3mPVIUOOyX7NHfLvVsO
SnGBc6c4MnmiQaRMiQE7zpkE90aq198K0Xumg64DheSt3ug/f4T/ZfNzeni2WsbT6f1k99yPN4NN
cntUft02z1S7YBGdZaiBNhnmniOR2jmuQtfLD1z2/64gkQZPhdBxQIIU1FXRtJYXjbvwX0HIbGlu
IHmYkeFMnYlhk47OwOW6hwmPPWA01sgsbid1VGlh0lqCseT8A5hi5koeqWAtjBPCG83IAhjxGmjU
fFYR9tyDDd8Au0jTQtL69925O4+Go4pZaiIwsPo9bsj+Qy7t0dCipMrE8liKl5xM02MJbAFacp/1
pjpiKKVNwR76syA/AJaH7pgjmLXQchK2wz//4Vlh6z1U8/DUQ971tyrv4MFf9dNHmecFenot533P
dAwYxbDvB/7LIaJvnW64MqYf5upKSJeV/ZjJhOWgObBsOEYD2OEF1mkPeHboIuYwW/tczUiRJOnw
hlMeMUs55tdK66q9zRILeQhbN1H6f17cPdSrzMqP5bDNw+QAnKLKG8YMs91ABZY6aTf40CyqFzGT
8t4qn54N0yYy0IKOsIfpV9Us7A1lqPf2dAfu2yn8iPYHm2aIKc6CMu0HzYupQPOLMNczV3eTobOX
Exb3n5DPfoEcIz0kWD3HgEl1murkJUIybIISx7ZkcCZ4RJHr2MnewXkvXmXbjPKnoDK9qKw2Jul3
D5gHFL6QPTKFW3vGyHTN1NKNW/EXjs3DULTH5B5Ma7j6v19qeKEgx/SYgpDKYJFn8TSfWLMGXVpu
ijIvpqwne2JaZMMzcHvz2gitEfGpayOrqGxxD2rDqrezgOXxAlpLfnWQpZiTg92e132dSTIiKBFa
QnVl7n+PzzDCIkgt8tnBPVKI0lsVEwQ7tD/fhI7fkoltjN8oY2AGLmOd11NNn8saBtmypmcx1rvV
dEoeEj/JDKVdOw/iDNa0bqi3b+nXiWwwSBoc9s9BpVuVyKhFhS4pkRpns6k8H20lHFa3CJ8dHigK
AJvvBdOBY6BvpaCc546CqBUaEV6FlrEaB26wI2vD/Nyl3ebWknJ7My00NxZwKUQ50IMxuuolyDtm
c6aHjdVEDa/eCrT1FuAfnnO1HS1iEZiNr4BfKygbyUjeK43i/q+yfhQZHbGzafnUq/BCYjdxGBn6
uThirO80H4XMmdxzLiRqCGO4jqiQZ0zkCPO10CZvgRGDQdTABJfDJBuTTRbJGCqBC6H9UVqXhwl6
OILNgtcxukyVT3iOT99dL6rw9G/bIZcSONklZjrPm3MNSYBfadrlqABOwRsngH6wCpILMftIvAl0
wbg5jTcOI/FDGfhR8VfFo/FC/kt0MuUV2/O1O8qbaoKj5u5fzArtV7V4AyQvQ4Dfh6SNE0IAFNIi
ClthSiB0LEW2UpcqvnROeTbWqIDOxsopFTsULsRgbHNAJ17SaI8Gufb6Js+gOh08623PRpd7OPQa
s/91hFAfKe36y9DYxaEqE8bct4ceK/Xq1HVZSK6BuayAUsSAg0SFwPgDn5L6WiYDBC/Z+HqjdW8F
wQf7ei9/AdchZtxeqNNDiyOSoKDZhDse5t9CQPcOR78lqonPftyqM65BEF0TjOz39Hnk5LCyEvpC
ntKpHdS9SvbVTgqLo/If4qQbHdfgT0TlnwVg1pSIegfUoSb0HT/x6178eXPktbSq1+2FCTAXbJ47
ydnHqW1bKvhaGoaOcIenc3YzGJh4E9NiunOoIpmW6hOMMTasSD5xa5pGdQpbqeqhqRPhqTNv5OaF
PTveXGR4nZ9kuUSk9qicR25DhzcUAd2j/2srrbaLQ1GVhvEbPzc/Sy2U62cgxKXjxUeMTtVuWVzJ
y5V5D3qiNzYD9NJwl/fOcHCf2Fn3XZUa09yuCO6avrPagBjhB5XJhl47Xt2rvdYG7ACzBkQLWfPK
GksBQQuPhgT3KQ25fDU08O4i38Nu9oQ5dHeB6gAO3J/wGO8EmX1pBa3brqpN5ZNxebj/9t9B4l+b
gO1Nsc4wLaHPi5ZPdRReXJsJSdxY6d3JfeS7XZ8mZ1Oq/381J4YyQTTgjB3dGcBOEYM/ndsozRNT
lSix14eDoU3TFhJ2y2gZJp0eCOX0Ki5wo//qh4kNmClx3GWkddsOhwUdLce7dsOP1gjTNeZl016F
5dxCw1lOsGwmw0Ty21A/DYy6PedvUYgtVE20sa+m7VOkmtqH63BOAKTKMQYekJmqLG+ZOP3zE50W
1G3NsP1/HZTgYjg+TPgkdOlUvz8VJVbxkdcl9g6BF7xatkEkWrPiny/lqokLtlBVEQ99AkmSIxAB
8sbgNXz1C1Yono9CKJFvv7ufT0Y4Nxgwv4E/czshrVTgdJt+dhvH0PIHncE1muCxMr0kN8+V9ywC
YP9Ghp+jDzYbrQ+OfoyJLg7Y1TwWiQvzVUfarhya5IzvYYm3Qtv/KGJ7gV+RqCAKZQUTkbXsGm+P
Omo4q/hjnOmvM3Jw8Mpmw1nHnKGS3bCfCKxUsHrXOK9C/tL4S1GQPLlwR/aJk4VYCtLgaOGfSkDO
IPJeO1j0vmbDQvHTLfoKcYCIUoib89G7aRPUI6NEFSQPLywk0ERJsogGtwhWWSBYmCajJrJxexj6
hdjNpsCPYtxXjb/EmUBRXnEvWIBe3aU4kqZOvcxCtscTG01mF1Oe5hWnS8HGWXznhE0kqDFvoend
EyvrTHjyfbVkzmAYghzjmo7XeEqycRe0/CNFvDoE3iPLSFA9wW0lFgHxW2P3e18A2yD1iOgiQ+J6
K26ZiU8lgt5Y9dr1efqHlKIUR4kllcBilrzv/DMVwh9j2h1LgB2tR5Vl/hgFVll7Ep31N0iS1AMJ
J8PiK8smaET6oWOb3Fzfh/vTHzdE7YHBqsPfTGfPkvUsO4hl1wulbyRM+oGYrCyhYIRBzutnpkbO
yHYLJT7M5vpzu6Ne92yzT9idSSP3Fhj51eb2TUFmLdueO9z/KBoGs+9/CkDgA9CRXdmDW9TWGlYe
u1y3hbET3i+GYPQp43BHkxLiYSWo+uPOUVzIw5weg2UgbdgcV7+qXskc71TJsUsbYI7k25/DH+b5
Nsgcdgecr/bceuuCUWPOOzB0YSh1jdT8pq9V/m7TS5sqZhUfPgSnftw37/NWCgpAwF1nqf/dvZfK
UbiI4v/LQ+K9u/FOQug/UTyT6R025qYjZehYg09/JBa3a3I+q8iTmYPTW3qFKZorAp0N9jToBEWE
zcHqogKkTdZARfVR5N37hVIrrPhn1ZAjfVodxlhjm8+Nw3oe813L0CZqBiAsfhAIYvmz2Yhlf25V
GpFWXRNeMs575M6KO1pFadbEtesxXa6vKwuvmcM+1Pr9WDGSbHKzgZcHMOA9gpcZKiKekM8PcplF
e38qfGq+qs4xaz1ZdO1xX61CbNU91ykgpsVhU6ie3Zdh8nncV2MJuIJRrK+YCFwcTw7i5pUQX3Rm
TkeT++9pt3ELF6EosW1yLxpLUP0n6PB+BZCu9I9x1KsMl0c7I2eWaxTAlW0C424MWTm532tlMKw7
TxFE1fURDHF9F4l9T/3Sn3GMi8mdptv6jOgj/ypEVIlReT8dNs/GpjBw1jf7+wyQCgswEidYAMmL
FWEfaNk9mVHIc6CizKfoz1SVK/XCUoD/Uurg27AYIoMqwfyRrEstxTgrKlZhUYij3k9zFzlu+18t
tb07LX2b2zW1hN/BZ3S4H/uFwCQiiQeztZoOW5j2zlPT4PkYehPOnUtGlD+Nf9Zzy/SlD6ijgVrk
GDEY/B1sMRA1qPrNwNE/dNK19vuRr1Lns4MYR1iojMsDKVUOka9NmU3yHSWBFm9R5EGpsEAIvjUS
kDBoROwiiq1s39lQ8s8Rx1VBc7IUooXm5nptV8G68+OhbyQ+LyVj/33m+xTVjKJMZ5jlO0VcfRkL
QudYVUI0kn8HbwmsFHnYG16mdinBSKeKm5plHiwDRSAoaPn5u5nhESwla8AktnA9DFkR0yoZtq/k
GBkayAN4Yt33o+YPy9IrY2HpshsZ8zn4pjwi/D/tuy4O292DRfpJmNpjjZIFXMD3Fowl30bNhuDw
vca1XUHK9P9aGpjIIJwPaBbeVL7wz0pztbSRhadyw4S+XVSg2DymmlGw5Jn2nyOmIUhIsZa9fy9Y
izQHWJuyLZE9K7flmsd25Is2fgUu2OE4x8Co+Slq5WHgBWhqpcKgsRuFV4Tu2Ml7EPXzYfym/u3X
9OyIp+QEvw33t6VodErz0w5yGlosndVDPM1Bw2ZfJcrMjkAUZcCmk1oxT8cRgqmHJAk2PMkh5pL4
lQ8Vh5yeGbSgSpCGABUCGtLSzHmzJlN0uehwaJHmUZNoLc06vsU7hnOaqjBtobTDNAsUFzb64wHl
an7wEzrrtZe0aBpo2W1Sxu6ORTEJ5QiGE9+oe0o4hDOtHnoWH6TTe2CoLTq5HiPh0qTF4ReuHCpu
g08A4bKF9oyGBDFzgFKlw1xZnNObvUZyHGMz+vMsfzortUTrNzrSDicU5IcnVlHigphfPCzmxKU9
QUtWCptm7u5DSYj+3RH9Bceq26+/p4b3+JT3SjqRNV/DK71h40zo9EzkcqgHP6za+pIC+VRUOnWI
dwGVVY7+HUSivAnFFqi9nu3dZA+G+oHoxRTGTbhkJoc5x7c64XZ+Mu4kLt3jIOvXJdEbtBgudyOV
+TnWeDyd08xA+AJ4EnM2uKGUy9e2JlajRFXUjaSGH7CMVGHi6+g+igdwvk1xntrOdFk46Gc6iJl2
Ekb3M0BaT1nPzTazGLXogoJLuvlKQjQoFstdIO/2uSlM50fVaCHp2uScgDoANG3Hr6VPoXHgz+xO
gMT+TUSaBRfvNp6ImMlevjEXS/efFm9PTdhrqpzqBZDNtLp0wHE25DofQ5S+O0JQWwbGd3mj3si7
d2mTxiUuQY2iYA0OHKOUBC8UY7N7XRh04aepgts3ZlHIHTjCEPe9WiqOJOApbHsjwxWR3etX5ZJp
Pg224Jqh4DexcnB/I8eWTZfpfCVrAbSYLCmJ4tqc8DNqOgxciRjQtZDmtOX3/TotzsPB7CssLE9l
Wh39yHwXqvIyeiMsX2CSMg8GYO/gWdmnQ9+cc1P2Pnxp8JOWT8r2lyqUjV9EX9edz601XST0rO3N
PlI4Ebx0+WRTC6LyO+h4QbOlFlDlzZMIYWN28wQ4VrsPXk6cP5O+YQu4rMEt7E4QvQBbYHLrUvvr
+YDdXKEBC1TMh3wQVjlNRmxWBUWPhMf2ao41AosmX9IlqVyA1RGBhgmx2Z8Oxn8CRaktU0i1wKip
dQrTN9B3MKtZnErlt97KAWq8eK7XLZgChIiNLm8FnX00kJX62+3QtgKP6OIcBke0Gi7Q9B+q7tqE
mhfLh5+lTXvv4IYEbEzHFkV+OczH4VLu2jx8xqOggYI5EwAHznJnLlisByAhO9RqY/BQa9TxAQ3j
47pbS9N0hOptdJOG13abECHzvLvehLxPI5jxa6eQ6heNaKwV12P2n6LncoCX347szE4i0E18SFaA
eEWfXcN+/zVC46H4nYkgOnmFyTDh3aw3O3yrqmQwD8jV1Wx7mPSVFhW4aAaHd1Ny6ZxXsZCW63fn
P7rxRq+j/8+sNh35M9dSQoe4nd4Bcr0dy11YplpVajt1KDsdytoEqrWOeXaKexz2H6AIaaJ0fM+l
5kSsdVHPaJP36xNkCrnbWqJvdCFqn1W2cGGbOTOpqH2LkUxCu1IBBUD02WIKea7EcjKLAu+mA65g
hpWyxO0aH+5U/U+4+OyO/XzXHLv2HudPLW7I80aqAWzU65m59PjQ7MN5Xod9F3nI6/1IMpsafQPT
Tp/mhcevzxh18l04n1T/u9mMSTXX0yQVg4so9ACqrs5LuUE7f3IIY7nXmqUQBHeZeieOmvTV8Noj
yFp2Z7G3uCvjSzMKI9rbj7irMo7kqTCpZHdCIlvsv3yv9lsIh2Y6NWell9TQYvnCz30NqQHhCb95
sI2hRjV6qfZejPh5edR+/p8sgG1mri95l1jA6XaSIKm+Bz8g6KyRcQCI188fc2lQrCD2MEO8a9/G
y5lhzmSGQSIveGtTD58/fFqvxoVH5NfGO84nJa2vfsIcGzqHiBMcCvN8P6RzLNYkBPbRx8Z9cOQr
Nu3Eo9s16Q6zW2YjjapXgIB5NXp9xwwbvVJLHZxikhBhXGDkUELEO55BCp3XQww0JxhCI5Z3KT7l
dDg+w9aZL9OuLyrvDf5maPSZ4itssusYHF71DF2Xs6JadgKCe4z+NcNV5WPObUrlNjknipAWYIXq
ynvUYRWgB+hhawSeTX0RrKoCSISvdqBUOCkF9/xJHJgDJWvWVJS8fmReY1kSd7xXliGTQxJg8+gL
f7iu05StcVDIrUF9+1PKwPMIRc6n/NepjPpYWxW5b17MXygIBixLUGEe13PI1YJnodh3Qz8wpoIs
+nhKdHRBWHaysejOaU8Y8VG/Bc533FoeXDYTg1fTGKwaIt4D30C/BS1a+1ORI4jgRviWpiZY9alg
kxyW0AVggXypiP0XdLFjPMjNeiCKvhBAgbByjsIaGgVgy/50d76xEq0zDzaaAnO1Q3ebquqF2nJs
1d0r5WC0qFCozZ4XtGZxuUX7p30RombPXkVAPAf/qYBnD53MuBGzB0mT1Wvs6LFrhRKK466EMuCm
P/U8wPYoplGRUOn6Q1rjOSvXTnppwBS7E5zvEcCJss+jTjb6XvAYPmtxMr7QtUakJ5sNRPMSe8kC
wsjmx8o9kjiTUyCJysUnA/q5+J9C5fVs+ujjKOzOXRoviTCx/hi66/BlFsZvrVr20uKu78n/UuyR
KmlMavjRjVFWRPzrzeu2qdpJJ9cj9zVaX95lHjmKTLaIkZ9bSrxGvtoFMbdqeiKS7ArGpJThoHov
g/Ie0j0l6e76HmZX2nR7V2Pne90+jKU0bszs4HKB21okc+vkmutLrzj7Ls579xZzipmggjduygAe
yUtqpFogwVcBLtgGOty4th/2yywvG82iWZOJl3fwaRAv9pxJ9LelNiUGp+qIGBkSckNCAUVWL2ow
x2Fwx43pWlnbBgZYODpDrOWju6MOm1hkwSj3h+o9hv7cnUl+BNJZDB7/+EYknHXE+kqTqzmUAoDt
yU+Q2TtLT/ls9hBNYhLaofo8MHfla+ExRHRnUBh4e7yC4yYadv7EIBsAtJ1hiUfQUpaOVquxwO9w
FCEpgFv1GWtpcNjVt+zvOENUr8Wz4JNRMkPBxOSs5XoqHAcwEnxn5/Xz3DZEYgaU068Ip06SRr0t
K5rcBBbieCe+vlxw08x6qUgSoxxYyQaSXQcm9rD0212N9/ZVwbfp0d0nS1S3OjmHuYQIvcjECYUT
bVvpFExEDD91WF6osV4WcWSVJ0IXJ38AAxeHAEQ/mkrbp1qUHus6qBPBzsEs1UepwZhTdppg4Cty
7Z+4Rs4mlPLGViORjpc65KFDiMD25zWopMwvgWB/9lYGstQEksGtmMJZQA3Q4be3Tnw/Lm6Qqhsl
CMcb5QOiCKvrkaNqlrWXnWFeZuqvGG9/J05AvT57aED2Q6Eq7wzLtsaEUP4jTWM+tKv5UrkUDrtY
bAJfkC1Q8GFZySRCRHLubcRYJ8BEYwQh6Q01lm3qnIAmkQlL+QoSgUts6KLBu/qxFGN4WX5GZ4Ol
7ALXRgphNtKOueIgtxUJSiJbbJQXPyr34HRsp00bGksjqwg3ZFyLth5ejzf4KmTTRsnSxwvjmeqq
Xs3o7DIctRjWHipHSDnxabEO1vhF65/GbmqhRiXJqRRFvD4c/T/8c5tGP1nRyTF81YJVYLqyZZaM
tstcMecv49LJKFBXK09tBxDaNHBb3Pe/ONpt1BLn8Mq3/bUIFSChUp4W1ThiaH+BqEwcrMOfuVsg
miNnytgxEBvvq0hVHjDnejdeh6ge7IDu6jrHhw+Y6nrANVHQ5MoURE5ru6juD1adOKOBTdVm/LKn
T6gMe5mYEfiku7whFq1wOxrknHc7kxrHO66o3MERheyeQbckLIdMMDjFF1VtQOs/QlpSymDPqgBe
CDxGWCVIMzScLZMb9AfcLfE7N/uCSrfYmrMqnXnbWVClOo5/EzfIj2eE/cKWcGpI21HWyBiCg2ar
mMNU3jzcLurYfFzQgUHGq15ES0aNwn0DJddFnptOcbBwFOQCYRxXIognqofeAFz9BsTLD9e7t6ub
8/fzKkiHkceWsX71pIfxDqtbQtxz1To4tsiKGcKENPFAjDYTQvuaZzUwI1J6MJVZTLNOo36k0Zml
hk2xhBDbuiMjzeDILoJZoiC8oz18lJrZL1amTu07d2mMEZIul7e8dnrc7CrWJhrIlB4PK6aYbNvM
w8/MDONa06IITVSwC9bZi4eBDfOKcVeHH4xvH5Rbaav3tn5OA90kd30yw2i79HgR3KyWBCpTqoWe
J9hmDrtM2bW7A1XFoW279+dsYADHf/QFurZHMKIQVuDNJOnYifaafgClE8uGCcEkR/+U9mMpBxeh
/rtmxqGVBLo2v5AimdS8m/iWsfalAAZeyv1jSs0f7G7RaSxmhG8H4ytUD8JzwJbTFGgUo6wCIH+T
9ZRangAi4RNpV+59Cyrj5fOwe5rf3lz7IBH7qDNQZomqr28/wD7/iXQ8ZMvw1HSJY5GerNWq408g
F9ZaIFJO7FC/4tkyP9HbVicSvf9l1Z0C+cjz2omiUInkk3v3rKED2fuZsqEfJ+6RMSDtyCnBvFia
EMlcNQTzsWdT4CPMZKPClRkkrVDhYAseNUgDtY+HXd+GgcRA8dSdKX6iCMtGxRpnDkE8VWah3faT
6NfAnz4rtRcQdzcOTNscI4+Z0eIw9hP2zT63MACDM2I5tQiY6ChchcH9cCKEbmUoK5ybW1luOOrL
ee/dcAmpawFY/3hq2VBFYDVsy1Ew4hLDZgb/ldwKuNiYdDZavz/MzyRYo4oGiC3pVO+MVYb7SISV
WmFjxCWmht5zJeNpGj7jQE8dIpM9lMCZmNRG8WciHHShLsBqBdRTzI/MPUyQon0FTTXwhXUh/faa
52U7/KVm41J8d2K+3qzlZ7zX3RL6Em5CESVrWxrJnHcHBJwJjKowfCKcXwANQKmHJ0NdIfW9w8V8
SVMB+sWFrwrymOn6gHhPIsZkjQ+hu2T7g6dFicBLv5JsmaFGPK3465HeNmHWeERKcOOfqKHIHeTj
XebjRtF9DCq8jiEHshQ7U90E8Qhp6A/frTisVCdmf3hi5EFojL2rRYirQYC/TaYnbECm2kVVYpCj
aZZKHTqEvPz7uJRXWlZXFkstJIpfCFDT9M/L/bOjabdKMN4wEseUeYV+8lkqNiXqsnAxpr2m5Dee
YlFfcP1iFHkU7vkzB1yl9dCSja6VL7csCZthQGItmRyDxHkb1fKkOCFGB1Uh/HUZZtjvlvmNCV/l
vvwIJ6ULyCFq/JX1q8W+jF1Iq6DXzkXMfEttozy0t/lcrER4PHtc+DS8W3Lg7aMb06S9okiW/Q+x
wJ+dySHwD/X68dmtBnPFca8Y5tqAstL5b5mjh9TCuXfPERQqVAaAL2uebVX8RiU3MYPSX9RGcSIg
i9NINx9SHt7FGcfJuVA/RVD/9Yvh1FFkVpNm9ePNVWIoDmrAYGV0tTLfmQ0XJJXVg0xpVkPD2IiT
g0ary9bZPFDqHC5u8p5/jHoJ84Ac/KtZMsH1X2TmmopFyXwSaVKBpsv14/60wIFNJhF89iCYz7+5
DJ3WdKH2GHiB2JJ/TQy1FH+DuDdxO63WTE4UzMzbEx43GIML3LB6wB26aVQCGa9ToZ5Cbywi+vPf
zho12yDkzg6cbz6WRSvXHRqsn6vrHo1eh9ssLA8Kppus0sWqGn/SvSjAprl/6GzBxI2IQHO5yzwD
mtuvqT6ZdqsnzpsXdT/o27WtfX/ao79/+4fKmc30dtCiuhPrnNnVi6xmJh7ONhgLiUvIRwDqoKpt
x/dvyX2jX7ZoT7MtblECiKjK9fZ5XbMVd4sNKDGZFX2dYA+JirwwhokO6Z0YW6td2RgUQy0kREYQ
74YR3lgkpLBvBTcMVdAzJTsJK0VpfxmoFbXMhEcOaORKBBSLAhNYH4M+Ullq9wY9LOE2hUowClMJ
PDhxLM9Q4M7FnJ+MLN0OluqyZUq3X4XioXy9yj1fk+aRbu/lK+WF2CIXur6uoDaceCBjBe+7AfSQ
CgOR+eZ3v6s8ezKFN6/69V9hI/23wydcTpE/b2kyrPx+pqRP/VAJBKRqHvmbDuTQ5BCQ/rG/q++j
GszGMaJdAx+/VjuSwfQ+bxCNXkhMVGTbNdbhKwn931UZF7xO/+75w3dLeMKTjUuSiWT6YWOaRfAH
U8eB17kSnCftTpBvdaQKV/4Y9GposfaZl6eTpBRXMqpyRHtffLRAcQrZMT06zu/38K2vtHfj01sj
d/8Ra1esCembVG/+mkjUk1yvK68yRxzXkwCBqoYA7X4L4FVqV10Ugm34En19zo+9k/W6XxGiCJWf
TqrMkX6OLtDEELkELlbX91VLgtNXr4vgvcybaXHO/ha+/a5XvWlAkz4qDa3PW3QXvt6KnsWY0fdG
NLm4r0iPmMyhw7axKItDr+qiGOPRo5c2nM936T2B6L0bVn4oS/iGoDq4ZHevlEc9IZ1cy1y8UXsb
aM79EgtfVIBE9KrfHOGhuseq+ObO9rBCrk7kjrgSQtCfFhHaOS0/dbypc9dP1GcWlX0MpRAW3qTk
dlb+piLzAtbUS7A0TCqb/hH6MgjTTGReTf2XMgNZlqlTPMmrZUSiYO3srrfr7JNLDnimpDmN1CWh
rMxVkPGeGKsJQWfIpWFhJQKme5ZoDBAe2UP+hX892Tt1g9z9h7riRIw1yV5mzD40t/xny6Uxy4bq
Id4UputxZvZ8ymY8zJvIlMejQIk1mtyy+c3SBYDQIX53srRauQERMAQNVEZnSdNHuRf9/UeXLLFy
ScOh7nH3YzQXc+6kofKZf29ctkxnaEO1m6yFaGAVTnJQvhLw+LbxjT73qgTFkQLfkShXFVO2POO3
gf0FYkdW6uCp839baVc394mTQti2pcQ9hj/CUCfmqwh4i02xFR7H82Dk1GMZ5Fy0rmNCBvViff/R
kxgKeiEq1QYjwImdEiyWVdnSTJ4ZGkL48bApT2XD0UVuOC9SQmXag8YPDVuGgqD6iM+7vOEncYKs
6t3a636gqG3RuuRxliygHLF8SyARL6xx4+wXcWqaFQyYCSJY7uVFie0BRieskkIbOjGkO8ZANACv
lwg3jSCcErt6wHc20mHEeAbaKyFrwRRXIrK8BcYWtC2CdLKDn28RtLmscw2jSisa0D4IW6ljmxfD
UUeQC9KfP6kJUoHDl7Y3nPScGzx4cQIgbggIjRrqR9IMQUon0s8SaE1JUHHaT8L+KZ6xqD/MTxX+
cpsnkxkSFmYfmNY8YUDB965JhMO0JAappQfqGa9ryiFLdsCBDb9qEnwWDW9/5mFnuGCt0biBNnz/
2lAtKT2kadOYwL1xOXdqNaA+5a0dxmXK8lKA8YVSRxwXZQKnVaWhbxKhk19uIfR3+4/5EodVIucc
44oSd0XDkFS4GKyK7x+22gmg15DZb8t7g4HALWcfq3FCOWVfwT0aB0ntDdoUdaRg8JJDeJGHcyOd
yAdrwENv285pF3v6Oo/CqVa9GigHigp/HO7JVgZitclykxiHNqKsqDqQ5alBwKySChSUhU71U0Tp
PomlxFx547fLLYO/yU++vzUUqFa9mmEU7uwir+1rsxZe2qa/MRZ8Wg5uzS7QcDQa3/G/OiMNe9fn
RXEfXFgINP4eJzQfSPY5oX9ccBGLDEu94n0eYHGLHw4rhe/ZMauNqO5aHkBdWBz+Uo9HxJTRWmPn
1jS+LvXFr0poGegIld+711TzwUmW67z2KAXIG5MsI/H1rPBFDA3Rwdw0VLOk3o2kRm609u4LCEE9
9nVDSyo3Lvz3G4+zuPUBMzcP+x1iqlM6+tHzuzNcaURUBPkWeP33Hw/U/2jUPg3+uUhMCCKbeO7B
+lgEOKKYNK3ZmoQgHf6JWg2oBWNe8+TLnvVmnzvi98JXNw6+N6uh0kdFeMb/xP/Otv8HTlYjN2sP
fxEV57Oy1iajq5qgV07cKRpLTNjll2Lg6j8LRwHXrAHkQuSudSkCbUioKim54f3n9XsZMMGk6e4h
TrESVXM0HpXm/NH9TFWaYMjXDJruAhnkLYbKMlk8JzQmHyVvdYktX90oGZFOEhOqT3WWMDUaZQmT
28sNQZBnK0FtgBuC7JFCiRJONNWB7Jt8K3xPeYeHYBfq+rog20TPFVxnuqj+dRX+j9n6GZ6tskBp
yS2npkjfeDBYv4uNxaA/ErfUiIrF6TfkSX20ZTH3VmfwK15idfN3bdM11C9N+Qu3PzN6nE70a8P9
VeSI0P/WfIcc5ueUE+MXhwxiVrZZZdMHLKNmYO5TIP29houCZkIAMnxZovUhLaHJMjHSjAFJ63J4
jpxbBJVNRrwoWHhEJDp+xQv1uD8YnXpHiU3/ztBM4emrxKjymgplPqU27wil0jeYMpUw33/1YAN+
P7PIRYYVjm0bqsgxFaspsUWlzAytfAUyctklsiS8WrISVQE7BtI4RWqtFKvEspOfaRoSNo5U6KaQ
Fn7gZzNeMLX6ggT5CSLkfc6pyfKKTfc4myN6WiYtY+bUa3IV/fF7ku5qtknUuke2+xTq3WqKcKtL
wF9C/075gCCX5e+bYtp8yavIoG+AzK/tIXn7ML30+qjQKhD4JReGqxefl6ljf9vRVpw/8rLxg6qh
EZTseG66fZsX23yKZYoBhMBSZzrOEKutQLnzT/doIDko6Mnp/qC8f5hRMkN1VzTE15QPvzkGnWJd
4ZOBb4t2dl905oRKne3KsxDrWNORc9TXk8kyPikS5WvlNlb9VC9D1BZ5bO1l2OkLnSmgKpX8MoPW
FmXj5ODwxbmvivvDiAsCvzS0xigXYt4Y/C6fINNpDHv+rzxaLVCMWTTAQkfEbhr4bLmW5F3wL03i
WIs46oQqRDqwNQGpjqze+xS/Uc5+D2tqZXeXRCM6L67ZUMIbgJLmhm/KAb8QFlu83aAs6ZJgLUZm
Uk8JhPbBxL6F0wzLYfP8WQeFZPUCH9krGVgFLRcTdxyMLYO3ybhmTLlrt5U5PZNPn7T70lswScs2
AcYtDOQ94u/tkRujshguw1J9zHx8tIL+kM+XP8TlOlxEBOmcIiGV8r80MShlhYM9yde05Uyjnbhx
1WGO1oLMwKObn+pGX18lfRannj+1vNUopOEyigYcCuU6Vfw8o2W+x/MHqSu54icVkGBMoCHOLypD
k2cWRdLsQJwnkgyuAYqaIB0linhl+7rmWBtGJOohgsj3JXkjUd9TM9v7jIrVc0BFSJTHAz2kiyt0
PSLl17Lr12I1olgv1x8tAOjGc7Z1m+IBkAy9CtqXAGGEFPhGojNzwVwQV9OYx9i22+0wbOXO1N5H
4jaWzKQSSdQpehJP7loyLugTXMGIj4f0kIkGPT36tFiWuCY9w9xtlmshql16CbBhGDN+lye7sfWa
0Nh2oOtcpuuEGM67jUN7o/bgQWSw9C46lUbOh2Pu8/WYoZxysI0yVmSbSAkuQnoXzLLp1T62IKDy
2iB2QVauofKQoIEHQgfLYrr44M/TJfnQgbgdCgs4190jfBKnqZ928Ss6/5JvWEZTlvbsqRmRg+sm
989h8ifrALHYml/xW85B5dNnpNDeM1Knv4M0+f+ZK74hO5AR/Jx+MEi3fTuJhhCcxrOp0GJdsyLr
CMEhHNEX7dKZT/7Oy1mGTZL5ilX/IT9q7VUX3JcoN8/NA8A9+sXxDIBm80X1k5/KqPjEfrfSq8Ao
MInVxCNj+rBR0xYQwW/0fJuaRlGiqWsXpBj0V78pyDfbLIsmSc4rkGwqOAPG+loIsD9wJ9H9q82t
UQHXGs+0KQNTQy6xPEfDWheNFmAyBVNi8KsZe7tMPkbZhR6ecDNXrcLN3pcT+hxVQWEAFBOn/sWF
D5XzY5oMJlytA1b9EQuiRmhqZzbBzsxDs5Dw2ZTMGvbnjVSi7TwgoXbTlN2B84OCH69Jga+H/9so
dkAaeJAONOVkFkFP8VZCYxgxJkzLxybWTImK7N+hcsf/cPW6BpXWxDDvMWu6jXzlv0cAd3Cyyc/n
DvYkfuXAxkHCiiA1RltB3eMxw+7s3uv9EIP8VY5afAcnOYyhFXdLP9v5bOi8ls0Ig4ZRk8bDgC0s
l8AtRrSzTK/oHe9VlX72eIdRA/WJo8fiCsjzKgJP0axPiq6MGLRMuc4h1w/tzItDqtFXgKE018SM
/LKlUroelZD8k3jVd4p8XXmCrIItJm6YwLEBtXaOHw4sJjbqMiSt6khVykXP3ZIAulfqZIUObsol
YRYnoHnzut9yT5m5y5AtAr1MVy7qx2CHnQDBZRCuJB6wBrSlsttZ1ACQikmVVUP1P03vw8sdRsjg
k+SbwBQRG4stM+qHVVFbeC3i/KXEnXRpBE5HjmkpRq/ca9+CtyJzR6dTTZUXfsqp0Bcbi7fq7Ga5
bMcg/6DjezFajWateoTYPI4G1Gu/91iaPhxHoEdgHj/QeA7NZa+mtANO0lrordCU4S5N0Q0Euazz
QkktI/CUJSE3Coxnv1rkjJk46NKorwWwwNaTeNzecWWD8ymV72aqH0fhTgGFA+kF7z2qw/yGLJaK
eEqyQiFlukNdi2KwBn4Ne4NON5gg+G239qCFQ5Aagu4hJ3VhY95nSyHIJROwgPIZy6NkdKgTXLOm
pIjauv6bsVi87R5sxVTLw1bMbGTkskRaClgHht8+XPg3V00b9wVyLbsT5p2rsjE9OqqxYdI4qaPt
y1lNCqYyNu4+hKl9vJ1FzPs8s1jcdWxRzVAZsxUypYgxoAfamaKpvpHEiqIHa/b/H5RZtNrq0s14
iEO+HujBJ6GUxygH4Z0M1z6z0eTgFiN/k/L32ot9DxEI/OQKESTq3v5qDffxa2YDqlnm+upvqdrH
eKywZbdyueBmgOSUCHcDL8wt0Mjb9HVS1HkSIIEFogqHxMnb246wAmKrd9mLZBXJA0rS2PZLeBc0
e0VNZNLinYawVxc9vlSHf/qaP9hCQ2fzO7pRZkLCX+Vq+rYGGEqm03DJEaN8aXlV0N35agVQYUBD
cHn6s1RKSARePGc1F58FfMpz8MOzortDwQ1VO1aTipZDFpVVbvGw+vvi9/Z/yXTDJoETqx6vNgo0
VV5v5N9ttlRyOgdleKcc/snqWx15TgFHD/WjiCPMxhMDx+IBrzQyu18lkybqvn0jP59ihV1AnRD7
XYkszbhXnpO3gG1O6ivTIbTa5A31cl3hMhmyckbmB9BvDL2Lw/xRP620L1g2w5J7/bi9F5ac+oqN
NEi+ML5/gUPIV10T7NCy9E60Lml4f75zWTEhwBNv1sixbxPpU0G3ixqw1VZF4vAtj/SnMBJrPnoS
BzrbYLkYQ1f+shRP8+TiPWHDUcDdLUsPmdoVG+G1oI1lVjKeZ9j/QB4D7Yh1gFgWW58ktu3VR/5d
fboghjHdTSECk9uFVlsR5PSh//9KjDyokV4Lj3ZGUXuJ1aGve6MWC0qCUXCSVMrfs3TA81yRy+Nt
3NVdHipaJdCG5bWXXqLB16oaD011+XuoWPvoGtuGLeyyA+iGJLxs4zZA6Pb/3Kqbe9i4jS5DszPh
++GXb5BB5Uv47sM6raoIcLpBCH/OAEbha1C3EiXW6lkUqJ7W18ae+sYpwRC4lnffY0E/4jSsdU+b
k58OUeNWCtOZes+D8t7e1PFd347w4lrAF9KxmRz1gLzmrFgYEeWN9pgb2H5qz3GD+rqgD1PE3Xfx
xTifpN9YCfYOQOESz6qAdfpzIfc6JSADNPWLKJVhQHUB+0K86gRydfAiD189pUvZQYJ/AvuYrq9Y
lFkuf/k4Iqyc20A51Ewb0UrhZn0E/vNlt59mAGD18O7U/4UgjYXRTZCFLkGZ4GEHJBZP74jYH0Rx
7Sn+GzuF8m3sZRkmIvXhI51YwkCTlEaOmnsJn62PwCyyF8BZQ/PdkTU2dsL5Tb6K88Bu3CADBdv/
gbwIp3m81Yt13Wg2QGLK5KpM3VrLuNlodBV//lf5grrQ3w7k/7Mw8xBX6dLow87/vdxHAGfzaa0h
x2V4eBnkLo4eV6eGJ7bUCAhI8i+WYVQpkoJrjplMRm43gyOUs97WG1dUrVcomxi1dS+OF4m0f9AM
6CdyevuCwAWIzeskiyN/WqC4+MgfgqEjYRmkFTdKl7eTm7vVZPWDfMPQN/POYXq/L3ZbKeiwh2Vj
F7K1sfifWt4BgHxEJBME4O1mSu3RiFNlHlCHCr9RQ+w6IX0q1KNBWzzpS/Migefg/fQ1IPvulmYB
VsgHB/pw2hBOsprL1Cwyx6HZAGQ7dZVuBxfjEBf7VigFdVOm9yVgIlPfqiW1+kYwbLzS2qTb97SC
HSMKCb6rTOOdq8OkIbpwg15pi1hhSFc0jy1ny/smRYb2RibG+hC87ilRxyS9yzw8//b8kRLJicHJ
Vsd6k78r2fAZ53GvbR3FRRZKwilc/s1xR7WskYpgBNwFcCXQ/PuqY2JzN1YxJ1SRluCu0keO5+eD
ZQwavZWmCEVPD+fSLaDSWuhbXpgb4wqGM1dwR7ZbOX8stgfYm6nmGOTL6smanwdFTqkQIalPMpHI
JBldq/GCBjlO9pkJuNisW0pF1osdRjcD5igtJfJ1dAjYSeaTtjkoKgCK2Gm6hR/BMmkR57VLDttu
83UDmsXCfO7UbR/iem5peID6rEMEbt03mCGbRU2cjTLXPsGNgVuFJ0R/drzdHN8egL8+6NqM2Enf
VJ3mFUWM+Fnm4fuXCewe3ECaVYDIjlLc7ea9nAWcNq9ienVITx2NJcDx/PrZJkvfbFYEOsvDyoUL
f5+zWOdnPQfO7snC9ybMFLsPUN08PqVmJQ3pR+9qqrj5AzgBwmzIXm34wu0Uf37rJ9OwNDSruw8z
2mP8yheO0SAVKZHEe383XJxaV28yw/9Ovwx6AhT3b2ktPFyrEmjvPw8qvQVD3y6YswN9auf2zehp
G4l6dmKmoPyJBcaM7SEBDODA4c4jvhu7fYcw/1vuxbkfZ+3s/ZvXeFDqa83iRSzQC1DpWQJl9fji
o1eyu2EFjgSXn6XPzmU35mGtQbAzMN4pWqxR+dNmnGOuz46uiIGrfBMMzcdCulXR5tNBs+eXdYPc
pn6PGKwXctSG/ZHiZ+JbMI87/6GWbBMuJw7uFvM0QrwtCsOY/fnqtcrb9pXK0EdVeU/XpeZ7DhvH
kObyHPwSPxxFCH8QtpaoNvZWMczOXN1NlTqTWd4LtaQ0OaH3Id2okOnJPtuLTppQfeHkVlKTY+Y9
Uwg5cYq+MAkH8qgFP72QUEVm/rcQZo9H/xOgtSnAVTbrMfy2HM6x42z5EZQj5S+6iTkTfxY0bbzk
neBR+PWbfSOr5qli+9hD3pT972psEc7tugrXJrcVb5BslpFtXqwbgJ4e+pvFqlOxe6DPuz+oysz1
maeYET7yXQKdL9zZWhNj/0761sw4/c/o8GeYlNwBL+N7nb/Z8xNw+gSNDCsqX0Y9eNjT4gUsSn41
3Y4X/ZpvxMrD4XkylcpCb8/prOrIiq/A62xutCbVLILUysdSM+TjIZgBF9kCKURs2rg8PGHfyQ9j
jJaY9MjFTmr1sSQBBbNV9M5fEPsmBMLyqPcGaFfqwW6lgypXqzSfjAsCmazGTZF1OJM8XgmawbHd
iIrDRbEuconz3SaEGv30++VaouHzhanr9EOtQCXU9wh6dpoI8D+TT49dxjrTgWKJZlPSJnI/ltF2
LnH7DBJC9eEW2F3tYEQ9Okxm1htVF2232KsnIvWM5BR/9W2MzXG2ZkpiQWmBagVCGsuq89Hs5Vl/
5Pfu2DlyeE2+wKUXQZOYWoGTdHpwj0gj//0nYcnQ9NVBC5FfK3pLKHfDjBcPE5I+NxwpzEWx4yf8
WVLpunkQydgOUtjva3KYvP0tWr2nKCwJ7R5sC9on2b4712gKp9RbOnxSmdwEr65IymIQYJ1D7E+9
THSbRPUZUiJ8xAezhB7E/PzAR3u6x6Djt9i/K4TBdqjlL2Xy1lteEy6yKMGr5CF0VRAxK2JKtpF4
n/XGZjEmOgXhmpy/1vS9W+UX23KJ+8mOY7/GaxjWymEJpvSRtllr9B+xmEPOe9HxR7mqSRAclhBc
6tuMsjUSMbqfPfMic83DtMfLQ4ibEesvS/SN0l2JPnf5tdBThGEc8+f0C0XU3o80fyHjVFd9UgBk
EWDGo26OP1MNg/F9qoJuUwhTlwi1J+9LO1Bpjs1UHmSSYFgYBTVrUh1+YjvFqM31ZvgyUl2tl/VN
6NNH4bd3aDw6CRSMT0peAe+Rxkn4j9w8/8hFmHXBHOEu7DURW27LDBuKs4e58rVmybfyI4I4HoZW
jlci8Lu2bKy7Bx+YMzKqRDZu91nFxPkBrL2tovjGpTVm+s5hnINxVHl+CIk0iVR4VKRqcrfSDhzo
Z5MQ4SKYZkZ/iFZB7mfqwaOxJbKmdiR90WZbCa8ZTWPBp1E3uHfbGIrfZ/DQ+ls6dSbS3XEzumY+
5sLRzqabXYfizDil4wnC4AaTYZTFe2ecmH/FfyE+UA0R4QxrnXXHEu+zODiCem5uytTMtHT2cfwt
kDZPuCungbK8uqxLhOiJrbUW1eowmCNQSfa/kIILRkSOVZjUUiI2fUr7ZRU+UHuCwKrOFWu3LkHI
Kh1VtJ8pZ+NZAGdnZaDglBz5hAhr4QbSIlLRB/AeK53Jt3kKdi/mfqykPa7X9ZOC9woWeTBT8VTT
3ElaYWMhty1Vj7Tg9RaQXepe5BzRBzQUmC52J4X0Ts+sHsLLnSqJxH0rDQ0OC6q86jaS8nrKtzza
TlEdCYAnSS+p/ufYkP/ziM3pM+1qtm+k9r3I6qTmI/QPGvycFpNbdsBjs/7FF0pzGHxBGrabD+W2
ZHUqMvlXcfw6LaFYSZ+98BXCx1/AnTzBuO/Qw+bxYAVlWM9wcYzy6fRGDTGeqhSXRqZRf8dAb5Z1
hc0ew7882Or/O5vuLOkwJCg+YB1TZbv/xSAvmvewAwr89haiKrqqIGJ1VGrSMBhKTU+E5LAtojfD
uk7qlJCFGVvaJbIiX87Gd6R+v+aDA7qnGA8uIlSbif3D46CHasHgaj0Q6o15ROwz+vWajo0aZlnr
2oSEVi46GukzYI04kOjV2XM3gOwNRXapF3R5dFIALLBn1ysz4ed2dl/LuP58Mistotue65Wv0f18
rVCqbTAYbekFEsMDmkm1+6Uwm2spPi4bhsw7vIIvlfT+Nio9r5nbG92vz5JsSXNtggZOJo5CyAYc
epVe6Xi9PpbOVPrcf/1zSlD1KnTIUlumriu2ajjzu0ZjJl3UZHwF1YTo0i6jElViz+Fqkl+0alTf
pLBrGxssg2pTPigOe5VvZdp7PJJjQgpeOYS5WaJt8T5lW6ZyvjhO3mRxFwOmi+PZTasqT8cK/loh
c4DTHFxbr7V9nTZwm9qfL9TjL1yJ9s5UgDXZUAzYuvmMyYU37zTy1/Ikkk5mH6N5Cfdoj9DGUW6R
fUJhpHy6WYLf3VEUG6SB5rqsY9OuXc0XS25Yiy0GKJOmQ7iRumA9nrGU/dxemiAJoIoJHUfXUhVW
22oGopaCuqMxe9X2JcpL82zABqH9xD4hfHJRpwRRCxVw4Qu+pz9Jx64fzfzkP+dbVREyGI0hFGVt
1JvjQIqec2KmWOj2I++/BGS/pJakByE4dcYqmPkWYMS0166NUuM46kEhMxYzz5SlrPqubzKja8Az
ypnXvqzvkA5dmx7b4E5AO5XfZ1TbuxNCkxL/Hb14NOF9yLyZIXwRwMaN15KmbTemAv2A89340Fqq
Qo9/bK5ISI4R4OC8IaVxWTGVSEG0tgloPffkZ9V8Im4fK1dfH89rZA9MTKAIMlDRT5T1hUUWcSib
7A5YSsHs38RHIrakw/Pgm0KjLpM+w3ZG21Zp3VRewxj6fqyq+GKUDpqqST9gyQi9tA3Fb8q8GQci
8veb+VCOKE/Ac/uKgvfBWBDVAvkG7u88rZ9SPWQ43ovE/YAyqAEjXiUOADWQSe2SqlbTMPabG+xf
q7YPCr4EvJ8Lde6HZRlU8IHr1TZaQ1wq8l0+5GA7Xj+yXm3Om0NE/d6fsIzLbJPd38oDRzURHJUX
DXS6LXEV6/PTM3doUGh8lbBYlR+Q4uiaMUNY7TdG87pgbulwsE7Gs4i+G1EpkPBa3sLoLDDT0630
nvd/DHngJbtVpCpo+YWEUbSB/RAKArsFLK61O88mOEJwPIgwxsS+eURmalWvy8rWf5nqkm2zr0pv
3RUTfyGSEYFcDaJCA6b9V3YsYBoOKRcsEZNQpyn1+BKAl8lN3bk41UQiN62NWDhAMMjdma08/gwK
jWbMeOzeowsQ6EmBwpK8rE4bbCMajYfAnJrx/8SJVnhtJTuhLQsq7+UvVGBkFz3x2nVFSGWZK6kN
s0ADD1uw3Gw2bnJXDGOaX9XOhhgWZLVye/wxHyPtfEcznJo19vSCN6nJKXmvJYQUnNcQmE2+SStk
R9kskwD+8TIv38k2kQGMWw93C+z8CFIwA3Cf9gLSksAVuD60v+2WD6YENDVTBaLVicl3OKAoTU1c
vzXWxsCufpD7NRfjlhtxEpGgvK18gddJUlGCZxPY50TDKvUFQFdKgcsAjll4Rx7CsDb2DujLJaI2
2Tx4SOzFGBFv/rWR/K/+0tyXis5Gdc17CT+T+AbXb41Ym9n5xkuT6OciGcoVxEqoi6isddjyDwbg
SmBtkIopqcf8wVvsywwvDFTl58DwUew7l/yE/++2vrPBVOs2VBGu90iD/coQiDKpcMFZkzLJqEYt
aU1orVQcmV2b0c0F7CWUv5t/UtpyTuqK0dK1tftn7AzuDONJeR3eFLDEEVuhJYItxZxhZZFtSS6N
A2gv3crnlPLMwtZkSa8v25dIdy/kwQklzubAxPsrHWishv1x0X/YTVsbvdmHXuVfDeI/yVfKZYd4
VpgBP1dM2Q8NFURCqX3Q7l5gvYGGVqu+MYyBry8OUYKNHYbB6FmYZCeFmyIOkmee7cbCzIf65Uwt
EafGufqDiUddaq5SPUILX+B9FW3+DnfE65ID5jdGiHINKy+K2/aBsx3kXgRapWrPZU48YU7agh1y
JSsNHudVU1zYo6+ktBl0K+EW1X4cprU6tIK+uEJNA09LYtlHJ+h1Mu3VEdnjS5GMD3UO5FjoxDLg
g9SEGW2Iaryth772wqUMStuHWeMwXmDMNIt2RS0B9ccdk2hGZVKMrz/Z1mqZkcQiQfhUF6zYRpT2
fhNh3gT1C2coiPGsU3dmwpsSoEP+0nM0NylfiWUgIJApO9J6Lrp6fvXJYsMNLHduBqTlmH9ePjsp
bDJMQk5v9KyKZtZawqPCIpAT3QevztHkS9ImGyYbM7Diiu8xknFhYVokSuBxMw0dj/eN4Yrmy2C2
rujS53R0aCzgTWsd3983DfIUjEGmVX9VKn/gwTOTEoATR7TXpcdopsZS6gwn/csTJkLCv4K59Dzz
Kis2p2RQFjsCFyGQRYirsRDwBzzJUODWheDmdTQaM+9Ow96MiA11KOvgNu8gIYlhGj1ORA8HvTZk
q0aHrmWdFG4YzTyy+QQKXFTrJoKXvb9R6H8/p3FYox4wAUiq6vNy7ac8j1rmtRSrxWJx8rRZbhsN
/aWf29uhuMIIfrvEEYDL7JT/dSLECJ4OEaCtd9AOZl+7b7l9Bf0oXF+rnIq62Lb1NL3/1dKJaG+q
L6DTZPOYSj55/JUW+bDjELOpfm4KztXb99SHkk64l9wmNwAljoeUqwsAH7UBJL4sesX9LfgNaIxD
5nXGk2t2854E89bYJVJCI60MyRvnsJna5bYSmDCQ62nut4lgA0m/PDpv7XAUj3iyQQyOTYxdKCib
1Nosy40RiF7t8d2ImO0QZJtzJZ854q1+ZOO4sNqGdbpLEszNP82FjQr/DUO4b+2IDWtkqOBzXCqY
0CHEaGxzZ78AoyXgOg0lbZ0euJmaMlpmxONMtVB7/PUrLrWeVKVWdi/VvQzOux653/Y5Ss9YEc4I
qJ1AJxnWQuTx2TLlINNEqyy63wvRuk4vgMnXOJKDYpq//ArQCFU4XVzW6rH/7TuFizI0z3e/715J
fmi8FJbeb5qgwTbE461gLEV0r3XgRW9lKKRbvInB1brN1mf0QNxf+Ed85UmH11oFThBsjRGSkORd
n/naXRZn1X3iMSBzw8hPt9gh9ziF5gqYn6+v7k8E01XIraotvK8U8udK9LhH7IrvKwArCw92+r0+
7UpY+np/oe+aYYOUD2ykL8py3gJw1UCCsIc6vbpiBNo7ygOGhwt4QkH6VygPH5h/q7TJ1nGVGN3R
Gx6RtdZaSdOryU2uAoz2x3jCIsXHwRdwxVKq2Ddy0dWZl0ZWyROcsKNb/XsenF9bCE30zSEvC0p5
eE9X9mAcUhgUym5uu2MqDFRzIchWpjr2NA6vQOh7+Ajp8AE3dqQo9bjJ1eB+ib/5p5rtMTyWSxZ1
LFYdhqyeB5tU1PgY8FfFNz0O36iWpz7nOffCMy5mjzlZk5jDHxzs0oQXbFYiAmPYQdL4cBw3ptlx
zKlZnKHKwkphNCvM4oFQAquFpMTpcpGB0Bad3NDkxIdTd+baMs91mxAUI0c8NMSmw82grbpcXsrn
3aGKWA8GoE3MBqs3clqENn6cY3SxJuHNybyLcNypeNw8WcetEuzvI5Ew7ka135aKqNN59rUgQao+
Ewa3CKJUZWW4Ld+VuMIiKhHq/DzjcyFHfHKb/kuD5N1tvxfivu7smfrBp6F7hpdW9Bhfe8kgIGTk
4xwLYxtP46Q5qJQB4zR4cVblivj5Qalqk+aV8S16hOMpkEWLkspyJwny4ZFOMnP7fF0hw2adkH59
VattTQcKUxnS40hbPOVSmJPqHi1s38e20yXlJJvOYl7eZ1b5quBhcknpK/WD8qxOAtdvJvCzAGfQ
raSDZ4c7otJQ7m6WusCzk567OCeXUAxgkUElCe/lQHVw5/9fN2h8MPIGbbQCTeAeIRFXHyKGy0MY
AYNLKIGjIukVv3wGUgu0ey/wkW4DEdMy5U0G0j3uMZeDkRBJPA4tYjG9z2G3bGmaLRoo3JFJDQ89
hg5hsEMcQJ/9cYEInGNYQUGBgK5W2pfUGXNexfM49eRnWGUWW2fLSi/Igrsun3ya5p26NRy4oUxy
t+M8hs/QJ3sg6mEZF3BM7OQcI+8WeaC4qZEUnsw+GVcVNW9qHO78pn1bwPOpP2hTrc/tWP8+i9vM
IJCQOz9+j7q6uNcbuzfszl/ga0Q9l4tLn5/H7sSurlPJx9oXNlci5kvl3kN7+vvRe/B+G4iyBKHN
7On8IZPPMBbf/asbzlU/6KM2wUNCdtjiUHgsgZV9+e1FPiq2Wt07Lirnd852p98H3tJoNgu0XB/n
4ewO1x2VD/wvBYUhv5vOOIH/HEZFAVtmT5T3dHyX2mKmOdxB9gqRhWqBUsYqgs9BfDenkqzgLXJ2
qfeicx3UWxUtWiOJQrzG7yVfLtqPN6t913Wip24Mj1dz7Gr4nnVlHS+QBBBIQ62ryVPa1FxpzQpz
CjH9OCYyqOObUcqp2C9wgk7IZi4OfyfjiHXKxZYbm9UIpmSQ/b7rNG8yzI9y5Cn3KRWzYvOYoA7A
0DYEk6AsCrc6oDf2SAYgvyV7rcL60jIXX6BrTkHSDUUknwbCcHc4e3W76A7fr/eS6E2dQNYlhnCX
nlvUQBcGaslhCG26mxG63EZaaY+xTYDSp14I/J1pb+P4xdLpUUQzaMTNeKJZkTyzWxOj6IHlswBV
8e9sRies12iaZzgvGG+6bV7Ca8DfPGLKPeY9lAivRrmQ61IDs0csMStnfFFpdng+Rdf+w9C2MjOh
zwbfKWhBJq4SiiTPTlSvJPZsKkG/QAB+0fGa3w2Yw9X3GvLFfss5BXxN1XfoajySVfviZoEbmI9H
bBOtU4KmfQeOSlfDUrvTiTZL6RR7lHVpoOVhbTWdIj7r5iwucAb+UZoH9DNYVW11cTYDxHv8kyMI
LK3JF7bu7DBPhEgeY1itysItogyjMfslbGaRSrZz7SwWmz8uUodLWREMoBqRxoEY9VVVDObrc0bH
hu04z5hyZRkkNQ63/l2muvPqbHewgpK56PY51lhfHCOFHySQ91CWcbKOGDCkeDeE6N5m6wXaM4ML
NvAibxPLxBgnCeYJV1oArUpH9CtzUrYNPwH6s2jZUVUv9vGlcnptrTT064etsw7qzZncbBwwER6I
i+CqR9rHEzzQDjSSoM9unkKavSxZwnWdT6BDJ+PRvu7sEMWhd/1B6F57WXPnMRyD/iad9Fql9rlg
LLLDofhKRPWok0KC+V4NUlajNQmD3cKb3M1+QniiRN0zYMd1FE1SUNPKYZh+XI8O+5RpOtqzekry
L1dAao/WmE3Fx4pkZ1GsAwAyrOmaQ/yr1maKKtkESi+fvr6a4QP1ggN0jmNzFGv1fyp9uPOBXNKp
SP1jhJsRcpvjitzdIVDKiYXrJmWmv+qb4qXL1Kra56WAuCWZkItE/5x11sqWxUPKu6a6/7/msZ9V
lNQlORaF0gAI6mBVyL1+15maqhWYKFce3V/WjoIigGu7tYiawoX5MkDd/Svkn3i5Za2V0N7bRdTI
Qo2XPLsBK5oZFPVOK17PHo9Qt5IDsJxdywLq7dxsUi4/myRuBmgR9evp1mwht3aBht/IYJYPYQDE
+wQCyHthzWwtBOGxXv0mHrn1ycmiKXX4ZJh0b/vqek8J1VlW/Fu1X7oNdKPzpRNevGrhsfqr9f1d
Kd/JnbggQWL4qLrjmqUrVofm/UIPoXgFQvyYP4m/8ea+Q5jeUnNJieJaDAYMkjFPv7govQh+xZPr
1x9UfWGV4zBL8COX6Zp1xCdtfOyRp6EX5v29Wk3T+zJ4sE3A4KiuJaL0hHiJ9LV1q0h7KW8P+Cxw
iBQa07yCUnqEEADsg+NkDmdPA5H9czoa6Ceob6h89zU44LNqqnhasM29SeN5vjgTE8yF+8VZw+aW
9Niwun1UVCMBbepMVfyUhApakgh4o6xmTQLoypV1EFzLONVICjCUKfjG1VI912G1EMo9V4sXrw+p
4V7O8vBwlMBZfsv8woE3n5Q9qvhID7gufp4KEOulC7ReUCVh1Ga6Zw8ceX2RoYLRWZ0yxNugTjYD
KAswS8/UjfYYp904YH3V5srRPnIy89iEE1XpjfjDbl52Ek4eRjOuacN/rNjcKwk8J0aVBlWMQnzN
8Xbj2sdfSy0zWa8UANzl3J1gfciZwMb1KGDx5Vv8Sl8Xi7OFBsGwGQrvrxHoyRVBCvASdGLvkl7k
/EsLznwt0poDdV/H+VpO7KQmX4tQdMcfle6shdPCfrZSk+Q77NAUXjJCKoK1JNdST7gh6G7SehcB
OoDGGB/Z+BepY+i4tWXQhGZFKIUujYOtU6BWc2Ud4AvEdwrC/n8JRZFgkUZmipxYq7qrAlhcHzMN
1jt0u7T0f73J+a/3mlvmwQ95DSclKF9t+Vo0TwOBbcHprigPiQPHc3acKLG6X57ao4G0Jmt5iqRP
G3IqAr8RHhf07a+N3AZ0Fk70+TVA6uBwzx33x2atxYOp8Cn/ch+Ts3UoMn4aWTh7/NrzPLnScS4k
Kw6aXNCD3VLwwKEelAFIvepdWbGPG1ofqqxlixjkLD99JCUFkez0PQE9KjF1zu1K1k8WT57bPHxK
J7XJ6xtNMM1zeZc92fKGm6n/KSlfRQlOXUPIMwj8LX+zgekQ8FJ6LQm3S7GJf2ivdWJMN84rK04p
0fT9cEbuKW2lcN/VIODvomMOVzIUOaZl4NVDqG73Zs3LRx8OAkKpcCx7RXTOam1PWTxEAUp0GurC
V8xJF7/XNReBZwnKm0pRskLd02ksHogPspbxVP/u3xi0bcYsKYyx5iLOVcpQuar1g+bwXrn+8CGz
paUqvCsXhsYl/GFWayYPDFPqMzH1RQUT+d21MWN8zgXCG66/gMl/j0v2uw8fJTUuTpWDL5/HLo44
mHY0fZltJyRvfcaogGB7U80TUH3YRXuIiP4ScWrDzPNjAZsfbPQiEGkvD7tozrvTjuq1ETVNRWrK
DqeVj7NQIW62KnkJaSHiTOvZnUjWhZyg8itzfFYlGbr3SAmSBKQsNqEi97xGeInLNbjoyDwzDolP
d5oPudziuTFGAhnXGD7AQjofimKT/fvGYdc4lKMD6+VgZ+LwDDTCmnZ7eVhg3bwvq7zCVluL9LPu
5daOWKb7wQN0udbrq32KkPccKkeZDM2vsn7NxAxaPQoC6Nx8yiXeNm7VQq4bqd9T1QBF/2GJNwaB
CHC5ldMlgkedZgI7DEvA1NJwga+DEsjpqUw6Z12GXXFbZ/4aFh0r41sqUiuMqJOLRAM4JrBPkvG8
ojiCE6FJwaP1Q3M/1dIPfJ+SUV184zvckvZspOv7Q+kI7RVSXVWMRgF539aJWjuVbcJGBpIZWwFw
YscUobGjLbCB7vFhqT/On/DzOeAnXGpBzkkjj3llCMRgUmeOIlAnRAL3UCr/TIMbDPKZ2cPLqogR
UPs9hH81VlsZHG5dLuTzhDCh7N3tQlVoJgj9+efXIzx9zeS+krBs+G+GchgtRiup+B94VO3Gyz44
iPzQW05CIl2CEk13qz7WmZpU56UoDGKIYflvdjysLy7JcKDk2aNYikGqNZxKlXPXWE3c7orvEl9h
cVmODpxarh8LqxOUZjYz+lzOr6OglXKMjigMEH9XGiGHd4gXDe5gtZlO65LtB8jxp7HDB/MXeUPf
3Axy26EJhXQPM/AzDFNldIC7mehvZZbu2yNlwEQVXv3MzBK+gL8yIXZN5I6lqxju3RkNEM9gV0Fi
VXecmcn8tmpooJdh6RpqKDbX2imCt0p+NfEo63/TGt+t6h01iD9CyQGMBZoMxtxjvRlkgsnNlbli
P3mVoFOk3TVYLlx2zU6Sxskxy+vfbcUHp9XGIv/FDqCmKNcCbKzKY7Dd/fAeenkyk2tvmfdqzkoy
1HS0oN6WuqKQaja8GqeryRYREG4RKJI2Pyn45OnnunViH406erCGcaVz+D9NtthYGKDbo947sJ15
45X8RY0W143PoY5wrLWHa9T/yYikFycKABsfEH6BIzylNkrA48BJTkSP97c1yPqdcRO2hJwIPkI6
WvzV9T4qfFRwWFcP1gOJJ0NISx18pjsus1EVKIZJKI48OEjTzZClXiX+jBnydAJd53Tp4oLJq+vu
KXbitIE21L/srdNZLUL10+cqIKkh1IjDotUwYfBK5Qef97RtYlvVlEgUE4AfBHhYv4HF2D9qN3ga
SlJRunKPU6kLrqG/YT4aqsLovDlgpshtqcWAOmebEcLjWnW8Bu1oIK4EDN4xMfB5m3H65it8lfmy
IP1DHxjj0nxdLhewlX1Nscj8RRPmsqin7K2lzAy9nfuYKtfCR6nAiZZ+9y4MSk+oOq9zHw7KhyaP
hI9Bqn8lhFQg/pQlrXx4/guAat9QiVQcGDxVWUUot3FOkWz0fSbewfDFNMizOra4ZqDmE5lmzXac
nUfGTmHdJIBq7srnccKh+NXonCOhszSnmt6421sqx8XnZ+ooeSI//ln0Odx+ZaYZGfwtOIRa0BfI
itHBM16lXDSDqkyTtSUFPUast6fAauMHfeg98OJGIYqSyZLlKbuVdWg4WAQeEGCRNkXXRR1LNLC1
zoXQgmsHhyx/94ZOBvxGJy7GOOf2T83d7RQyQxQErj3f6gVIffMzBigzRh+HYwwtTp6Af1bvYSjd
bOe1T97a4x28728FGvkOybp5gT3LcJGhiaksg571gpgg81AuFbWC6Qg6PMRBDxNMZ01aU86TF56b
KT77hrslx9vihWLKtaw9MhEkZCNSmvw1MiO+dh78yDrXAYxqyLSAI0kx3LTq5R5m4BsthGE8T7JW
E/1RSf7uUE/cQgiIvv8ZGfOEbKc3uQACVv2LMXv864ScHScasBT5JU7lJCkDX9KCFpKSvjMtQC0H
sucXv1CWsSCH4Pr7iGHwGkhhgNX5oqe6RyGPkqK2Q5HrpZc7yVSLBEOYLndpBwiRBb2Lu8OleWmj
SP4Pp9XtcrgaU6afTlHioq4stOSAx0xoWoXRFETGc1ahkHV0R3QXtY9OrPwZEDUUWOHbIzo35pAl
pqBu/xWqj+TSdKgd9U+mk+5Beq632KpSl/ZjItqFGmang6R18J+ztIYIeL0pcOQW3prBOOZ8VG08
4yea3Qohieto2gh9qSumaKo/VInYJiQcxSyMGbJ8lQV8KxnXCPmVHKblvLR4EytFn/0TdkN0VLoo
gGSmFkrt7iP2Aqb4ZxnA7UIByVii21Ib5zt6GGVl2us9LgBQlSGAXfk+SKiD2UIx88uvj9mOgnuy
U8ZBxXohsLvjxkm2McmqULGLKw80ICCFxko8diI/gzjyB4GDMP9ABgDyd4t8t8I35/KM/7opmDth
w4j9ATp9znor4vuiSgfyCAR+XLSO9d3Pmw7fY8uUthwv1JD61NLr8bpR9QeC4g6mxCIaOJipzVV4
UCSEAf+8j216xrFM63i6rUygfwuYQRGcp6MAol/gxRAId2sm/wVD/NGFhhz8fhF4IaUYfEi0dN1Y
ry8QEk2OZqxJYWXdrnHzLJ8ZL5Fb+KEhEpGRmnFw25kJsIkYWJ9jmKwf+KLcqREmC86pe3RAYYxN
+JDnBG5bI8coPlskZ7r9s/vVc4P+xFbMYUmZlfZmsEKyiDHPafka7y3BNdeQxlhxFqDh0Kg4ZU9K
SWmRaTPmA03BzxhO9yXQPcKKig7tkDujwFtVOti94qaf/PZdQMWnReqLSjGEGm7qTd+Kh37bIFZ4
+xUL4GJm7AdhL/Kyh/uPUTD4fq1NYX6pP/GFc9Etp6KLswSXSQkFMkp6riPg2cRxEYergaNOGBhc
wnRU32WQknDcsv9KRA2gS/zGMY96whMrivh2Pijtbn5yJMp2TNg22Y1K276gZMKRmLey+fnSmKOU
4fjtzwfwmdqd41zwUIGh/e8vwBTxcuB/TS8sAudhvT+twDoF2nhj+odOjYcb5ALMwGXx6aqIDrI+
SY3d5SWbkMqgZ1FXTnpsZmcc+fUwLB62uU+iPXtyV99gMtp7wbECCv+xXlcUNKQcTUloVsEk3Yag
oewC+X5QOT6Xjs3rkSpko4SYPMsCYRyrFgCAWaA6srM/mTw7gnRdcRmF2Wj7c1xbkwNGBv+87h51
tRUht93H3akYEylCgJPPH/xW+ZQpzVoJWNHtKFKi0ei2E4qOhvSgKEpWNOop1UZFhZgO0zaHxCx2
sYwMY0SPDy7FkLui2fkxPu70f+K+lmPUShkGbjQxcfg/R/qER9KIrpC0OCv459nSy6oqdpMIauzA
asuqYAaRDTMkH5u45KxnhvH7aSEAFwazKW7mFmmbQ+38wjluNGPTF1Arj2CNxQAG0VdRbr/PFsJi
v7Q8yQXO9ML9arSD6fsnIFRo+8pDKAtiw2e8F4MkRM7GEK0EBUAyUcE7yD0pJtKSaI0ojpKxVQAc
KeBKY9gD9biO2ElbKunhTvlgtiWXBkKbs+ZvgA9D/F/ua2/VD0jGVMYCZ9k4meSyVm2uDa/kVHWv
599Sla4+u5538F1O7WS/oDhY63rPlsWakOhoVz3p1wZULloU5LPfXECLyHmSNheJWeHG4SM9LT2a
YF4YOSJN0hptIo4bBkzqkdUv22w2IgvwnO0krVou4N7ijs6mU0lV3xFXnw6OXYBhDR5bjQjtBrKU
qBlMFoXfBTkvaZ/Hgbd1iDvWDMzmuVhEhNqoKsujSN70Id9OV4U31uZgb04QSILIS5pKbdHN6OrY
vJpBU4UmmaKvdSvRweJ4t3szw1nDHoe7fCpcoE1U+QkUTM54vVcJz4eyezHwBaqU43kIBv3p6Gvj
BGwc84dz5tzVSxWYWNK23X+CR1OPpC5jzUbogOpu5RDg9thfzWYv9ES4+gs2tAjB0K7GNWeunVFD
TQhJkbq+wcWWl5OWZ9ac/p8hIx4s+h6iHg4zAX2iCDMaQk7o82BqBxdkp6QHxPY9dRoKsC33ubl4
xC/pGPoh5Fa+IUSIm0TffV/kVaTPQtZADC4HNXiCvjh7FfbYUUCLlBv8XKp8GTXL4Pnt3r42VL7W
yOgaBDhPdk7D2TZJSlnk9MLASz4rmn1KEmXxwBXI2/Di/wnvIbpU+qvm55vCKKSCrjlA1Kj17Wk0
hkRQWfq0aym8vE2QJHk6T/hUOfvG60gZiLV2zTAW624dSDdjbvLtwMdqVw1EiK7tZC66imgB+4aB
6Qm3JZseFQZu7qkiyi7vHxVkTk91DLSKIHzM4HWNVGPfTPz1h3N2OkoVkwWKf5NxAr8O1CdKSCAv
+7z71V5HCUdJWstu9xcj5vRiWVbg36RzRK2McK/3jWAaxKwtaXRQgYCzi8zXHeT3raYR0PWeYPfD
XSDBZL2xXzWBihlPEpWZJALPA/Gi6q5vZJ8dVcDAgIClxR7D72/34FxdUKEHI0r9fL0EZ3Q1ee/R
nkSBZfcwBIiXobIZRQyjz1VZoY9iaHPQbeZ3JCm8E3BkNxqkMWXy8EXC0bwtnVuGuz0qlCtlqSSQ
qQKmUirXuET1YrX8D3+2LUe+I84amc6Evn+qZO3XcIuiM+9BVdsMQ0Dk+6+A44r0Gu0E81+cqQWV
lFf/kLmrJblvZ+ywOZm6kqZRXP2zxisj4qsPMhYn3BYyrBv9ksGXfPe/GstDEl9gXCQy7O7BuJpV
hf7vDV5JNbL6+kKfyCUs69DD4DqB/r477sHzZUW6ULLIlFkHiNVZV5j2D4riK1o5Fum/f9fpEuz9
7SQfbpm2+owfLfWY7nnufdDhn4RF1a1y4IoZb8d0Lo4JzwD7cNo/8iC7m/JwmfsINhXnloX2zNbZ
BtO67NBVq2f0PshWSBBDblHfXjUEpU32flvgUKOUga5xD2lH5AEoEEggNdFqNZPhGuGSNPcnH6uB
YqE39xIQUDJkuoIYx3Xy4/8QRguR3M9sAKjzJZFTQlfUuKBMKCOSx5T3Z1i92doQpADgEGvh6QRr
nrQ1vHJF8nMtFCNxUHEMZJ7x4hj5ZDb/Dl9IiygTP9TnUWZHgB+Qg0gFqRjC309liBk7kD7MB6x9
gIMwSQ25r6rTOvLS+m1selOCGYc6KWDRHGdlU0cUGEUyJfTbDqlpS9JusEOQPPa6c5h6MBKdIZxT
VA2WrIL7tTG4+Pbrloj3rryYl/f6L8ln0RIAMSOWky9locKdamsr7cOSLsldQ72ZRzgOhVPAalp6
72f9Cqu+HGbsDYxBC9p+HpL+GGlcbHbEV2mxjMXmTKPXDfN9Uyf8JegqER04/1zQGOclzmDrNnTt
Dd7Nwm932WwNTEHa+pRrm/Pk93hUMJ7KC3N8+5nX0ZkASpXo7Zf9SMAiCFZpMMf0dQbZUC09bhh8
Q5lnaChRRdtHrHONmzXWUR7NggpUHv43swUuFFB13uA8nbMW5wnFtjfkxQ5I7lRtvhVq2J47Yvz2
6lfp0uiqGXmk4Y/sFaoadJebXmBTDFZpAEzoFhucZs7SRL10odp5FRXHJtuvKCXsRxJzrdzCkXek
kEJ8Sc0EKQJK84sxGA7i0GLj8ZhUMPMzd48/v+0ZpkWIvMN3LGWuvtxRJz9sWFFIc1GeSgBLNWPy
syZp+Z8qoRy6tpOkyrr5v1zeuJeVG0dsCTUPtDuB6oUqpXhGNgW23PXVRk9A0SiqpWv1Up9dWHUm
Cwpljz4lFAotJgN6ZS0/WdajLTnZfsQBFtshC3J0ygUAZzWhwf5//WIhgQGguz9nVMT1/kRxekA8
AkfEC947LIQ8fO28KCprBA8UvesNq8Scs9WRK1LmQSzm9mxP8rrC5pbqFubiB8/1Rdeug8FJwafl
UO9TEYgQHtJTp+014RU3FL2OVYz9hwiao7orkveUeGLHx08MmJXImL4Zu+d19XTp927iABS3TL0d
BohelWdS1L5Z5xraP9t53IwgTJsvGJInXspPM8Nv65+ICzluhPX2PJCqC3ChnMhhVyJp1JJZYHvy
4VXZf9972D+tdNSqxCazF15NJop2oY4OIa6teS9+MwkM+oF3LLbdCiaud4eFwbwht/kAr+0ULaIS
7QXXLWi/oPwCAakG3HWISyXY7dRdHXOLBXU2P4+giG/l+RFhL8k2Oh0Yy8FzJfRq1Xs/g3vC0GUc
V5u9Wux7FVSJtuBuu7lKpEprWw/IDfMw4V7y69MWhag6Vf9pngpeGhFnR9CyintAGlCBhHTsyIvB
aIOfdFYefwuj3EE6KDK0JWQSaJVuhohEJMIGs5H6yszZ6IHs37UJI4lo4gTdUocpix4b9O7/Yn9W
/GXmUOoKq54wOlzD145kEKE8gVcZ1t2Jnr/RosR09VfqYsfsgq5XrL/qRMDuNQQnq8XqI0MdRUXo
skg6dqdvAbHzAKC9aAgxHuHCRXYv1BxAGqHyulfpVLZTYyjiXpE1NaYKKJ31Q8HM582Av2H2KAon
RNNLn4vL0+u6sSELf8bOTf7Smnxoo06KigZyXhZbxRMHVebDmKCxKfFfhYjeMFcteUxuMJYmzt4Q
WjqZV5s9wR7myU+0E20Ma2RfJc1GwSkFXzN7m+LMhA1/T671euZOaupOj7WCyXqPtieU3+Dpjq5p
P6L/wNbPXB5YhTVuR4PqpF6wsFq0CT1ejP/N2J5jhJHX43uEYZiRb1F4qJzkDX2BiBgHCkRHaCpF
8G4EDOFvBZCO4K+t5NOKONOz6m0Fm/siodrEfGqRu9rNUJbKetY5NsoO87+LwZ56fVDrC+PBSdxb
0fc0WUkQApnAsSlSVTCViVCvTmoxkj1E56ahpgUvHEQKRUruHKEaCA4cyXytVu+Blw2liyDVGXPO
pZjU5apRnkVhocRNoGut8sflcinR1GGC/fxuZ4X1V4KSASoPIAyUekNc0GpBC8HDElQC8SXShfgF
87pH7m0uLhFMuvwMchqoIFTHOG4uSI96fm1e8f2IZ6sb7uxBCUVyDDCklCCQ9FqnN0WTDprFSTU4
8SmuuHv9VwgPmuhB0BxKuDVmsHCpgnzjwOkN5YMF6ZyH0awxGpXu+EMF4JBIq59+nWMR2LqY5Fw+
is13b1+emEV1QoM6vi426FkzrusHYI8sTlhck7doGb14QtwMcuX0QUQz+DkTkgjuk080L7JGroVQ
VKMancxfEGG4BIIY8P8V54LRU6Mma1y2hzkgU856UTyKt1err3WSVjvljCKcidCit5J+vimNPaaB
s6OWQIQ8qVPXNIFDOdfY3iH20nznR5OSBxFzJj3ORlUBaPiU+6hSeOd+p8XZxkG0FM6vHkF+R6Gg
GlEYBCO4N7qSweNHwMI50NaOdn62OvYSQMTljanINDcWFNEiu62eqiN/g9nnRbf8sQexBdBI6AU1
920w+yq+GPF7w+G9xAx7XpXC5Cb3W+zn71n07T9UF1APxpUBkg1fHVI4kUsEhtfRg+/nm1A8TgEz
dJsLFxJ0jRHdB0XlBW+1gVWs7GnUlu7ytjTybk25JpIk883OAt1jDJfEFmQxhv9hE9q4vBt2YiYq
82DBL+TskC0W7oNTTK6grMUu3+qKs1WoDkpOXCS0P6aC1cxx0Wnp5QlzdGIMV787XW7W+5LlVRV/
zM5ULafY8KDfiC8PWIe42BU2H/iYsG+rr95vYRsg4GtwjZwUuO7m4b1c+xdgkliByWJfg+Mda7k5
JpF/K0CERS/TmcVafTwxBJpLHuz/1YzpzP05byb3yeffr/mPCzahq9qnoY9arZ5qu0AeQF8Vs7xY
LcG9equ5BE3Nrkd6OSiBvNDK9v8z919ATCxaxKg0PONKPlVNa+4+b5pA8JZXvEq2SO1LcqhotkpO
T/57XgOUYFHVU98W6XZOSBHFh/+Ps49CQs3U51ltnRC8Cl/qbyKRZ0KEQAueCChsNlTGAN8hVv8m
zibyRt3WPBBc3FkMeTocYY09Ua5QH93kobbmX/+r45iZcoOVG4Pc2hw28vYjkY9+Kn+0IYpJIBl7
3wOhCSZNjF3qTIq3MSO+IWjC3Ye6gxe1Qn/Xk7d4d68lbFnphJPc9qO5S4JGsIM7fMQthpufpFPe
Lnh/IlRDEEtcDjGjDHmlB9EiMMg6PsusJ9j8eSdP6DS24ZgULCy6MzXMDsJAUCQpXcSiJG05Ppmy
L9OdrS8gvx+1cncFTGMVmiokhRiMbKXpitqNt7VdEKI57fSe4UNMUfC8fyY2R521C/EEHVQX6a9E
idw5bfiS96qLD3cDew8AXcCFkL79n73m0eQBIwe0PxdWYrFCRlRCI6kWknlVHSlAlugTL6nRG0OB
rAljwJz0xGvsrWZdByb8cePPE9EaUIqS2WLbXAGRd5PkBLXz0e7miK47tGuIiTFMDDVR6J9KwH0/
/+UHcbj05AN3/VEsX0U7qHldFS43voTx76rpFAUxYIgK+9ofjEzwPw10oPgIRJIIyqy6xmijZj3P
LfeOPCaHKu7jKX1cv/jtfKgIDGHfaa0dku70f96PCz0SCsVtBSOLupTb6y7s5sPC+cQSqOXC5WQi
5dnmmYbyH/BDr1bSuN/G/xmguk0/VeFIZwGQs0MkCta35UyZ18No3D5IQXMA0tXNvTlxXos3l5ft
cptmRVLe5sLBqWa1m921LlzNDK8lsnS67XEld7IxGV9FWMsp/Iwln27GbNZgv6i0n9qUxZf+Rjhm
PqRf5+XUatd5v3m8zxZbV3ksfmbNFrUN067g0xE11ogSvIv81/mv7cvqLz23ZxDCxqRqwljrJYyY
tNOrlwosttoMqci7K1LnNKxAVCi+jr5CXrLTahThKpXrswHcZHxb7jWsnNjFJGZAv4cjnTRWr16B
0B0zAUHYU9bvE8Aa1AvmKg7wnFsfiK/+QBipaQiOJ/YjaTrSRdTr+ED6BVutFclQfQACAcba67qM
D2sSqY9aC7uqcXVGQcbtEdiPSVdcedtaeuN3u6aW5nLNPzmBYJNUvO2O+wd/4Hboq95YDl283tMG
/SOYDV+rT92cbGRtSRLVm2xBp/+rAAAb82qBOBPO+rayAlYKzwLLrGL59m9tqNmc+no+dO+nlsl0
xQemO6i6QCubkiXEhah5tnO8e4XVxqtHBuxl3Xu3eeotdympUgRl10u+G4vwg2lhkC5HZ9czO9Gp
0pMAD8bGC3q+AgKZQwgnlPo+CvzBubByzPHsmxflwzb+h/JXVcpjIttLYk/AELTfG9lVz62YaKdm
HlMmcGuXmOc3u+MFwy8ocTNZYJifElTMnn2niAcMkZFA6W17FNVnDklgnb1f77QSzp8q/wCwTYtV
6SRmNzzMB8AqirVIyHJ2tnLEMeR0h1t+HiSXq7z9zrfLX8Js06FZkUVHiMvuj+ZTeBO29JUljWXt
1tj6mjFMpz2RiXiC7vx6zofNJs3HxkunXM8qt6tDTpq8lcO7zfBkI+0LksasWwizDgb7ePOlCBpG
QcMON+Yel4NnhIHjbUlbmdhFR7J3VP+cidyrBPlhsTHN0PXDXnlExNeePrtP5ZVA74L6XrQRDM7I
fE7UlWrDYi0Y2s3zVLOKIDwDMYCjXxwI1C+i9UpQo6tSiqffAvGO8IRbp1fxFAWkeWAcB9WuFkCG
QT9dQvh2duweDX+A2OCzgwlTM3l5YgLkwTWcF1ukJ0k4MW2UqzSzP4NnzpAVolJbVaRGUlOU8YEx
utTxrLIW4IEW3mHu+iAQ9IJvF+KgBEexgcTLbn9lZ/GYb/hKBUlLRon0jcWazzf/fD48m16G7kU5
83c+LmrMdSA7tfTllEnF4YoVh+MXJoXxZbHESWsCML57F9+jytV80FKuGEK80CSN3wOEm3oWXouL
M714A74z0pOwxxJmHzLuod8dl04tm5HjMinEE1yj5YKzm9kRKhGRsV+i35n3KoOdQd/4rw/PgkRp
jievEGP9C3bWvHy9kLmvtZpLKVuwMjzMfqq3Vf2VpPCxSFJvNEzALQFyO/Z2maljhLExMMuBaz15
lhxSoL4dPppPruy7bXFD1K7IMy5j9pxXC1vphvRW9TRWDoNYcKazzDPMxat8hiUXH2uUmQYgB/SR
/EP25mZBqfYxnDkotsqdC9oaai+sJ9nWrk11rV50lZN0ofDw1qbN4xejpILyKt34NAGVSI0L00w+
UwsBRNQ5lhAjtLRkA8pJV9zxeQfiXgNfZevDb0tyXL/2rAzcAdWHs/t/Jf6kgMbk3l6g6PkPrxos
nvqnSCfero5bJXkBqGYqFH/hd18Xj3v9KiCEC3DvMYRXqmEmt6DIEHb3ExgPu7UMTTbSEvSDRTRl
NjLuwAiTv1GPUAsCkhZGm09BsFQ5pmVdMnpZBJauEYzaI8Dalz+Yk/L+Xg+XEiz6XipOgzmJsdqy
64Y5aIvBaWl9Hsb9zLwENVAn9dLDGXL0Lzx+DeJvgjcy6Xqm7T3qpfiD8flOiH5AgYZ7nLadmp+L
aU/ys/oegiOcA4yN8SANIiiM7nxabjSZ+i+TlIu9c3id29uea3DQ+X+jONI3su0Kyn5hYhlnCj2Q
IVqAvuUMOrZiqAX7gy50bL6tYGSIKrZcR9gTEt/iENbdRsACPTmUgmF431/SgtWYJci5sxDiRTm1
mIgos2BTXuwXbKJvGbAY68VDrmDMg3ejR13ZP4AiCi7pG5W50L9v5JHYNlEFiTIj67L45JORpyg1
B/DAciMNui1u716ZDcuUbs64t9DsjYuBSw7nKCOwD6h5xoLwWGEVfObiE7AFI4t7u8C+XFYTJgFN
Vi590j9x81eYm5OWZYIFN7Y6GubLrqbvZd/iI7wZ/hUnGflLYXkVb1HAIdX7N9vD+Ba7rjc4eUA1
3BsNsa0F9irFz5ZvgCfdAoxA3+0R4iy9kWOpiWY3m7b5YD65jznBMEea/1lZkPmiF/yprERMe2Xc
qBD4QjbJPxtyAStlnPawTTe0aYq68VjNnaeY2HlwjRE+jnCk0tV4GBIA1eHh02hsXzbCGWGBPlur
Ejz7YCLx7xQiDC5451KqEQWGUhYqRKZh1z/N5g7QiSNgLxNoZR/GIYhCyLKmCZTHaTWGl+cj0Ny9
MdE6UZdLq09250fGTCHeYBOmUmogyj73EZV0+1697jN5IwU7cl33+pN+K0L/6wWdZhjTTL9P1NL5
Z4Ue2AV9fRk0wB5W36cH9MEAPgACmSuaL7sBBGUK9rEDUyH4fGGQMvozabAOM0y6mfbz39KrR1AC
wObcwieH4hO1VUDg6VqJfMqEA80ALIa2tnAQAt4atKQQmJM/0Z64QXPIAr12kvuX3Fclv9UKeRbp
j5a/AXTX+8qB/+YyrNwkY8DbQNvkH1f9BTZQ/yhHF8hX5CMkSFd9z0ypYmGOkIb99Te6JLYWhnQl
vXUangEX4oQPyMIcA5ZXfhE67UUlU0rnNK4aEpO6bDfkdyZM25YtXBQySeeJWzh9QVylLfJjYIja
E72ocJBeRB1IRptlHV2+EB4GndxagN2VvaCSx7pVU8PNx8tEhCe1Y4jq6Q6qg4ZC8/s2pgrftG5R
o5QL4BpsqhhHojN5eLLoovop6mcOZ9YMWcE5PQNT8tLM5zhsz97nKRB/GDaaXdW0jxEOLj2GSrEz
87vKt8RFPrrcbcy8jt4mk9R5OzUgSN9eDlacJ6vZ49ip91LUif4Q+toDzcth6u2PDWNwENls1cRF
qffwGRf6O4dvr//ih9fuNyKpS/eX5CyQtSHY+/ihqzK4DcS3igSPx7Aj/XGlKoJOpjhXkQfqEOwg
U0PQ/Dg4hFRfPlE07Ys9mhc8SM2PP9Ixg5XlOmX/M8iJDW7CZUgLKr3xzm9UMVGMkUGIQlG6Y0C1
okwY23psYD0eX0ieMUinEYAX6IsnwRLGQpZGwsAoLCqn5FqqLVl83+PkHrzoU4uV0pHr3xmzCfuK
XgKDzEQR1wmhoAcNa0EsvvRyxaXejYpvyPquzvNFQ4OcvzYhn4ecBa45Ixrl9lJO1tkA7wOoy30c
V8OjDFjcYNWHczbWGaPirW+h6th2oCAMVd1J4mSrQzQ6AoC6vzLKC7prxHWi/saLTkP2z7eRolwQ
s2cFpdAAMuevaRXgNO+6DKoABHL8aq0Qcg7zwvqqOxmSbHZKP1hjpJ3G642uVU9Ldc1d+RO9PNOu
nBbGECHKfg+Z5T8Ms7bWZYUbxheUcxWqY0PLNFaL5gyZd4tC0wmVy9YiVob0f+7LbXZcScAf/tf4
XeqLJVuAOkyR+2wAY2JkSHi5TyGOYFEE5dS09hJ1Acl1o5gi0NAyekBVTkWZcDfwUi2xsRtpnqF3
Z6ttKDLJhJS7uUZeL0P5wIAq/3oG827JaeMSBQKlIR3Fpr/Duy3aHQwgHYhzhncc8/81K0ss4Sc/
z6iaUGmOJApKJFTwqa//UKSZj3LFexkhCveWsa12rQg7b5DyonbElzYE2JTHDvbKAUh00DY91myV
bX9vFcmO6VG+zcEX6XMTzhVugc5ZdqWvnErkspMveVqJHaHbf3NR4XLGmvSZ5LRQXUVY0pULOGEL
Y52IEt3+4eWVQpJVbwHkhZGQhjvz0Nt4Jhu8D+4Ve0hfwyYouAaNkOfnCmY+qVPTmAbmOrb5Idft
N5C1pk7Xjh+odAjgMCHZd01TxW09LMmCtWEmEP3JF5m38o3ZURQV7pZfYF6C2fpZsol1o1f73GHq
QLePY3bZD96WQ7iAlj5DJ0ul9PN8OYJJcHkVgquQ6RAqMXFqkg6EF4utHZY0CURdyKdm+vmtVeKa
Oii11yK7AFYW5ZuBpyAEOtOYElskNUf7zL4k7avFg98YT4yVKfFN3PChVitScdtULwlUS/DIrHMf
DbSksJMtzaDulUaa5Ohe3qmKe9TRtLJAt1y1JR07W9pLSCtEEbEoK190/q8snMS2BUwJU+lNtUNv
kmeOGRxmMiaUB3/OCQp+oTSrCs/ADQqE7aYDsgHfZUZywbQIiYMPIAA8VnTg+JSf+vrK6S7bGmQf
j3PXMQIO0nXWb+d08teJqSaF6N6Ck2vrQrHq4CSXkzQB+e3NpD7gbxQQXlAvaCN8WZb2fCQgXGir
eihFXwBrYfoJSj1XxrtXEfdNd0Cfd9oPT5a9q1cUbsC+dOuYYFpKcR7229NUzwINhkUcane2+Ogl
MSSztOlf1CTEOTkmG14vWG1FKmoZeA2GlpfIhp0i+dt6SSRXUQmnWE5Y03sNU9QLklpdq5CRtAGC
IGvDfti4fq+EvfLvsC5wIYzUEa29uzRI/Q0nPYP23b8bRnv2IiNHqRojr4Sm4d+ORRpnMYZvvH7X
2htjF8qZeG4H/I4r+OMCO1cOzwOHjoOdoQ/j8X6On/gc3xSybyh4J5CML5HfQ18Pk1y700cMLoF8
M46ZB9HyFg9NpPV8pA7JPmmCDB3XcwnDW08bTGWi/W5A2hgocNhmWg8mVbk1NLDMRIWHhEbxKMQy
7V49hRg2T71wF9Htfg7TrSI8y1CQSBvLwYE1VgWELTHM7tT4IL+4vhS8T0fARbX9IdvEpiI7bIv0
g7CH91FFjEzN4aq1g1lQ1rQy8JgUy2mM/mr9WF8sNYkX83W64vilX1UMYcNgpxQEpIVEIo7p7tOY
Pka0OyOjNNnpcqbktnoUuUcLs2chjthnmoJyEgnGb9Ma7kiIgXXqQ8iNNvssu0vp7nC6PRxABsgW
1LY1SS0uyhKlWRciv7hS0z+kWH8REULw9lKltvxyXbYWhnAzgVbLAxQjkCTE7lGbo/osJFUtkmnE
tD1QqcDahkNWFMoVwoc/KKfUbcS6FTLlMeBGMGlPpu6bbqW6sI3ciZZ6IFuXJow5uvLkNbC7w76R
FQC+HJEYR/hrQdGzdXaPe+Jxf0NLtOAl1wzGiR0lnA5yXs0HQiYne9RPQMtOCxoyrfdl9yu9DeUf
EjFWQ8rnMd5ZVg3DJrXYN3LlP8qV2S8lQckSpmiEMpudu+gDT8EdxxQnkQEzMqX4RP/e1JXDMnk2
DaeVenRF0YQRB2YBLXAJhPKH1VSi2TltiOXxFFVM1wPZT8vLRBvUu4+BqgPTdId8ShjnvBeMvwS/
p6eVcM+5dxyqHpHNU47kMK9N00y4DitwxhY98UC7TIQu6zGzwC5tnLotBKwv1Dw85iWZa4woXye4
1XtwobmLf1yvNblUjjoyA3t4/4sb7GzAADVf01M/sptlNtlvuHSuVJhbL4ZJMrbT/euKSdIlhbrM
hsKolJP2kyXXvDtQiOu7mT/tz0cuHuZGDkkbqHJh2CvEL0wbOKJ9Xb4ukQsvhK6J/8A8I56vhXeu
4XxJbkLdh477GQDdLQvvb6i8zzpEGsY3eHVCaFpQ9w6NrGDUVQsyy6sA/fEF57gUmOLkM9dcSSrl
IDpjavhdZbmI0NBrBVQIRbSqCnzEdCeLMQaN15sh6TeP7hJX5nnSRv/3fO2GgmZy4qp8ZlunmlJm
qWKUR96gO7YgREauFn2WK76b8JvQQuj3awACTnlWhNDf0swzvqka9VsVaYm/itawIesGlshJlXWn
koeRRoHq9MsCEv4gx6qd8tKU2marXHYV2sY9I48MaZ7u8zI5WLelaAHdnVMc9AZNIk7bflHC8giA
6oXVJrCRYLyNOCoHkCbFQCDlLFZcUmcdLBpye5ehNpOGXh0DrT7Tr6OirSQxN6ybnTB8t7Zx4PT1
iO8ahh+IQ54zrBEg0vmj8e8P8anVZi0i1WyCKFVsa2IF864s5HYGjLzCPYKFEN5tnQsTUFirKmiF
3DZN7atEVymUDFD4CazTl+kyJa/TFCTMB/vme71S7Dqb0mJTojEiU5cjWZJp3+Ik9jsUr8lR4l7P
A4YwRkdnqQqCv6gA/sACS1rdHYhAtuZ+2NRqdn4zZxnFCbryrNtfLCoV0yDrlw/lDDbWKGztcgiH
UeanPnkhz6/zZlVRzH4ydRDFL1L54AMeSJ9jHXoFf1VNGJMQnRB86P04JhhTvXTFEpHNUHzKe09g
5JaKnHKMk2Q35rGTvGWVWEdtI297XvWc1W1KQSnMgGfN3RlR3oHy4K7xXtSepDY/pmPydQOd16MO
/mthwndNWDRc8k51UHggbTNMe6o4kbZL07GBcxcGiYkM9g1Y1ZNfO0qlnZDrmf0ZCaTZpWd9bdwU
i2Z+i7P0jrFzAGZ2OLOSsM4avFW6VUchlmiqPpfj0pNjeAzw6um+BRvsa9zUitDUeD4V1Y98XcRY
bdxDtjo0VUNQOV6HGMZDNUGKf3gb9lg0PI08gc70wxdwkeImrRMSCYYxbG5I6KPeW+wv3X9yGwNj
kcmPatTEa2Hkcb2gsm61pMkAdKZXlwcAaOewFn9Vs6rxuLmeKWR2MZ3DHQ6YnuiWbWZhS0giMYHD
hY24tzaebe6PwIX6kchYnXeDv+MQ0NOV5qaZC88JCUtUEmF8FIWnG6K0EAD4CUK8DUuripLAL3pa
BmEpxvcGbBZW+aNMHN9lf5Pef0QNf6arEYYLJQRI96cYNBvgTx4YkU62/XgOSB6yb+B923SDMbo0
KLs7kewYmscHQE+QgWYTvbjreU9MqP9hOs4h3i9EwFW7dW2/TPGQ7vUbzkwpLf93KqcEZR0zReTM
9W0sxHiKxUkcVMnNkirIRVI/XRcuUnwgfIHiG7YeCC8vniUmOlfIoqNdtmU5jfVGaMvMhEHlBSLE
P0cQS9DnsUee3pfdGrdC2CG3ZtHuDI9ea8I0/d414oC2xPeXZ5ycjdEFH5t0Z/r8bUns2OjS/3rX
lga/d+LLYU6Bhs14BNDbt6eLQpPAGHwoApNJbifEyHG5QQuP9Tk3ZYcH2psrEuQiWiY+jwx6pbRo
BpBNyGN3qXF+ox9JMo2Atlx7OyTsQdoJs0gEMuEMtLUcTbZLQIA2UoKIOBvgcM4FsbQcKxHKrc4p
dB3oopYaNt0SXgci33t+/HNruueZXDJstCqPPeItyiooed+QVZv86HqdzzCQTkGS/OK4GDvS2APZ
kTkPmma/7CVEe/HHTHW/BJQWsEMKdoylLsqA/lnzkBHnf16PWlwFor2eFgdGMweDPibdUgD/tfBd
6o6+86jN3gNmjevJ3gWJ/9hb2OD0FRaEpvg6i6q3FJRmUixjbo6LJppIipQ3Qi13t7pCvEjLDWVt
FR5W6jMZ7oUP/atpoSQrWoEy6uQumv0nQN7JQZ7v+jc2hmJ6+Q9za0qU3mfVgvobVwk709YJIcJ6
cwBLbPXc+WuZEl8T1SE5R9l2EDw5Au6KNZYNFmklhHziIvwdYYV8eetpDlPZ6bl707IhnJTRinKt
qUV77c5c25A9sYP7H9DMhIv1Gl4Z2aMh/vpDo0WdAdzB8IL8UA4XGww1dREG6xaLWNNtGY1bCXRG
FUcfkCmY8J4XCXmg/B8M4EtNRtUkoaZWFg6pNUdy8mHxk0L4ElCAFdpZ0DwB+edNvcPm46XBgVay
tgdNPTon/w+F9WXnR6wHgmPu3Y9+e7AJk2PmHbCzAfKUrvozUixna6hEgr3eKjPx/BIyw14J6HI5
14iphfpVfkrWgRNZ+Vrxjpqag++MuAi9R4X7Pxq9iL9qqxEAUIv23yllKgrTYbUtI28fN8NKlLIZ
AVfZCKI7Ay+5sMx7LtCaThDOTEdZsKscUkfnfSbxA6CKQJWABA6o8KtwrZnKB8/4dXhrH65uVEi3
r8m8cUPMwmp+vwo7hKBWwV636cKWM3q/Uupo64ynCbJNG+7zFPISjxctdHjiZmT9hRqjOauDJKPA
VOlDh3rBVLE2OtxIFidFjwzsojnC02DpP3Z56Jiw83uo+XwBBYdcqaQzfs4KeB8ADHzfixB1EHOW
ytubE0Ai1qeQCI75NvKkkCx5LpbFeAlKMhkCng/kjbCULduaAEV22Rj6FIR4Xoo0UJfPTxvIDW0/
hD3i8YFJnJNTrkfFv8KwoZL/7vzNeTynSbxHgRlpPMGih0t7kxDeLKnDJ282mPYB7nWcGuwLe9H7
CY0FIqo4Jj/vqczqZ3XOA2phenNRnCspp3nHS1C2YmAgbuc6GdMg7d0/yJe0x2Aa4w9OfdQ3JI7x
l4eiNayVV0F5wo7d9lUWIetvP76EJjuInCwbUYAgH0Lxe4LOzfhTbSFCZELpvngZ8bjQUNkHkHLR
bnCIPRbpyjMyR2GSfmdAxbF8Jy0RCqboa39PuduzMcjxNBD6N1I+fpKdVZc9sAwlQQboKEu05vxR
VOoolhetLPkdUHmMN9lgW4O3RXhM8o9Y2Bj+dePqn7cqf/7Y9bOFaS6D/FpnN+ji5578qzMZDizz
iZCzBoCj2xusJgZ3qqcAeBjG9Q7VvKBs8otOfJvf/EZCyE3c6yu7TmNe+A/tGUs6X4WdkjCUsqyc
TG4uman0LYrPyKLSn+9kx1khU0xvC/TqVFhZ2mUeWnZ4Dw7dJHzTVtGP6j1HX8FCFMh5yhMklqC4
sOg7/T6QoxATY9BGRWahAKucN8X8Y9iTqqsXuDpNNNdQ7Qens9/KVxFcqTr136UOir9G+31feevY
nt8aPg7WBDEPOxrNyGrOPQ+5qdDpl3Cwvmdy1+FQNC0EoHUMHz+v2uJETRpxxFVQ7gn4fF0yevsU
NYyWZ8aLzALdtIF/qN2rk9zxuZoEJIc7OcPKBmU4ldaxQCf5P/GZuv2uBLiYAX+OND+/8uOUNK8p
ODEqMgX4ziS8psbSi0cnZiccg7rmVPlmwiBFVaiOvsB65033vb82yF/3YywToXJnM268HHil4JjN
9TxdhVWQnePehqc9GPrYqHUWxYUABhVkmpsdCp/skgJSX/CGSsQozAGsfTqAf+N94CRaWfGsE3/W
19PJd+27F+weJmmVcw1fkGySU2IlY40L4lntZiQfd7UjrC6mC4W68sM23u9xFZNUWK6CCqqmu5Rh
RXEXA4BfxUlsGgIP6k2fYq4il8wtLR5B01oAbkK3RotEo+QLfW9m2b/TzX6cBu+0MJyPNSYYP587
HfnnOYyjogpo1cvVeFOc1FyqoSac/wBFj3CgT6RREfDlzBrtzryFsMFoI4ViyOwRU2xrG/5ZR2WK
UZ+V9yc7cENv8PCTn3Gv1OC7thZZaNSHN2aiULu3/rFRwnAnX/D9C+o/IJmpMNoZsEVxypOzIuqv
4ARxX93lmE4uhpyAeASu/mNI/SDaDW1qRA4ivafdsjwSzDvE96wMr0t7Rr4lQwmKOSBNygIab9cY
vMwb7K3DVNATlGfSHODlsNVBXHiC2dSKRH+CLqhv+2k5uTCysncy6y1EvLvQJugoWggYF5p/TrEt
lbBTPt6DS5/KDfFdbER2EZp+Kdw09k8FGNO+9YdvAiVjr2K3zqWX2BOsYuEfqlOE2uavLEP+PJVA
9lhSuVncCnUtt4hZdaJfTQEiBfwVrqrZXJpbSGPUHlg6cEzKqHnJxVCTPJxVh4MlQmMSnc3czl4k
kuDg9KFaTbVFxmyCIvead0lGH1lRW52972DhDB0RRMjPbZ9mAd+UinPdXXR4eNrP/qzAQ+CODjyr
QvPBw/TlCMi7kG6AT3vQRNHkbVDAy59mbGI9oBMExl6X/uZBrV/x8MPbdgqGCxOi6QALWlKNqL4L
ojytY73r5jGYEI3M1k1SYiGgijAaw09igFalZDbFK9EpjF/ZibrBep2UrHNXt7JJxogCp4Z73+oA
PpgcIIUos9y4pkvzlSOJBAogAGKj/wS4ZQWLSLiTs95qh/94W82IMgyBgp+my/ZbPGA+WOB0Uxj/
Yr2OA9smrrsQnlB7Zk96nyYlhjmFTYeKzgNsQL9e2kYVbmRSoq8KrpnNFUPlITGKUPvst6578Ryj
+cPtGfsl3Tl42uXxAxabONAgnDENRQ42xZnBre82k2dP20ebXLpiGGSAQiOqSo8V18z13jiIYjvZ
T/2CBinodebw+YzKhQ7Cj6EWAJwnTcLvTkTHxQbjuMR0WUCLIpcP6Lt+I74V09vM1b35cz4eSSVa
IjksmuEulMEWFJdw69/ycusr4kfhYJOexT+sKKSa8GJtyxfqkegY0PunPgXuurBkeqIBUSRhoP7E
lTPOIf3BphWDr8ij8B50L2ttCzPXsfWOeeF5SQe6p3Zhi+oe8xmIPDaciKBAcJJhf+7C0g84o3nn
syncLHmkKXLsYouDV4RCplfFGTAMB8clUBe0TlkT4vm/17GFAQbOYlsr5Lynx0+bY/v+ov0uWlXt
VFzos9wjfhec8X//a0/EgjC9rtNV/W2mFOE09KfL43oPb6HOhssKnS/Bro3i/YYU5Kl3tnM33fnA
iBwSxjzMn3jZpOjEP4MAgpmuUcO4cmT0b1IlUFVfOTSvUp+3s7htWTN6wclb+Yd8d4XoaLfVj+kk
8NHgN8HslmuB9G6DCO4TcroIM73Z1yF6eP2r4flUqj5hYinwChbXYuRg+qQQ1pF/XrSkzUOpcTpV
coVuTQ7YGvcU2gaw7A4FgrY4xmn5IyEB52s2w6rY5E06eN+nukqHV8D3D4POh5r2eEzh5yGrotzU
K3plQUiERR4T5IU7rsSjtZgLoJ/e8ZoZLob3AfPNN4JCmG+or+V9i1KjVpowy4kYi8oUrTO/hnV/
I2H1vFoFAY3VRtLqbzNWIpt3Bbt80uixBAWgqGCtmjpq7QUF9ZpCfCjm92diF+7afBOLhEUFmlWG
4c4Gbc1FqMC42jw5XDQ0OCJDyhJJm7MozorT5Z3GTbGGdOhNQ7tp5cyvWq8asmAPVXpU3pGBQt5+
JOPE/HFj7ebtgKR9E4xm1K6o5XQvwibCvvxD7LIk+rkq8T3SAJ9nJSabsFYTZdPVeTFYiCug/use
1KFDJODtZMd2+DtOo01D3wZtUKSXGA8K1CsZHEbn18GDs3t01FKfoJ02hvP4C/ACssTIKHD1dqtR
bGd2g+buD7E3jE53JvbcF318SW9IQyVIkn5KxYCH92oAV3tzwieavpNXbvob/c+apfSp6HUnjnxN
rusbq9UcdootKwEkzgit1IU/QX+3RhLBuRJNc7DrefBfqTrWzswJ3S1wI7OavAf8Q6mKasbrIdhF
aIeSEFr3Y39HkO389aGLg7Lb4tjzhfyF7wuzbzxujO11X1pD9pS57l0F6NjuznoszqI0QugADXTp
U4/a3jPodPCoGXd/VcUnePCXtuWWI8tWAqA2QTQhtKIM+G4ktHAYbev84PvYuMCgOGpyOS1BK3O0
vxROY50S3T7SWf4rvSbeV1djw8K371CuHaqlUESz5H1ldU0+cPSG8oDbavDg+f3HjbnaRek5amFW
z/wmwt1GTVNvUg4LzwXmEyd80AVK93ixGorainBdI5bbVE3xsd0393kiQxksyW7Ac4iEEkYWc4fi
JuZrp/ClMojb78/pvMO5QbdD/4DVFDpmF4jBv+tKqgsSuVAkK1pc68PgjOm1GYafywrs6Sh4rehb
4210nW9W7do9NdGMqre3k0fIX+MD8Lu27IAwSU9KWeJSsPgvWROa1UkJOwlwBv2+IJ3NkuUel5E5
DCVWUDr8eKaRkztts26DF3t6dllb5f9uxplEtrf8W1/f6+Wsam5ZQ09Lwfs2h6zfs0b6+n34FZiA
d7VoIGN2bPm8vhlRjCQ8+b2N6NtiM/wKdW0B0+qMPWhHh4tZ7K8YFi7v+xb6wKfx4W1luzP2QYtt
TMUrkaRPa6PEYBWbK80LWjArgAKTNAauRFhGkEUiwbUolI3cNw7syVb8j4QnnS/Ezx0NUiELwDTG
Z8hB1+sI0PclNUZAZqcpPAawbI8XOu5CWXzFwBNpcZ6Q8JqPgm2FfLg870WzZbpmNnfAm/FN/Pw4
049pqZsone5A2S9AVWVkeyTfd5uGOAuH6IQfEeeWSJVtSG/vM580lPRB9s/1gd2rBoOTpZirwHUf
NtLij4uh4dpqHxLa1Mg7xIktReBMLzWy/1zt3H7ACNiREWLJUGJgUKWsAqZdyb7r+LbtU5f9cyfW
4FnkDOvBVccBtk/2nuVyPhDW+AzOOOsky+pwf3JMTZAjKKpp5e1VYzq85kQZ+uBM/Emtlkz3aCzN
SRz5chosKvMxaGOa3bCyQYhi4GV888JWa/anpYrmPVUhM3kfuq12Lt6zLGREZxlivZ8vgZUGFxE+
hzlj6jbLTVULeU0dA2GDmWTFcdvArdZ3FVScxinxblO3whzz0j6Dosxlwc7mn5a7Tw710tU0Yi9V
khMlv8veYEjqQD2dFnCnGjDAffGbD/teO+o74oel5Cv7o44Hspozt7WojXSNe5U7r3AWlpTUo7h0
krjwOe50SCxm2xcUaFx2wPcyLCz1p5LU8owNfaqfgLBxLHj8tnk/L6+VdkbivtudT/Q2/N+GZP/z
NXnG1xSeTebYSA86E9RooFnAWQIuuQD8lVLM8Vq1+yKVPgPs2gQ8lkOptbDg/lI9dQ/QQ42Hej2D
+L+rJPTA5OAi1jeRaXYV8D2AuSs56/QXLjiSae1USRkdNg3Up8N9KDaDf4kXHhPg0Xj+5A8UT1me
nIfOGsi6QhfFYcOrDn4wLxnJtYJAFDH2skmQVxRtSfQwMqp/zi00rZWZi5E8VwolQpqx7jnPOq4S
2VF7HUbsh+oxs69s/soDgnLP5ljr4X6Vcl9wrJg/YnOBr03yyx/B6p/6iSdUfP62lzFAJAXGrFri
hWkWMBcB2lyVTRv9j8lHy0eF87uHUFXUtFM2+ruTKUYl9jxVBQJnmfXjD93gxiwoaGXdHi2dHOhs
RHBPkDQIHE58LNZTmQy1x1W4kCWp9ixLjv2E6YxATQDx1tzAap54TYGmDByVtgQvLPuE3CGcTy69
36RB9vb2qI0C4uEVozjqGNDXvONH2LQzmJc03OB6Af+QAv4MBn9fgMpI8KXBsg4UNilFUoOqhKdP
uO5nQNv9xUEBBVScYHkcx9TWrjKQ7WU9szJlDf5qKjXub+yzVRHrfFRc/jVHyMYL2LVapOCRAcG9
WypMu4lzlJRiEj9zkNwkHSMuPOPtX3ZVk6UQIZas0g1Y1zMoz/dpnC9a8N8/VDIm97yezmleAdna
Smcx04PqUQ9bp2x850hIGCCxeNZsmVpItrAPYbfJ5WNHV1+kTd7mFA8v8g38UAXjBhKbe2GySYdV
2rAim/1/yN3+VvrCU6wtP4WzxiZdL6AThm/VTOnOf2RHdNPmHniZTV+xbBl0Dwd0sE52UELws0Pl
0UQikz74YrlxZRvH3gt513PlIZ3RVZ8EjXirr3N0MMThYh7W0ypnL6O4I1tbjoIyaEbVerJKi2TJ
DpzbQjFPSjo/A2tnW2NKUvupV9dPzpE63U20njX7Z7MT4tewZZ5PFy9slE2O1VSktxuFCYJyAC6s
C7CnsbCl4ehWm91QD4tFWXioH2JMFmRgdRbJ16KGkRA4dosJvgjWg6kVPbgUlU8xLWyJ/dYrUtuW
lJv+FOAeWzhnAt3Camdc298YLKmoe2JawHfM2fI8BkkOHBuk20dppEJx/VaT91mBelddxShYL0u9
dzgsha7stwjHI3MQfAAY7pQwHo75C+UCB1FC730ReWghYn2gD2K4GeDCNzc5gynj2yXflDvnA9UK
ZceJ88HBmGH2U3B+lK6QCm6L2dnZpQcxssiw5ogZ4Ir8Xhs02AiSe4qIWTPrtMvlmG7CA566H8u+
/l6Yre24VTZ19wfx0Gvwe+9A7XsqzG9mm8ZCABysSfzZWgJmeB37/ZrxuZqE5nAB5ZCqXbEgNmv6
i6vtCLSR3ZhlXxAmhe1w+t+TXYmNnObYF7BiP4GM1KT+AXlQkhNSGJsriGwNRGZ41EsfAfy0owEQ
/rs7SreHiy4Pz2y0KR/8gZQ0vcyTOlMpimdJHzU5++WV7iobs4RkF0LUzH9ooLZmxeJv4gFfeEa0
uAWjwVC2WIFJWFzwOFM2uiaZh4N7HB6oLeNKQb6yYJAsP2mIpWIxfkWrA0SNdbRXV17XzIr98gQ/
wJ8By4LpLp5NBqvszQ+lVCgi0CalqKlI8hbWWghjcRgnVRMwdIoLVsYdT2BOuQzm44caTDbT6Tq7
A4TzvsQyPX4jzrq6Jdc3eVo2KY4PfgTtW1Sq16WCGFWzP8+4CLUeQX/RMnPE7RKRh9cJJ365zm7t
EljykxtGhUm8nAxN35sBo77oVUXZ2qKX7G7f8ifq7H5fq1INwAnWSa9bEVZsSX88543NwJEkLvXJ
OJ069f8mkKAPDAFhBBOOJW8qYcw3IiqS++FF/EPwy1JpyhfsJjOu/e+RgTMdpniWgybkWQAEO9Gc
aLSKQSE6e+2jHfyPcTjIENMABKdNOERNHS3ikLcmohFBXJqsC173/dDafVz+DTGoEM9bX55zw/hZ
4bKheRtjigTf7KNCExEJJ7p5fFOao0LsGz+OJYcIY6rLtQCNhmNzHTu+9bpvijiCkg6+WPqqyr1J
ZexMlgho7rf+knlZe5BUIjxgpn18PHG+BP551FKEgNURh+lZQapmfQIq8FXOJdfsuHdtma1MReF1
R2wCugDzzXdWFdRLEdADdqn+gtGSiaipl55ZoHUOTELgWhGDFAFabnN/+zD0SassoeDHgrpiCUrW
HF1caSFqtcICZkMHRndk/8sgBGmQ0FBmyBKHud9agO4JocO4VbN7u6SgwERn5BBhAcY0pZyJ198E
r6vglgRJTBL34ENSIcBKMaYcmtWb5PDmeeNm0orfPV3SWRrnA06AjIOpZZh99i3aMRAeL96iIk1m
g26eEr9DFeHjsvah89Qj1pUgWjAsurYTvPmEKxpFDztkLAtW5BXPZhJeWrYsdgsmH0sm4Q3eQ5pJ
zvdm1nP8gfBg16pguMU+aKQvrEW1a3/P5vHKLPcahJ7Mbxprt33m02S1p1dboIDy3b+hkqu6qsEe
Mgm62iLplN/4YiyVylQknFslw757ECBvmELa1VIE7xdnEMYxDVTMwRBuOiwU98M7NsK/yLKvkrpI
S5F5FiweKh8SPY38FMvzPa/7QCLAM/usUrabcT60gVnsHMNOToTOej+F3HdQW2DQb2yiD8OpUx8n
lCc7wrQ/fXVhqv0huEFiaf9YBKWnAzCbytyXOE+83fGebhfeM8aJpkjCFDNu4QRRuJDQoMhvOrFh
QrV2faDXGSjf/Pj42NHpJOtX0S7mHcGilIYEWv7nAyK4CIUMH9oMTdSG9YQ/z8iFziWbMALYhUG3
DGXDdjY+upZI8o1RrVQv0Ll/Q1QshbLsT1hze6di/wsMTqxCXaibkvZU1K1eDt0V6isGKzStCKhi
iJbN0ZLM4Z2gnSyfsJXkocGTIkSum4iRCzvj9DmyLHXYO7NJECZzHRe59htebkGixgZvMMpms5Tb
JRTr6WZOIrHA3JfibDSIrGIfHsQMstjXgZKkpRRrXcxa5BawEv+GpYvcmHkfxz7CTyCSfw19nIh/
i+CEuI+cLumDNZb+UMHXg0f73ktgUIwYCksjCaae7NOwPmYYJb1qBjLXbMviQRjImwKL2i4eRGsb
SoYp/7nOF5do1jg7Vh6Hit3pIOUwC/5X0Idjg6CMhChzSndlRbo8UTipzRt4tKkoboabG9Ti4VKI
1WtBd5Fd7xMQrlHijuqSdWhEfVPXXldgksnMTLwzx7p6OletKbd/bhz+3QTp3v5gqYIGn/1o5b7L
DHGgvJuac9SkPD8DaJYqrfI+BZHvE3/C4a7Ux53uXwY2rHhDUOlvBsuvBUhrtSGGdH9oX2JqCDXc
LPUTOU+yqAfh659EblhrmCzYXY23TfHhkzZp2Zwjb0Vbju+wyTuyyFV4UegsUqa9oY2KMbrEsrt0
oiaRRMEicgWofJaoXT5qlDM0UrmogmYoOXEDseqzp4VBe7eB6jYrn2XH74MJBzEdvYXCGRyIzN7b
VJ3DtSBq4sfjBnDRgH2PEkhgwv2InkMTymi/LXRLUZIdnUOzk8hUnGXHn3BWE+ZeSVQwpGWIPaxY
gCsFOiaazyjWYi1WPqq0nwjVdJbtPhWSQ6Ycsv/GQGBd+SNzbQEGY+yEQDG+5oQjlPiegg7Y9Keo
ZAIlrq6rQr7t8FJezYUkncmcas41HzGkgDynX70a+qDQ58UO2cRWP8Dx4sVTwbtXWIhzgKaQMNP6
cpWPeW6yO6owxp0QPbJWi8RHvIx0YlddjPJa7pwck4Xk+PbmqEe2Vhr405GMhCZi1HdXZp/4sedA
nBf8WwIf2GFrQKqQd9AG4DG9mTAwyEAQa/tSkbkQNQgp3FhrETfvJLbAh0bE7dH91+WQTHmqN/RT
Bz0WDXdCNpiCnq24t4O1sLUTQjaIJ/CHG/9CBr7clk6p1QKizDU4J+kzQihlkaXh1w/p0gtX0DdV
oR2TdqvFj+HaYp4O5lCrJGqasmEQXl+GQmc9lZkKcWvrjTuQnKf0gtnvIJjH5TbrUNzwKOqhfmgs
7j8ispnRzUspjAulQezdAElRIbB2eYnEPGF6lAybl0UHd1D0BX+VdA250YQrgMRjDmNpNQYewO1/
hgZJxplSr9daRHAwVlLhB+BUOvX4AW6lSsKq1z3c/n8/o9Yik6nr3zZjQFHK49UWij2EyiaPzpK+
cNpClFUkx12UatGO6rnmHm7cwZxcTuYkwLowFN06y+U5uf0oCUzzEbjwbq6xzshLMHoz1L2xWfqf
Gu77yOdkT61S5bRbvG18Wl6+OClQbSp6HaV8Up0MWAthcF0kaZUaqeMMoBB8u5+h2OOfB3CbIQBS
k4oei76aWzVdTX5JLkgDUjn3lcYPUAatX2Hrs+6hbXtTFH4H+wPgA5K0ZS4nj0L4IOW0+OWKifn4
s/Ge33tbpsF/RkoPHFf166FKT5wIS4p7R4UR7X0iaKDDTXO3HPJIZ/xZ7/O+Cmdag5iNE+gMWA1n
QGun4jLGbGzqYdgTccvnnousHq75sUkuFBBJkKfIOd8VrC+N2tnvGe7gAYaETKFbv/avBmX3NZoG
0dpgMGVRSmTIED/Ct5ntTVRjhmRA6IidKUkZRDWpnu64vvZAFYJ9zRh3/wyuecK8sKaiZV4aIJhA
t8UIj6werC8s6nY8ixDbtJsybyCbkUXJ+jL4HaftfUOwjAB36l4FmpgeLz1yXN+sxidIADCCT4L3
SO/bhLZJrNwQ0AJ1HgMyHtO86LN4H7HWUsaQi/28tBs/jx/GKQJXzFrbV84Jw5Rjd+mkIMlhr95u
B8YLNoROn9oKbrhLT9cXTciTCyQ7aSYnQ3SajgMeauy+gRytPAcnA4o3pbvwSkMWkHNk7DLw1Wqv
1GjeTnnnn5qjd4z2QsSik+JLcbIodh8eZSgfDGd0gWLS3ArRHbzsv7emhPYm4W2BgMo/mEVr2Bln
FE3AdNueh2jyUJfybb72d0Zx3CiqrRGrmabiIpTHtCmkrOZYHqKFYp9aMTFBrniIX6I0uaRfX+o/
3XLwHzfC+CkI0iSafPm8/QYM2zXAwlhJTzsZlnBaDeMFuJ4U5GgA2xeoexUsh0HznatwOKPLSSFy
7h0Z9lkOP+IiB35qFAbo6cFnySDTEtej5j/MJiEVHFeIUvyaIJn5mm9x/4UHNxycKyMtBeSdcDcX
PJp+L65dxyhhArPqYauqBmgrUksOUdE0J3l5LQFreSpN2biBd1EbGSnexVTB6QB/dMJml/0otwq6
RLY5RaSrRSpt841gyndoVafYxdoJokkkhSrdImjjJ1QQIvRmv4XYVo/W5wb08QbHN5632rYILdW1
HX8VjpnMONuRkqyV13pGPGUro3GEnm8/7f9wyu1FriGHFWXujNALPCz+hw7xDevQ9L5TiY3rvlsD
4vs0ceN3chdAHc2YMzs3Ss9h1Iynm12oJmhvhxAqBOoSf6gqJ8wXOh2Ni93AyqocrrKHLECjxy9V
4IgXZ3X3UnRhvvX/qKqMbUHkZ7OhSiEptSjnQI3NepvHOeEuPdtoUURJJiVDnAnjdctrB6SwooTX
MaSS+xIzJLEffo8zupKZgO3I1BJ2jfggYuRFfYzEKYtJv2FyPQf9SfZBH4DK0B+jV/xRNIarz5Dl
B4yZpq3PQJx12tfsPZxUcs2bwLMPX9aF3CrG9vcG6rhtZSn997CIg2w/DuyL5Tjm1ruJn9wL/rtG
jgChkf9WiYOpz5GKJoYmqbwJD96fmJr+gbxIna+sJX4kP3iVlUQK7qnr9SdMqVJTt+uw4NHiEnu8
hzmQun0ahKuksyIktCtfzSHTIzGfZVyJXCiCVAIRwgO9ZAuTF8yBpegYExSKR5vUIcPuf8GIbgNc
a55O/MSqpmcDIkqJVvKUxSX80M3fujgY5gz3jWhl7nB1gCKnaKsrHzO7Bjzkh7XbLZhd4MhRYmnj
D+BqtkI5CGdN6ZpmBIvPV1dDDE+HtoJoHfIFocHoRDkznT+ima3dhCIHlN/y+/Tq4CYddQuZL3xt
bm3ereT9HyzLwltdzFWmhOod66WNwIV/3Vl/KG2hdiFn1NBiTSZwt5L5GUbAe84O5ha2qppXTpTP
jhrnyhRnx4mmDFNrJq0KrLYth6xHO2xfLo3y0/86vThIEEugk+AAoExrWfdxkI/KaCEQLqUs5ZqU
riFIxlWftUPzP682iqBm3nNLY7EL4LRr1cmGvMJL1ZmyMnkZypdJj43UyUasDi6O67Oxit6LA7KM
gmDcgaDv7BG/4JsXnfVuruFvbhR2AMkRbN2omh3UUO4OPo6hHMOrymLj1cyh2JT6V08ouuyTiALs
u+wI4Gu7JQIZUcYOyPnHLd7EAEd9Eo0a+Az/lefHzpGU87C7PESoozru4BvMsGCfM+lGcYFEyUBL
Fhb4HBuCgJdbWYwhyRWOSwD7BtsuaPyilkYftY8JROdDZX41zIU36rrEQIBosnLmksYLBEIp+hUJ
gHpssjQihINigHN3G+K3KvT/kmt9kISFLdpybNVxth4QvyjUa7pcBOL7PUk4cfjIhztaGzCpzOOX
hj788/N6a6D1/8rjLPHdoBOKOP6oOC0i77RV4PiqvO79NmiaQabDzltFiOqvh3szvS9qj5ur0ToE
aieCkpXKfCjfIDkEz3V28Y2jJCgOakTrIpAtEwTIZJ7auENHrs1XnK2SU8xYowHyc9vNVM9RhIo1
7J5phSCX1AVUzeEug8cG1RFdVyME9xHmpvbERYBHrJ6Z5Wcdaa3uQm46xjv5soWx0fsG/HHBYFGY
9J3jJS0rQ/0FtB/+VBc/Du2aHCvhKRRu9PSwyByHY6yFbRZxmDpjmTez07uCIE/Mx0dvDVA9Hdh4
b6pMTQtjzAYo62+NEdKVbjRcJ6J7DNmR1UQplUQn76HKczjELtVByfykdlij43G/0vSDL7FmEFLZ
mJSgedsU0gp7HGihcC1xiPDypvoVAOBKB6ADodywNYGsuHguH0yKtnjna8z77QctzpEY2Svr9iaI
/1hM7Kx8E8SnbI9fUl+BV59+v3+j7ZF6UZJ2QpNHgSDvw1CfEHw+JAyoOiAty/bgRgcUnEk6QG/g
hLTj+iXXKyl5vISiPdfrB0pbzvBoX/gOpSA/JBJ0EVECI++kZx/1EepJz671Om4S7Nj71FRQO1lV
PbQbMqUPnxhHdzyaQdn8+Dv8VgiQSl6RGq06FCzujZ7gXZjyXfrs4iV/jFM8L3h7aWSEgHQFYAoV
Zk+NteqiV7Nq6QmMosWhrRmb2O+i2Qa0WsSwuwT3QpKy4GZ+DfOMaMKE/xjdvnqR12N2JUjIVG+v
1Gq6oGH5IlranGptEgVYCI7Tv1cGS9/o5lwSx2BTLdbxBJYexmf8luOuXU6scsvaNi/6TSBlsu6z
xhCS9pMhDt8jiIcIOeN59fpbAhhKaZIMrMtLBzwq+mlFsRY2SxNT0uY8djj/7U33PmYp5OjbycxA
UW7TvpvezdT0tu7U/YNWhJfUYOF/VJMlMDCuWWbRmXQsZ/BIcU2yADtut2JFNLQMFNdpr7Sn4bou
olOU0p35kIiaOClesMGAqSltrcwudff4pcUPEq09RNM38k3rNWJ/bIl7LZQtSTXvyXEGhgjF7TOY
71pvB8NeXVpb3kqPJwfAZgKt90YEU5E8plNDPRPJsGo+cmaZDXfyYmpxmPGWQl1mfYIcHpesD1Yh
IitmLFugF3mCVZhYXDiHuZPnnguuyc7KGJ8xW5j9KNLjLp33Q4XeW331MSx25RSx96lyTfR4E7F+
Geq191bFajpn4sevmwgbNIqRRYStIBHmePsd3Opfl2Yo4VuwmurjQlddHtjtaHZtjpJqE5CIP7e9
bmkw2MkZFcWSpM6J2RCGp3rrEpHUoI6gGk5E/4N95kA4wMYtnvDpTMDNrsrOl5pLVrDdxOYuPUQx
Mr+sNK/2DKTpfl8joKQZBOLHZkyAiwcfSb1TPb/uIEtZKF9Boi3kqXpHRwiQYbS25PxywWRLScHO
SDm5gsTP6WW20ArXo1emp5Qeo8VcvYUU1PntW80qo9dEcZPo68lkLGaZAIF/zZtdBmjzC8WMhjN1
WKCqzuWuqv5SaptKLS3hwn0ln6mBzEgUCGYbQsBzY1yKuWkwZU8UnGMgynuL4VPB2yG914A6hLBl
NcppjD2kuJ+9ag5LRh6kxd6CrMUXlgYUVyR1X93Uu/1AhcrpU5cxXMCmEGYesECIdhAFwxztcQHs
tWGznMpIDkcQsgLAhQOLuwo+VDt/3JCWK+NpxX36Eeo6g9XgAA0ZBtMGXhE7ypb5mDS3Nvg8YbeK
d68LqJMU5vQebJ7yLeXvy4VojAduuynh3QmUiYrEWJtoIWU2wu6vJ37Ld+peiRYYOnX0nMgTus4q
VHA2Hkg5HqXsfiNFNG/7t80bPTPYDjDxCfiUja/eB9IdRhkdlYpIdL3XmX/5wzR1M0pwpOKqgkLM
NFHC/NGfIfa97N1Aa4PYItJzIa6qvmMG8iNEtLfvtIiInCY02CDp8VZRJ/IV4/3pq+oebVFPzTtY
ZAQBQt0XLO+Z9ETIAn5WDVJWeREwvw+4DJQ3q/KMVZNW4OKeLNehtf8EoGqzyNZqgIpdtmXrzBU1
cSzptvMJUGP8wrtqv4xoo8LZgM6Fd9bs9hyu4uWTq1FX2ivhhPBij6xtTcT0+qtLZ2yi4k4NWqgd
oh5zGKokxmkie3G8PN2PZ7LqA8CZc6QvcWsWtVymQN07zlNBpcaKJwpUJyQSjlBVUB8cMlMNZeuW
J165VJdYEz2fOZd+lOTVEmqL1Ll9bHY6ZlnMJGttCkOonOkmB5aiNrQ5BYAW4EPpiv0NIvwLObPH
wylgCLrEmXWUK7CB+fO8qCJNZTYj63yEDZVEuOTj9OIu/w1UJDmdyonLyA9KHVTS1hjtT0CNDrzU
+IuKijm+YZI4wzCU/7/jbZsJudMz41mL93cSUV/+Wg7RmNj22bbPhhQkwP2dqY/9KGh9FnJobAUc
E5jn4HE/iEOOED1BXdyBdS0bqYhVrrpi4PTZ4fa5Lhl1dsvWRyfdxEgCmFyTNvU7YlQWLQpWPA0l
g81tzZxdvLYTwfLJIwtPskA96Sjmq8kxOzHpkcqjzooE90k6gUVIPfE6bVTWdsXk8968ckgmkP9T
QAFkDnlH1yZ++9xh/JLu0pyhoP0Oid3+spgr6vUpdyhXtpWeKFB0vBxRxcsKZkDTTA2EauukdvkZ
c0jTKze4mWg39xU4QBmPwk0SA70ehzS4QKLII24mGA8DkPPyGWg9sPznb4WPr1O2HUJz+Sd267K5
XO9uqcKdNjU07roTxWI1CVpCs/OqFpuMJ5QlZU5xPAlD+BadNiwEjLhDxscHXfyB5ykX812nrAEG
BY5NQYjgfO7Bbtue7Ez9uRe2j8w4SaDFk7FNbvyOfdx2vKql5O7qtHAxFE2L/VEmDEvWSt9+Lwsc
y+CCtkabvZtWnyw1IB2JQkiUkE7kkvDbULfL3I8PNl34ybD3h8H/kSA+HiGwa+Fh+rHoqmWwUlmM
u3BZ9UpzoxGy+xm78dRzcomOAm7VLn5iokNSsEL7OISB3dVXBWxjId0rmBpCmvKNQKzlyVB7+lr5
J1MEc1WTvkFYCX9ARaHrnve2V4AAbj4v09RbsXgud9ikbL/ZolmIEz7RduN+dp+a7kayE3b7XuNx
vT4ZyS9uCCyFqmgu34+EKpzKrWrC+s7dOPRBjfYUNUp6ougpX4sASa1VcwSA5OC9wckEQp5Msrh4
VMAzjjhlxD0KV1SXUjw08VK1BOUWEIj/bxvfKxj7m2uMhyozneSC5JlHN8PJLYlXnaMzwTzRT1eQ
DQBTCRC4uLegjEJlwVvgQHh5ZuqiOzLuM8lr7QuxQArFZRKLHDaQU8bN5FBRmbeNomz+QRBl+E4p
nSkpNUGWiyoXWdNBn/jQRbhFVpMCe9HjRMtAtXwHdsqikZXggVa9rXPO2fLz7PxZo68rkGBWmhQn
30dikyI21zaXvOFtHgNbeJA3UwOXnHRPu/RcycwH6pYy4xzC12iqAIzRYWfxUUh3YVlCNKPpT+PO
kjtV5k7uCSFCZ9IAMgCnPtpxyEM9HJHnTH5AjQyqySyFNSN0wv0xQ516TCniw0scxQcvaLqW5jhM
eSWd3BRo6DZgb/myIGZu3JrkZOzhvn32mgYXZQUHRtjVsSP22oqpS0KN7LaIN9vI+Eax35G4bpb0
38KyX5WXd+vXS9PgMAtwk99x9u2wsMi5Umfpg1Rs4b1jFt5KDFoQBx5tjZs+rDWXE+IsA+Hw9kmc
ZytS3mLxYZ0JTo0zMUXgjgPYKh9NSeAapjN30C8kvaCjWt+1OwplfUaOftRmhWy8gVlaNfD0Xg0H
VsJBKYC5MnkhiuipY/Fi572TNtSKOQRjQxyEsYqT3bqN4cU449YTRhhfOK4TufVkqcE/HWhqTClT
HYJ9iVr3p7N/mbVHu1Gt37pwExzsVtOgxAIGQxZCb0asx/sDEdzzCsmrkBTzCfR0+oiQS0pg8yCc
1KQfI6eypkxpUUs0NrcUelS+V2TaOGytwg2LmH86eqNVETVEJO639iBnMCShV+IdlYmPgzLDkRMq
BHG2ogSR+HufK2ArpMJETDtY2KwwpCGYG3lE65YK8ymFPEri1F8alodbXSP3AUk0jbSeQMb1wfRZ
UsbZTafEUaofs8PIzlq7Vos3v854FCewAXgm6ge/FU+Zpj2pPS7VHeiMUFG2sXOT2LewYbHi2Lt/
WRUYwCAhgXE3+3b85yquaJT/qQKGn6IvPey7Jib2gkYJRf7pMv4QASnLs8K8N0uQpdkPARHUqam+
1mdBMayur/FG4CIyY1Cf+tchfW95+ScwBKEkm50CrasTG51Fw7RqZwB4rLsDFHUnYyfG+uFHX05Y
6Sns287fUnPJRU/U+EdSBknOcw5WD6UxXBCGReMkXfm9PC5EsrsF1AWWBof8gyI0bOVKjHsognyp
CmA7N5H+WMxAgHZmJBzpXVUASVnvqOCM8L2TR1EmFvDBHY9oogMmjSV35lnQZ4Fr+I92/WKFdtcs
ixo+rr8nedPfipJ43zde8sCyInPuuABZBZ+Da2g1V6JEij+yX/ebVMrOVtE6gzpAjEhob7fdLaLG
v8yo0Sf77kG0Aelx4aGMGtFq6Gh7n/nQTUpKs/52no6c89D6u9mHbPjqkn0UEB8brqKthqxtKBLX
GGKjRwPwhvRtGNuMGEZMWx4gGoDNcmLiQf1yRcGe2qVSwPpmDK+i7L/xkuoGeRVpn+E0KHufOQPn
2rSkzETDwhArI9vZGERC3iYAH8IVwWCS/miqYl2o+pdCBLHqYpZSRQNYHti8oXCQ19DcZZ5YyFEB
yexhl5TITb67rk0u9tFuWIlG4htbwmgbLWBuurmIsNKP9uPT4QtM9/f5iy/wDOJ2e6Q74RG0L5XF
ejKI7TcBMm9g1jyHbMqdtuxGeh22M/9kE7YP3UcozNil0FYRLVQ0vCW08U38Kfloj6QLxYHp81l1
np5k+7pI0Mt+Ji+62kU70A5bTtgLW5QiPU40ZwxUzfyyuOF5ynw5csf1bOhCnq7DA7QN4YsVCSe9
wg8yjs0twQDUUdUMNANrHGYaNlCxCtPLGOvW5sBLxUchn7kfyVhZjdCwpKu+j17iE+Pt3/mzD+5Z
rRBDmIdZ9wMqF37XT8yns7la/IO1Zq0gcHGEKH2oq6PECrLOjmUaYt5gatLwEhgpytLxqhisNjRh
QdLx9IO23wd7UZW1Gf2ESaKej9/kM1j/RWf314EqrLLuI6Shb2VLRRZDintppw6FLb4EFOhoAK1q
eUywN6/jN1+sfc3aGEA4Yk+Nu7IDLX4hmg4TBEOvwgVo71GV2YGYdhABytX+egJtrStjgF9EEpw7
cpPj4M+CvepsnAblU5lx8ew0HI+eZeU+iL4RLeCdtnIOVKdN8UDeQB9Zghq0LFC5iVGWGwXYMe9m
vXojCZX6tBJze3yvihMbeEni+i2pw3stmvWqdu16vdpiWCpvOjEsl1NKajSKzR/sqzxmKZYymdq+
txBtTR/m9LFK5nxFsT8NLreu9n9jQqyWDSrlenmJN7YXrIRLNf/FLNLFxY/eNtQD2PSjnrSRR4vd
1mNAfHl+N7+TNzIXqySOp6KnGJcCO9Ae6v8e6irC+gafft0cOj7wReDHv+xqlgWUL2uHXeZzUH0z
n26giEnGry9be7/q7MvKv5ii8m3Jv3Ox2PhUNmfXMFKt5oAMtSCT6wRdDoHhxCQfJJUl0JalJzeg
jergrNmVWbUpKHzBia32MTL3Y832/VB43GGt3LPRlKgjxFHXWsaUncLwYvAwf3WfQwoEbws/oDu5
M0eR1RocwPuAfW/CoSVstyJH1aX9M4lb7gQwIEOapa3ZFex1nW0bZoGiIPkOwKq50rGcDq9CIfO+
8USb8s99S0JVoa8YQyXqDjwFmx6fgohk7YUOFVlSSHDDgoIjEs72luY9xVA0+/YdniE8XH7XPqeC
d4cFhlgkWYoPKOBh3CmVqrxQT8TTwu6zkOnvIhNeE3zyK+Hozdo2IAv2ZaBTW4d/Ap05BBqpOZWA
Sokwrr5DrOKIPz0C8L6HIbwZNFkjprV2FxMDlKW7Z9eOYsy7y+mPFKQMPLqlwHb5bKrAK7qbQ28a
TZGXNx9mXM79Fhj6Oh1kZ6ynRLMXAcN/x9IMjtbkw9WfnlJ1V71Dh1OZBOBUEXT3EjWYGrvoX+uI
nV2KS/zcxoKaYTJvL4GWlQIArXuQuSrzzbrBKJSUpS2OWbKdQUmtHWOGyWS1jz91JJCnbUeX/Jrq
SmPFQXnKED+UeZ4EO/On/pfDZLx6BIIK+mKYMT6ZAOKC+eHZV7xYvCEE2svQbdn8W4kN2lCJ2gHF
5HSMmmmuaVLl70gI5e5JiohtwSf45R0bXMLgz4ocOyxXJS7lhJbrTuMi1wqFPWEHJcEYRr7+keQ8
sQcZDUM1nkdbNPqE5pFpWOGSeCPaLrWIdFu0kXI4UVYp/x1ORgMg7hSfZYG6TQU+YDIEJV7yrNnR
V+2eGfLKAwGEKJeRdScgcgKH/vuJPCnzkCdNRlcQ2NM1dUyR8Lsi7gI96t6gopr3jaHbuTarM/Ei
//GlhLKkUZEINfjOVKVoovdKBXFoEdvb0Y4etZcYepsmwqDqjg9X4qdQ8RuwBRq1ctQYd5Ky1ssi
3BmkHuMWd7NWOfQib2OTNs+TwUcVVTASfkXGK8IjvulWPZ5sxfHbdQulNra3mUJvZRjAxihlbqLh
zXLpbh4DoCZkxzIyZmsOyC8bgs01YpvpqfacLfLSwxCs2kbwSeLHU/Ql2AiXDOESmKRX8ucPw7A2
mU6wox0Y2z79X5ad+Z9FDRXwYqtpV56/OqT3MeYc3rsreVpexFwRXZK1mNK/O4wDKp/nRq36OKns
nDaYy2xSQc1pnHh43khMVPXMDhuBxqRCiosMwPzXqlH54XKYtS3sFTA0YHgz/rVPV4Nk8i2InNEH
ySr6aXDWWY8TPwaKGUaJY2U/nBz0jNhom4bUiU6amJ4ngYRxpPK0y255YsGcJs9JTtIqijrtDvWI
5CYbbK3YbefiMYRV5hZF6NWBltJZb/gsezPwx0csuDGGmPQktS00qy3FF520W4l5ZdRDHJ22vAOX
a5S+6B25fZAqQZRwo0a/opuO7yC5ax+W8L7/hmXc+UTiGD6GjZRXP7OJpHUH8NbzP94P6cobD++Y
85z57TFBHgR9uaJ+MO+uYQL5SfVAZs26uPGjNPBd+5w/TJ+J6RUvbq3l7MYZSWUSWUZ1pIcmCFs4
pGlpI7LH9WV8fnNPnMfMo0aB9NXjnL3SmEeiAtsM59joigNPnaaTqcckJLO9osAnRMMdS9CnLPG6
DI0/yjlag40jj8MjtoS0t+w9BvmwT45NJVGkFPDWeYl4EW0Bl47cN1iwK1ih8JMtpu8hov1HKFsn
7gfZ0eIGvuWVdGotf8W9VVw3Jy+BPyOZ/Of3Buuc0lX+Bk/ZcLvYCbEtQip5kmA0CxaY8kJabakZ
Edu9dydrSPTdKao0ab5Rj8hYcrEGsvMrdMUgCIwBs/N4de9HOQHyfvl4KZIzsWuj4YfHXob1z6EU
SC3LIXkNb8wLsaE+fuoMgIQ6WScUph2nk7cXJ6fDtWrre3jGODQtaNuVUr6b6tRKVS5zwaR9JLi8
nf7MtI9w28di6zZ9MrrXYYIzvOup/vTs5ze+bIoo7daFK0KEGWypXZzwLbE3FJLU+PDC6O/vmz2A
h+iEbfy69rbOEAP5MaI0bowdXzZv8xV1XBuZi8CKbjEMzdxZThnIe6Mq1oPmlADLsnyRvwo2UNJz
Cv4TYl0CO40cW1sE2Sn9Z5s7Bs+3BAOLzudDjApDbSfJJcF4P6ItILfiPf0M4aFXAWVV23J/G6Op
ftEYbPgn/4fuLmDWs9fwqkjaqh+GDbsPqRdViu1rTf2wV1rhqRwptlOE6Mxo/EKrzrBWIfjILFUk
/dJa7NYhsMKxVbztOoG+qSsqmjLVxvIzC39bVlxnYE2ogeZz6UvYc7kWRs8P9vDz49JMGO3V5XSj
RvCwq5Ds9QWWSnTC1BQ2dfPU8Adry/2JZSnn0DVqslysumb2LcSQDdwo9ClVyM1aRmbAGQP+Legd
ZUpd3+X0blAHAD9Qzc1hq7RJFmo3lALVKTDIdlmzFKjYA7Q+gkOQTQhsI+CNpZm1KWux/Fm+zIf8
d/BXkpzfSFRsH4BZh2dSsFvorAHDhR8MU0NM3biQ4w2Dosk5LKMXCpjkhfngYMSXLTefQ+Kla9pe
NzggBuKus0Nadza4rmWFO+vmB2DtIgHu+2SLjiW6jhRxkIOjOM0mqe05S4yLcIKsUNKRAvFWzXQG
W0Cba3Fn4WuWrKdMOjyJ6aDlTc7u+e66Cy3v/FHYVMjs64DNC86JgttSdwd/gpbbMAS/53cxNYSP
8o47UgdD+NgteuIpda6SPB25FXQoyRKmdoaumm14jw/5sJdIjy/V6e/ZXcu5btKgDTqgx4gpYa7+
YULStSUeuIeOKu9l3SjJ5YLqAy9v1JXnc+O1qYIyu7sjQfEWGXnS/5JCvwDUfnfz9Q1RUt3W+Z/S
RPNH+A70Di91t3WvgOfCBE9MT15DUsEOH4crgtF4+q/WKe3mPWiv//jGSia3pR0gOcZTQ6/fhz18
Gd7UCLPBKFFKksjZCSSVGr6+nhcwXoZ/ehZQPpLOShC/7WHvwtRDsV8juVh+oexfhVXngSF2NsH2
xws092ZCK9+OzkNOZRX9Yyj/r1/1h8fvDZjcQg8fUaDqfcvZm5ShnYExIuXh5r6NWsyf2mW0LeDO
OjsmC74ymdi9ArMl0LQXnbgeuJNF3yEKOyWQtiBDned2u+pfJc96B2iq/Iw63fbRnL/mCSDCv3UQ
bnKTO5n1k9nDkKLtyLn3B9CVUR+pZo0MqB1Kp67HmwiThLCUk0xMu88RCsPGV+dzbzwDJ1QPSwgI
XHgreRvmxsUj22D59tQO1RreK+n2fHnWnO21izntF8QjdDacZhOJAxT9wtD7CP5jBuxVgixieGs6
tt6AyuKFjqI7I2jbe5hjcREt0zHkTy1OgKN5qIZXN5gPfxjSWKtl2hpmi4GgYH3kAYOjwLCGOv8R
gZhMYq4xUQgPrJtNxo3+nxp2K1TiKXkEhHyh+fkpoLvPSxhFroaILyK3yAX1yB3pD5MHuo1F78Z7
iioozbOGUzyfrpRtthXjxp3H2WiCgocieFzxWd2s3b3NkMdQIwmX+uXk3xRzn1i7FWzDCXhjJEC9
K5O/ggXrB8EX7hETgOsybW/FylwrdFDXEr0I1fyeeren5glE8vL9umDNk02KvIt89XaFlfox4ueD
UnPtJvMpRMLm/bwLbeFacd9DRYGokH8HqeFaTBq0lHZCBV07rIHBN2HGXdVYixP9//F7hWVIQBdq
EUQdVPnwzT0blsm/CFKndRxnDIbAD/q7+l1MP44P3qOu1gezzNT95CLsS2U1rHZh04wrR/Ozpfi+
uQH4SbjXB+sxZcC4j4fnfij9zW4HogPW/f9CAf94V//x0/yv6WCOaGrP4mBwSoH393xJP4aSbR/8
f/eWFIMp2JD3T5C0mDRh2R/GiBlKbIiKr4mde/Y8Ez/sptLiz3ObhyP+10DREUai7NJRGDDbxtUx
/6r2ozIwle4Z9V06jGM/Af+oSdSf+jtCLbo2kv/kKzn5kxtBLQenuN4FBpMI0Zf5LRvBP92zYzwu
zHd85iySklEuZE0sp1KKaPQ94Tz77ZYVhQrlz6bn4WQd4zMQ52/KsDpyRFY90WI5LIVCrhxGybVE
iKS33b0jkQqep2yy5QWv8qFVjNS0pEVSEspZYAGsrukQUlXfSFTlkwWSx/cQLzN3056HAUtTySHD
ERc/EtLe/YFVDJ8wJS1hd5SQ/9x3FuNeo8GqDbCDn0jo90dxuLCwnps6b4W914S/+JrzWCnnx3FT
GkjjaWqhnIww9cP/OgBun4KxJ71rCqotrD0qu68ChU9+zk+Qu7gPEGIHPrLH1ndx29yHZXy0PYPu
EKpW9eZAhFh/OdsDZ1fe1vgn4v0hLKIi2pnsi82KCJt3V6OmLEJfRU2vRUOJ7gMWlMDyG2I6mRMO
PCkxXogR2bN2WujDAXXV3ZF+37vVFUzrrFQuLyDJNKC3phYY+rQaAtblyAXXdLhtEuF3xELpA3Wj
JbOQ0A4eUgZDr4ngVkwBcUT3JRdDhgsezhsHpmGZhIcR8VauF5QTQgNrFFSuO6D4/mkxqyezw6Kz
8+i4yUHG3/z7bTtJJQIFFAq1GTOhancqtqbS68ZjMM4YS+/hVxziA1h4CT4+Ffr6/sXLpFTsZBEW
BF8vh1e2Vw9auQ67EFzDqLd+CzwxVfpErltOmfA0lYtjrIA+78wFPojyXD2YdmCRxJMGE7V8Z1/J
QVDvpZEpCL1bGnY7sClb+B/foZy2zM16aYnJwU6KAd9EzQRHDE7kPe/2OivjFlwFpnZm0/ZKkL6A
TF6MuwGf5Vpp5pIp1rXuIFSYo+xJOWSSXPrO+8V4or7LqW0haoQPQJSdy3fYWmUuMaVRTIB4tILH
ZueJvammZhDSbVZS22Hn/B5II4LWALQ3taWBI194Diyr+z5drG9YYJ2qLCZZ4LECjK/p/ez1Nh3t
DQRy1/VueHAeH31Mx8A9CXSgjWY1GCBm2ti+uVnmKUhkg6109wG4AGmK3FXDupobM8go/gizn/qS
abkFIja/BdLQCNkh276Xixw5hsR+wlTRUGOID6m6jgXWv5tPyl92cYa4AwFv6GDlYFQXVFutTRum
HZQ+w39/Xxacw6Wvks8ugzUlRpwUWgwb7CqRmWTqJbmUbJRlf09Czu608KU1WAOuY02ieVAQfrBe
Qlq6gO5c9DBV1FoX63cGjZQNXabaQ/RnyXT9CBKA+C6CE5Dnjvr02fXbB5a7SUHjijEsXcNuV6BW
as0BKAjC3tqx9fy6VohTCpPPL82srfaJTRy01nA0BcwNfB2XtGWVT/M8gXGce5I7tf9R5b6woDsJ
tChH9CjsD9WIh9QGh+Wuev4zerE4yyvHb3vXYuqZA6qI60pRhOlMA4jV9gByYOmzSJ5WSgpnSeEu
hY9Rg3tTlmzdwIfA2dv5KMNWecivCYXvXF5F7zH4iSEvKqIIeRbLWGZLpHIaalqFOPqmuqAYp28C
Y4ILywcxLKKCmRr/nSRXtDduiiknliPn8NYbCrgstRq+CA4gn7eXY/VBaLOHPVd4/BY+yxyYC5L4
jW0mycOER2Ky0Ls/rVaJLyoCJrTvJMcGHG/wL5c3NdcHmwLe6dPvljYdybOLIrefkFMER9IX3v/8
rcSrSUkyeSHCOPtpCUV7JvMKpMbNdcARd0ULMPdofOo8uIQgBM7j2dV9AXYfp6xFYVr1Lqid9xM/
iWW4QiVUdNaFZUUETDVgrBbYpMZ9Keey/RHPA8ee5LrUNw0sA3vQTofLOMaSlndWKW7f0tuTKXQf
q+Z0mnySn0YL0AywaNCQtCunzBA8iEvK8nH+Bi1sIz31oU4g+T2JNVGX86rPAaeqY5Cvc8SPMMUk
1qv1s86BgR3L+LOa0ie4igII+SzYNjf3XMBrc0rrLpZqc9TnORyHUE4P8httgSbYg6Lb9LgsGGZE
w6rNvphaohm/PciadaD1oZMXQQbNiy60FH3SkR0O6IGfef6rlhdVwdd7ZUkHHkGDJ7gUN1E80sbg
9pPcztRVtmnkYXD2kXYZ6oKGxkSmC/5k/J6FtxVxyBH/RsLU4Wzwnn/GMvlC0NJfv94UaVSkNGdY
b9Al0vewyXK8b5nwre8n31DZLCuqhLAcTPQJP1zmZOKmfexLenWPbAxtyrLPNdWFYBLlXJAYKPE2
VcPnQLSWgfvz18CHDc2JJ+RPr36HO6KvPj6NJgAH1WBfIz6ct6LCtLrHdoQfyroziKUXXxV/6Y3c
OSsWkZcV427axGxxqNwWqXIggC0/ysoUExt/0ipc8f9Z6BADkSB0qKKAFhnrbMqWFeIqamELzXku
Q8J+THs2qCcgJiGpcRtjhQPK4tN7U9V3XHA7FHQ+qaJMBKEO1Z+FUXU96lk8qLnb10Z+4JV6Z0xl
o0eyN9k2jb+XavJJM3fPpRW6d3WIyaIkG9qr5PmSIzvJ2tpa8oumED/yrblPOQZoTTMaxeS7gznj
b4Qna09YsKstzRYfxziPi4/nyTHyOW44mryyN53zKtk1HKJOsY+qNUdCXSVB8wzwKl9rOl8PKJLI
q2r227nGQvOBruabGCtZZm6U9yGzZ27m7j5hCEBQJgt/mVTIJErtkYWSAxWLE2FlTlzNTCLObrCg
1wnQIs6d6bnIiMfHRHNtTp7hbogAxHeSDd90kq9chn0Fuvtw4D5ntNDJ/SoipEJZQf6SKLmVnVXy
a0asJRVu0QFGh3ZSl+QeSmGII/FkswrU/Ii+nU2JCqoqFFKPA/dO2nzy8d1q9mkcOg2TKOv5pwak
pgRZvMoGBH/aXbwnx6HSJxObHl/TbhjafDi0JQBuWVykWxUc0FhTnkc5E7SOZ1MGJOOpFELv4pD1
CgTHFVI4Kw4R6gZ4XR2rOVhJaY4cDtV79Xguv6OGy0QhyIK6u+zppQ7S35YUzE64NeiSwcQq8jr1
etGYouxF43aNvyyjh3TAnEY23Md+Aa+XbToVeGOS8Ok6751RnYvGSEYY3IZcaSQ1XJW/TldC73nn
dJ+1L03UH/ccdvnHr9KYPXWAMuBXWQ8KAM/iA49K9Pc3OWFup5v3SqoKsgJhSXoGFmexvmJCuBB5
p1i1B4gEoh9E3uvHmwUXE0PZnmC50ZrcBW68pUYxxbHe/Zer3z6+uHrZ0BwMTs6sMReNN0RjISjH
riSC64XP29B+WtkX74zpZNBbxEMx6M8Is7G2wh8UdQd42rDn2sa0DKxowW284lhXxgp8oocCWC+p
jU8/yXJhaYN6Kp+YiwfKsWVzv94/nGDCpWuILn2DmvstduTccSU33ByHz54zQnWKFTraY0ewFI8F
/MT41R5OTk+R+8pJgkYPWfpe4O/MtQYxA8vOLrfTeC33DgQ8nq2AGTXPumkmLHSJaSHIApHrE8b0
QDygK04Pl8kzqAhbAP478jvQwiZDboxLcjDoTunWiuhzXqyBDFeFblR6fXzRhR40PoUaJf4f6Qxm
PTxml19Vb9ZSutfNrwlfUo2oywqqnugbeJhkOXDOGVZ63YYzqMRTmqVgFqPZ+As2cdYUOkTU2mQS
S/2dzgqGlH1XjrWkTW4TPz2nTBZL5SOP8gSApXd0W+gByPJW05F/iq6KbeFqQHNTQV+/0ZPIv+/E
YrQvaQhCjklHlYIcRW1g6tIbP7cmqBjQHGvb9rG3MiBscC+2qlmitmGyy8mXz/6AyFsEQxVDafc4
LfrE/XoiCxYCaNaAv0WGTvUsX+kv7DMzPmmVXlxwdo4XGWobnGqxwK0aDPjuvhd4npiGSDI/Pv/a
ksHRJX3z9o1a637PR7pZJ2C+90rrheatRk+eV847wTbfvpz2bblmvqhmXL45Jji+NB2AmA9aXCMh
aVcSMu7Zr0Kog4HnKkva+IPizrPuY11skcc5GVPx69AHg6tDga4JEGxaM0fE5ps2mdPq7n1bTLK8
rfjJD/yKDfo8EiVy+314Rp4jDM/6+2cOrS2DBVqBpydTu+xIQkbkLvTXrCJl3q16cluzpx+O3vOH
Tq+a4EQUhvxJJ1077o2fTKnd68YHM4GUVd5iFX+A1u4K1wNnOnzqoyageeHovCuKY9Tlm74/7ko1
rcqKMz4r2lTaxTBEcbFameQ6GPnXIt8xZpIU4K389P8jK+VVP7xg3r1eMyfPOO0QukULgGlYA3Zg
WAxtFvEKRGq6L1VdfAmud+hcrBQRYCBCYUsRymixycc42bVUqX1lDCdaUZGw+71Q9XjN8Fp2ZDYB
DRcj8kOXDZYaHR/VTiHGSdAa9gjgx0ciVEZIfrBSP2c56JD/Lp7solIPyxKeyElyZootVMMR7YIc
a9C1i0Xciu2siio/+hwoFCiL74FgtmvrTEM8TSfVs5vSMKtxa9pKhMJEs4nhoUkBnvUMgNnLNTyJ
WGTb+Rw/hhi6H9nbT4s4LlYg8hy6QO6nOeBazcHeEtfYNDvdj5YgvylNbhD9/yDNWB5IPcu7QYgV
KhUKR3cPjhMULevbH7dWWlSO1bX13bPLAZMxNJY55rob3PIlCqdu8OVkJ9idmANDVQz59au4vlAU
HqilYd9XTBQrZiHMMpE46Nn1uK4kLlHNn5SZBfpRgZfGh93YcLSuKJnzMhe3Sk+heHmfqJwSe+dK
0ho0iKDo1a3h7uWzm/ST6unrN3UDiDbltxBcbUsWHidcPTzoyeB+fgDmcfAdtNoAbPZDA4JXzsKI
a1r2qXz+novWv3IY88XMN/90EENG4mXV8B+pjREaSkmfWFkPmHTv/2LNKEX3mNGUMzLWjTApSABg
WhgobBmriha942Ufv5BvDgiENGz412YpMDNlqqfv7SAOASAAvM9/gkTfgt7ipVjxGxrpKN1fDrqr
/tkFk7u+MKnVeVbEzwW6gBDm2rRZa2zktOIpG5oyz9HVy5r/dMcJ80k9slIEN79kUKA4CrGMdpVe
3Kx7NK3lE+9AIivktuqKxjsC+gN71z5FwS9FsRDw/E5S44I6qzZIjLMRc92y1u7LbZnWagXbQNQl
iIUeb8PepggRsTOoVEa1w0LT1siUzjuFE2BSOsH+u3o4oSZvSWFMj9dPYQ7vXRHksS6xrX6ZbZgN
3DRB3Xy6QPI4QbzgWJxIaRPikBo19JDR1wt3unQI7SO429/Zn5WQeDOIIvTPCYJCWloRj0oJqTZM
WYOiM7ZnDjYXnxm7rXbzSbm6JRUxekICmr9NkHFCRvh/u+1RFPrCZV0xW6bA+F1c3T4xQb4nRgZi
fRTn6aVojzF+m5Xc2zL/FaRIyOLkQDqqQvbZoM4BdtL35cnWKNpp3hWApxZwZXh5QFjUOhlHu4J7
7jvB1bXA0SsP1+kX/1CdfkK8yAs+3axni4BeixFZ+RaRmodRodPXwMl8pT3YtlTvXBQqOwVf/dx7
eIJbm5VnfVUxpgA6vwYACh4MxGVGWLRTe2JZIws6LdmCgAscMpuZ9yRrGHkVYHPKDLwpxGEni2Vq
Az9EX5ToawHvAd4ReqipzqHXtaz9E4yeDIetZht4KuTId2nRKz+voPpXUzuLnRbCtUoysd16/QNR
OtkkEDhm9Upyl/avQeLqFsPxVGLJ6gEcgh+7GAcHMpunCYVncy0oxbM7DLQZkpe0MQrKIYHFwgx/
NPKFjfq3zpS7/Vljea4tc+mGyCzp91LzBuuojccxXp/Pb9UU13julZbetD67TdqO78ImKO5UvAQe
jf1qyvRJBmZKKhfmdMZET/GRa5WtHeVbBJuhObE4Vsz2oAJiGqWsVSQbySV07g7snTxWVCKQtdHm
XTR03Png3go1tp4ayYfjge7m5BJUIXjVx/32LK6NHBDzjHKZ4YlJq7vvlhYuyEOsSGT7u3oSMgVC
NMWKruv+CZUugzZoC4Vcm76Z0KnGQHYDjUf/7kjSC6xW+xV3Ox2t1DTG3FWBzBqW/1L5HHSwuji+
J2yxSYWRrfa6Q7ZfwWDU6FAkCGJUzo6LGyPd0f4RTkZsZJ7XhRYhhTBxKWwIcGRya/rqMNNilu1u
Gq960Js05GS/xVizCM3e/30kvZ3YRg+WkwEIPYn01R5lE/RRhWIfNsQcgfX1H0HJJg45UArppf2R
/Dr7asE0raDIjOK7pdB8G1std4gFpBVnTRB/SVs8mW/EdiKyyGgrfnvV918AMQe0IwKhlC8ihnMb
y3EJbG7RzcW0illRz7BzVi0RiypyBH+psF0f5G2OsCpDw7/+OM+8iWmHchaWko13BeviWyfX5U9b
mTYZwUvjJOao7eFXKp/rgmvQokeFwU9Sqa8nP8o4zMWNKVuucBnTTofBu57kqF7Fz7ENtVehoMro
PKWegNcMPdad2tMgVTtuWxX+2yqk65NgAldmqaXReAUOMODaNUgSyIW99J4gXdFi2P06562wJhzQ
+fwhe2p/6cIcUFqcgiwrcsTSMMaEC/uB7YIjntf6jxMMNQIuwsdZgbWzQp3FB+XNxiIGVWjFkq5n
Vgxtpm3lXgcFDFLaxFjQfkL/gReR0DZaqfyEneZpFGVqs+18rF4GBxPY6B9i47WmNERYSAVeiKMU
Chba/D2Pi+LpoVwnXFv7CeQwJMenPzew6eMaZrkHE1WHNFqUjfXC4wmyz9qfm/++8gpD9QgFr2fD
jzOkGT4JYrV6YcV1b+JXnw4uijbgwwZuqh8zJM843p9s841FKByw5ZmKzcNIiatpuLEx1hie/6gB
LNDoz1x3MxiyIwskpd2aJXcdDPP2lXibUDtWUCY59+VEcVvFT8NuRLlc8EwVCDJFt3SBm3Vw1aFC
+du7a5pt//vG7ofy+6AsI8dqigMFinUdZPXgF8lkUzB+pzYY3f029GvVHIotjoe42qcX9esbNDOd
YkpQV6kGv3jFyrvOgI7O1c7X0qJU2a/2HdQRNVlKcEQhfpDLS9eNFae09uxeUmyjQ2E0Xfj3j+mu
K07YVokY/0JG1Yw2St2cX/91cNWxxhEtOw8UEDQW3eT2Ejx7AgvqzyjLbJ3jNLwWZCHArAkutVdq
cRA+jP9HMiueBvg9swKTha/Q5ZZoVjso2AVGn7n0vmYsEumJsl7HMbO/WdIztl/ki6Exj4W8kF/X
ExIeyCBn8kDPfJtsAxJsuVH8X+jew4T6qeM1J7cb21oEL/4h70yDE9zWLrbmziSwoYwqUVzwKX5S
/bDUaHhTikdg8XvYtFxDgye27+Ap1RZanOGkwg0Kv4BTl0zi9IjaSgcovaokuH3rBgIdq27/55SV
1u5H4+tezcYojQki+BIo36qIyyezuqYqD8r8mMcXdRu6e7eTPRVoPB3HtSkQvM0z2Pbdt2sbrv/G
Kq0qmCzsyE/NjCSwbJorVVC15dPuX7xZesTPdmF9EKv19c1spbIHYnZehT3DxD6w4p9stWCy2x6b
TR2wYrwV2HmJ7QC6gWwg9ExR1Q5zIanBYNu4G/s9bTa4FnKHoedFA3PyK7BC5oBKnydQhJcOB11V
/oW1KkTag2/c29SxZVUmzy5eYkdSCF+tV9Rtp3lBi0029FKI/KP3xQKpyccXlni6XdQKBwLKBBeb
ugpyyF5f+7SmYAmKH5ZdwavZzPePbry0IWe67d4FBIkbCeb7c2Nb3XrL9wWtYsWWrXFAzSEV028o
f5xkfi+1bUrxRnlBnVKCqGXixVQkkCFQSGZYa2Y0oiE6+HIRNk6yaKF9Lk2I+aVzJ+2xYIIkHFDV
lEaYYXt2rj4wk51WgACUoWcW/mjZ1Y2QfgWak0cnfZh7zxx5G4Wx0JgSJZjRyZ72Ce5P21Lm+ZQh
iT/NLusY+DKzk2xnsKExu3zIe3i8n0DRbmzXWpZ7TBI2r+BC1cYFqhbYNnMr91deRHzmlCCMSUQG
Tm0X3vK0/w9xrRXhxY2OpNcYpD5AeByL7dDSf9aJ8oSeKFlhFXwnzlQ9PDKoDdiMP8Vt4fB1DM6y
qv6eLCVanHOTLK0Eo4yNhcbi5fLX9WsgW9zKqeQk2BBQUls0mOPdqntyipHIPiAVtP/cIlYr9RRu
Ufz/8uosoaIG5bihkfCmihZfnFk/n0ZZqLam+Pbx05Pf5Si/stLQOak6n8HmNe1GT43clPpVfVyH
IMr1PesC1j9/OaGbnlJMTpKIoJ3vtF11npPRdEoktF0JGLzwh9pZMmHCPxt8VfwmToDimlcyrzPv
1wPyKDv/cUIFFKIl4t4fqOjpMyGho/8w7fpujDM/x16QtdC/FmGqqXqr+jJWP3SuaqvjAuSovYGe
uq/ohLAmN3qR3OQ+C25n1sSn0w0vbeZ+di78atArS53ztANb/h6pGxPKSv5jTRrIodoUjv/rr8T5
ZnlAdxZ7ffd52LgoJmlN/YPi+ckYkBAs8352CavYPOW6RfQP9UlC4x3iltH1by3HDeJVDGsIr0PX
pKAzRVxNYNDkhYocpX5sb97pGQw4cs26ZYng/yustk6L5gBT8+G8Xk5fLNcOkOLjUUMzkToIh3mD
S9EnKADfKWsRov8eRM847vy7Y8WOvdLz62VY50yJx9s4aZeVDlqo0hQMIqS0Mom8qPh+XLLugaum
MbZj23BXxDKQxAfNY5AKliN3XpbjgaFnkrb0xXw7ShymAmVvgS7PneVvgiJHoijDtpnh4dPfB8CF
zeUEvlDHeL0f/7Lux6ZxjZi/r9yBJXVmPtKcp01PFKITNdNcPp1p+PJIMjCYwtFMxgQvHiYtF5qs
tXEwtH1Q8eSLZMFf6XZpZeXIYpcrYqa5oOyvsKalseebmFCi+Ap3kjFxgZCmhPLtHY/bDrzioKEp
hGt7NkVRQBBltU8/P8dOfZpOVEobfnTaOOB5tp5K1Z+JIolGlFHkC11MsB4QmPur5PUnPCwRefFp
vZfMPd/8WQ7cs1xaleSdX9wYw5MUrDNp9+gTBzLWF9KqpHfvIB689K3BqpalKGx1bLivQQxMzi9a
Tm8hNg+TUTTQkxJ9ULimz1R67txLH6d4lQvhBYauGeJ4ENB76Px3VyQCbLghqq6qBuibuqVJCNND
azKk1mvNG54sSTbPOsTpNEkq5IGh0GKN88DzzFv212f0EXP8vpEdMhrprs6J+CZpkVOrXO63EzaE
ibNXCenXu7gCeJhYy1fp09zDDyXG80tM/TG6NvSIRFcsy4oljNKw4XjIJfPKPmNCdnO35fih36Pq
pDQ6mWbilyV2rk0VKdsLK7wokolU64ZQjdV1IQ3+aia5Mj7nSvAGl69KNVzulwEGSguIuFWlw5x4
QFdjw/jH69AgFIfZqq5Bw+AAnWQgvL0y3pURSoFKTN/4a9QhDIeCe1TRGjA7zPHtH2fkCsQwSk9P
oWR1g/suGR1+MUJJVBE3wP3Sp3weVsQMotxbn30Eb9UpBFve0FBM1WmnhrKk1Yo2CRGo0G5bRUSd
HQYhPfiqN3V0ZAYk5UzxQ8wAL7sQ0yRjgjLKi/Nv/cHQmDAzDYKzcIDUdV9gzoiqMDa4viYHZ581
5btD8Mr0ziMFfXAwFzYT90ShQX2fBPgLcQVD2s/S2KhZWZaXhJ5OcM+tyY1SzT1yImu7Ly5MgH4S
zGMdD5rl02rja1SB7vCVNj1NAZYnSX1z10Ep4CzWxwuLMbwLV+TmYdra49NNI7TKiEqX4NTYXsiJ
Xh5oMeSbt0a74cpbb5bDBbx0N3DBouv63HaJoiybVmLFk+XH8BCa/SJ1yqRx6EFJy3py2UVFBevl
gij6xBBn5y6o0yO0Of3jj6yGdkcPCe5h5Dm+IbrLD7dS26cbFB6mBEitinZvONWmr5Oy6Kkj2j8w
gDiaSOMjPDdjl9Um8wNAakOceys6kWh7OXYHaALa2Dz5lyNCT/1iNOPIeoQgHJCswjKzCco+3WQR
15l0M6tORpCI+qTbv9wv4Mj89uW8vbqkFOiaGyNpNYRUaSNWPmopNK8aR7aeobcNZpr+RhDne04L
WVGUAHKXKtPi61ctVMsfMeoVNs8WCFsz0hzVNrfWxmrgqthJPVIc1hvI8OwoXTD2gPSbonZbtVWA
jNLoIELCt+hGYVBq+jljQ2ksaha1yNFSosmwnBa6kPKe6GR34rVM+TTaKV74OzAA74gUEWLrAICG
nQtnMVNswjdO8JSeTw5fKLJT6z3yhkNVBZ8PZC0QN6bXT2BaCdJdtz3BheUMcNp1zcxY5jvScaPa
7VyD5QkYXT6TpewHiBMnhv0yT8nZT3tVm30epUFZAE0YDkGVkMO/72kQ4f9IsbLZthIJAF/+HT7u
MkARW+4D1JDPbZ6ShXH6UwO3o8bWmyJmpeX5AmnXiGqgm88P0BoAg3Lt0VsYYR74vLEqyhNIv4pN
XG9b9p0QDkmpM1i3V4YRny95SxbN4yro6qNE11mwVZAeeOM+2HcaLo/ydfLBp6mxzR+ie640uwRI
3Ltn/NKh37HrJ5ujezpCQtxyf6OTpARQLgxVOhEVIZobv8P1jkpFGzMjX82QuRRcQMXZaR5AoGM1
TrcOvpfCHGalDL8NBEeJxcIwM8ZoviLAU7WvaHlN9NpXo6MEyrhH1BkaZbdr0UEhDhW6Hgivpq7q
rLaodoX+mo1RYVbTr8jYFWEwTnVgIHM/nH08mdCgGLnbN3arzPUClcNt1R4gwM+2ByU0O+8bUYG1
T7UbxRt8jP+c/uQsh9o3NThwFemzEJ1/gg+lSad+r0THupeRzcutUkTmu9BeFY4d6gZEk+4NTugr
tcPSfIR+NjAWhLfmTiU7qi5cfcH202B5egqZpxqGd2t7ItHDkLcb7PkN/ZMKLH7l7bzJcFd/84SQ
K5wFFPcwUucypEBh+7L+4G3IdXOUpyFUpX7Um/Rpy/+hg8zcbncs6iM57TXPExc5D+1pNjBogLmH
ASkSXd5sla17i8AxWyKGWaHHR3SwWReBicUJL37rg0V41Z+u6mInuKDtXvS8F6b9cFlX2AwKxlUR
a9ZQZtHaPE/erK9WvWx8+yj8Df9r/V6ss//nImvRCtm6NAhhjNzb5za+JLi3tCjC6wUtHUKj8zcp
KYDGlqNwCKC2InB9RL9v+gvKOMqiBIffA5TlCj3wMJx9HXrWnT3Q+O/IDlS0+YZe41L46AQ6yCig
kPHhgyC50Cj1ghzkW2/kat3HBZGD4E4BCSOl+VwHhujfWrThuaQcjFBFiRWQQqVumUlfHwpbOOI1
e7tkE+frtdzknHkH3gACHfrmRc7+MjTXFqBrVbUZ/trcKmaWwYxQGCechBWLcYBjx1TzYIfKvv1q
7+jzLfrMLPm0yd1EO9CKZZYIkIGkRXRxy/maSpkGpB24RIPiIRezslu9LAw5dxg4Pftrm1rG/P5g
7I7wEb6msdQMV/yMYTxQ4uG1mPfHKp3DN+O6WDnJN5JOqZdYldUi+iuEC85BzogZBl4Fn0U6e2jj
hfOl9DgRCGwBzHz6JZapqzZKym3K9fRwvx80+YeNbfqUyoLt4BdsT5XMxBVMnSNRFSW4c5iQ99Rw
7fpgm/1iWoVd/pkXycqT33M/E1MoatrXVZaQTaBsCZ8cl+Vrg4jKOh7DK727jYPqDMt97FrnBE+O
1k9JQz29lY75lUfLnxS8s3PLZTJ6knDR/WCP6m86Do97heWyBuRZRsAln/nyx+WOJxRC9S+hYChm
LGNXHB0sYqEHRzZrzGf6F9/hp4ETh0W14p/IXM61fjmqLiZ02018uC1bax/TFy0e4Ja13hfJ5t5f
WjCpPJ7wcofUwlAEbflbigDvRmRmEPMsRZm2dNpKLQkZo9/ziWyqXTt+9F0VCDKAzBTbXb+PZZfq
eG1XuOYSyZPPbQvBN9ysAf8Sts4/6MEIDlzKb6hWFj+Zwv/4vPgJyukxXtGwDh8PftSuytzKCA7Z
UpjvLCX1/7SS+8ttE+LFwADHt8gvSE2Xqp/wPzSn/i7MertvZjWJ0cQshDpfhSm/irlja/8njhMa
G+5rceY6vNcfEj7rfHzciiy76BHaeBDRYeJPH4WANkVLOV7dnGTl1tu2uRCZIj8Zpw31mnid8g4z
wyAmlqZqYY+oFhv0EgOri9q/rF/8qJswRpNkUHhFpvLA+sRvEN34MpCJQ3OijQ65Ws7FHcOPfbxW
/5UXMRGsTPfbHwkQ0gp9AnWDCYzOKgUNcF7tEdLKUP1MIh2GglZgLXTD/1BssrGgnCOSvgHyiH47
XfAykjx7zsX/6Ny/A4Y0x4udobASn8yz/T/zU35fBvcf4o0uFhP/uYQJG16GclGKpXsCq2jHwiaC
z98LnhWVFQvXTRW5wkWyd1uTJwFsU+osOLF6j1JHHv7nRiJDJKhhFrs6yfsgkQST/hNQuAhXEiPB
XjSCN3TFfvaznJFhF116Bdy6NWsqcr16hbQ0udOtivOW7q+cMvcNJjqnRbtI1dEVjFEkPy0hLyk5
sdMEHeQPBcsbZSK+MUUjOGDJXs8H9LjbY2ip7Rq2WUnXmJihmt0KZXdjty53Ffh09UNkKmeSEQXx
n0OgbwGo+mlH6u/h0pElwzTh6uWHlTIuFEIjWffH15SvfMZvZ9fnU3ynpVWQPoh/yAjtaFH4nBPn
fvh0MntOtTLw0YI/VzY63ee3F2v5jBq49s9uwmUnOuhBj3wunKOzm6/AXzQcKBp+boKfQC2gMbQN
6AMly6lIToclV7Domc2WG1QUUtDtLSblrMw7lAxuuNHbyh4QbOQtvG9DirPYOGFrkw2sbfs9nBLe
Dqsn6f/7zh0pkOmUHPGqhDcB5jO0hCJa78CmkOvRFvp6C9lR+zMASTqlJNgt9LseNzuiK2VJghbW
BykDFRA4g9zQvSx85ivAglLEWXdZzh5RlNBwMAhXr1bvCFKlc+hv0OMF4BfcK7J+73Y075zsCd/3
SV1dftSP5aLkweSR4gwsnuPw507PQr0dCAHFpwAB1eYRdtYRWruSQwtOCoLiLKtil889pUvWoXGk
IN8OnY8VLlUocHKhDrrUzce5UTglOXx47WR5/n7kkC0yEKY7XlZSKtYj/kKU6Y3bScSFlpJMyHIa
m0WkO/xVZfWKNfdpi6769YdTWlitQKRuHpjexQ1ZQ8FYN0/Mvmf8Ol+reZYB5I4wywT2+ejRTomN
Rg2um4Do6luVDnVzM2U5xNB7SA5sdiBDF2JygUPSiBg8HAfKYpVCeUqh/igIZewhyBEqmr4bnmDO
ROXZdkx+USIj2G3F88ZWrpD/HCDmHBonvyXaAvPQmOI3ystBW6BA2XVLSjFGuvBn6KxTWLIBjV9e
sEWWU/faoyF5qT+/lwgJQ5G6gjFsBkysUNi8sIUUL0hahFEV1ADL9Gh9l+sc3FqyGyLuoUw7xNa9
VqQpDQPnRkfz7nOlNwX81hHLQxToPre9pKA37OvhVbg6/G1I85Gnb+b6I+AHpK6n+COlRMc6Glw9
G1owMdb9tIy72dOhYSjcJzDbZk2ufBtjEFL4jWDB1gC8HpeZp5VfStD8nBWeGjksWAhXHx/mfvhE
O+9e+juaYUrcu9d4wkCy9ODOq+kLffAq9UsE9z1cvXq8PWzj9rgcb4Fv3FlDWkfGowy9+8kp8v/k
//me65tRvNk/PLGe93QUuVb5uIqQW65hY+mUX2KG/SrgsrkXwC6NWDp1OaJESbOApd1RoTOdPa4h
V8PhMaAvS/mDJZOduBkqjLhYzaqgAv1ncTIlinVABaAZg3NnDrzLEzPvKcST6sZhiIMFoutKl3ok
/L32a+EWyfgjw8J+tAa2XhEXqQEA+82L2sGVR00jIhiBxz0wwLFKbgJS+WjQ6UwPR0Aq+YmuDJuX
xbwnDPh3vtN6NegArxRr7g1R6pEnIfK9a2Ahx1I4zVncF+hE8+nJ1RFGGhdXfZJV2sCTdVUIxeVx
OB1W3D42F27To/G3dEZ4FNQR7hUDVZX/2KrKJ5WOHJVCjPjYZtO7RiKVSbi3P4HW0GxUUN9kXX9W
RFYH7DFwYiJJHk7j3Xe/rItqlliGic39tH9XfGAHjWMV2EQAunqt+ZmtDGPg9+3ZspFpbVplZAz5
mc21va3P9RIqwiF4eeuyPyftxHqCyiUSjlFFNfIFAEwiTuG3EXle2HCBSv/KQltHmkbb7Ow5hPsQ
UwDaMH6QiLK9aj/i4+5bg0Ht9D3HPkS0DIsX7EamdEoRhzT5MetefGa9M2bSrWLKNSH1t617qDk3
AOxjOWomedC+zN1LWa0Drlwr2MTPsI75L+1oe/9NpslJKuplQCkGZbx/MDGGYEoo8jeps2qNorqg
qvWOw1udi4HFMtd3IoCt/ZFqXAJxUxW+ztrYP8ihqJciCrkvTiXQFqOjhr87IvTVqw1C0T3dYRvB
PBfwWS8nYYCF2aY0mP0+pBahZFUTmRCQbZC/RO/WhMKqLNqlvpUJ0JoJHI0hCQZbpYyn1gZQGH2L
L/Xp318+LjtAFPRZ42ixolHV7klcm75BkGmcgnOYdB7d243MtQcjpYhjVhdz9uRzjNUk6KmGo5mM
Z/ObcAiYv2AnBjPzUDUp6sT5YC1/VSLY92HaRtUapc/IZBJJIGJXJjH6BTydi9we/kQCRE1OOlwU
KBtrkTIK/K2OcttizC2AKV8cCyiexQ6poeYmwbcoSVn3KA6giUcXx+NY60+Fn1CacOBQuZQPSj3G
VOu3Cf47QmWd1wMDyjb34ZqeY7qZUa/ld8kRsx/JclBmY5VGNsx10Q3t4HuqOs+gE4IWrRfRemjc
vonet6ybt2FzKh+UqLLvTfDEvNOcS+WlSLwACrlzOpOoahKjcVe4yBJqdmtGgG9osb8Z26qApr8O
EfvhY8+bONUFp7tF7eUXEwIasE3YQFA5VcGCHTz6siLdrugMUQJmdX+McymKp0wuq2+k/q/yNtAY
VapgYxzZH7xJkZcRD/wcHJ2pM1wLvACdP94d0fiqO0VekP9I+iktwFq19WInpAf5lui6wQG9lQOB
1AvY0S4C1uydhMOLL/Bbk5jEwvElMTnZIrjEc7F5BWjb7ax6iIwREVPEkS9VYRO8SqFxHUJUAiQ4
iFv+oVgZ1tIH2KDSewgTNlN47Oa83ZIrOXtlFHefLYYZ21iD21grYfe3C0/M5kwgnPgi7OvvC7LC
i59H6iFzoXiML8s8u7jZvmxTMLD0lzW32uet3iZQ6S0TLJTFPUV2b77F3rc4OQj11dTpz8ELt5r1
k6SF8w8BDq8f1HevlyjL7LFOHhWfHUykpeJqzPEgmkOdt0Dt4oUqRk5nyxwC7uzWuSq+q9YHfqPp
fsuQ1lsdCZ3NYSHNbNjstV5zl1FNAzQ/aD1zuSAr9vinXIEEGlMy8j42whCmkljNjE/kB/G0cBrg
ztUqlAFdlzswQ/PHb5YNnPALseRJ0wwIdUk3VOCcNCsFQ2NptvbLhHtAsazCi0il5PNOEdcDdh0z
HkTMtMBfpR0itE5VkKEXHF6zj9Xjqurdv0AS+txkf3cxsGfkHNbujUB4KHNM4xJOX3uOpE8n/x+6
lkmkdYFojTGbfuUTWt0KMaXE8NSrbRicr7lyIuUNbR26CL9eiCazNmQqlvXOHxjTYyw8zL3xvywI
RzFZFzRpqg9p93dkUV+zH/H4/8NJ73Ba0Fy+ulOO/Yn71PWDih1rRGEOCwDtxyFuK8IRI87cVtIv
g3IE4wtzk1N18nJWu//SpsU2ULJJNd2wfkrNYIBiAh6wSNtZrZ8Z2YSu7wk1+EV1nbsInrWf+M+u
KrVrXBudY/zQ8JLLGIgOE0CmQKiPqXWbRmY+cjPGWKf5T+8tfGV3nV+kiL4cPGfBQB2sk9paVGg8
PIfdCqGu6odKftKx1nfCAAaE9CfG1RN6+efSWgXSHZXNERsyrz+jsTpEXMvMZEAAg7FJwbhzAtOE
l/E7kbs5RG6zYfRH+obCqy03y/VZcgKvYzr3z80i5xldpL5tx0614xe9RdHFnEJnWFndXcPV1HRy
cJMqy+GnTxB0MT6Z7rFdNe5P9kUQWkrVzRx4d3DMW9vm1MTu6cVQv5jl/4z7Vus+gJClR2wTDR0H
MGEyurVEdCpQHovzKSPFnM1FOep1rycotZKtwwghbKIKavxjDWu4QP7W2qH3qPT/hQYxrBZMTmYX
RQjmyO0EatAcaJ3NPQFuzZvvM3sPCDSQ7+oWbfoP0UVaskv+KYIM6EcPv7bAKAfSeOrjEmxKSXLv
8L1CS72GHbD7btBV3awiB2ThQ96PmQ5SHll9Iq7ngs09FeZ6VUcdAF0VWbBodPNdiLG3DoKMXAHS
AeuMOMvTmNv2GTj6ZyDzi+oFeeRYhQzK50RmRHKt4dsB6j45dGayOitGIXkdC9kN1Xxzm5OVnQOV
EmwS9waYLSsjCKv5/SzsIGh7U7ItrXxk995QjvZIp7JcqbLUtkGIUy+NIiraxBK4D3Gt5q1NC5pa
NNFCAssymXv/GrqHkf3geg46A5eNTjnNRLrPv80QlJaNxkYOj/n5ichN8OA4Kbnr7fnYxsdu5Qcn
Ve5G69SudmtMURpudLpZi5UBjm8webT1bQNSMEdACIC8ZRV8ccZenH4dtytFXQJps1mRAVSx5dTh
nJzzvxXCy8GX0/IJHuYoff/EE9ktwZTkVNO00N2zrn5VsqhBWTWdTzZQpIp3GDgDi5VqbtmL8xs7
xW7W43t4AmTiA/OmjgBBmnX20d6s92NcgVsrSfVGb+qvVI75ze4bGxETaARtBuo7Nmg6Ouu2p0ea
5DZGpqnCaokdmO9wyCJFg8vuOKyK6q+mDgFhq2XORGz5CMXF6OZq49Qo3ogGcnzPlVpKliYOXND+
9as6g7kGHwyuEZ/fQdQMcKBoWtrzZWiEkuIs541DKMOHOoW9gr2b541t5k3HworC/COjr+BiqUKg
K6AVKIyDz6Yh9Gh5M6NT+0xBE5Z8H3wXrURNLatAEqPECP/6cgDjFRnx6tHSMrC/Pp1Cc4U5dDd4
GJF0Rx5XKUkH8hFFNc9Lj55YW5zAuQOfzt1g/QC7B45cxR+97iQYwLSoc8bD3zOf+vRlsCKiWHUa
I/N+uRcVP5vTnZJfG3znOz2g7O/DW3Z0BcMgF8cY1ommhBNculTVcTkf5l2flE6ZK6+vonYD/G4K
rMmKQzLY61mU920UXNX5mc8iqUcvINRqFC81+1k3OJxvabnN/VptzLgasxIhnpmb4J3foAXug84R
f/AcRvjE8q2MTVuCWbNFBZsGAsdSkil1TrCLfuXmxuwxmvrfP9lS+f7JzU6zyVvbiISUvMtnR7Fd
P+2yNlnvtQdYNi9yFyk8BDL361hhQUCrsR15AriZLevkMOocEVTTjTzKv+SODGHoKKVNGkfTPzh0
V/KsDBY5ui0wjgMGKi6WGowptFt5Ij2ida2L73j7AfdklYH6RyBAIQXDqQc/bwNnIckXfZEgYKQg
D3By3PBLy5OuwDATeO/JExAuq4LACmZqTQBJQAB9GgiH0NgxJRuiZX1UOe9ePzN6tP2/6k7QJq+3
EgTIim4gn8guKGFd5kWUKSFWO9BZHbJRkziBlPobDstFuTdvDbYMPzWPlC/PNOdGCeAaX5dNLydM
4EWGYIjRU+pmfzFagkpwbt6WJiwpNMBfgUkIN/OsOjUGq0pePco7l4MS3NZBl/BWQRetFDhz4tE2
qyx3Ch0tHafM+JGVXemm254RT8Wr08bEfaWuWH8yPpuLraIs/H5CXQeOwcV/bdufzaBYyADnt6Xi
B5bPfiHLJ2VhMY6NJyc/tedO8IP7F5AknEm8IpGFuA2mhfklsBeS0TESiockhPNs+TNW3GU0ucl2
5OCYKhhzL0ZBhzr3D8HdIJXzRfxn8qEMxMrNlN41UDWaasqImn+43MJykXXL0NENMDe0KJis1/iM
/o1ShfVuatptFSMEPypsYhWwyRVQlZyZDQQF9TdP0gqO4b38ZpxtiAPK3WgV4tWlWbXBTZCfR42p
8sX95O4AzJO2TumfgwVbNcwMmBOjXvQjrnOM/xtdqwbemQpDQ6ONoCkNAwa9S+AxUGQUoZGKsfKY
OKTTfVT/6qKpG8OuatHjqNgta5UKl6lbsQJFA/KblGx3gD/mdHGpLc9n/k4ByoJAujn6voiXplPX
uC9P4K3CCslHjfXbU4+aABgoE2GcRsL1kS89Vykd/+d+Iz2FjlCpP2wD+KSqiqy+6Rbt9PrHVgyz
VLTOe0kfr4KZoFpFV0AymjUuWD4Hjq8B86BB5Db9dpOxtgmoFkryVIOZumJprjnbdjkcEfin5+lH
pifaS75HgXkJoz8rExi06kkCjyxuOG0iMU3uQEAoNvR0ZHXWHYYtCmXeNPbXERfl2HkT58EbYIC9
zUflg4Pwwh3TIxnANHB/LF4cUmQ30R2Iut5jBA0QXXL4OcXd/SAq7Aq+dLsj0uovNhFrxCTXiIOh
ElNEyW1+AlQCE7GaKYqxGSBN3TLs0KMXarVtzEwUzMmO0oICUPvpiPnlbyLjrsCbnW66pbtyZ580
PEo0/UPnXthkMSEAzaBRJzhNtD9aIEUMyP5bYKryqYnBBjr+saUN9D+SGy/vVqaiODB1R5HBb6Yb
xpsglR9kUjeGEf+aYokHWNvlrH/4JQWNqCMJqACycYbqUW1hUSpRbJvyAiM5C+ZM+kFWdmXYhpHy
BoriC0uGfqS7yFAfON7jCPymgWslR8SI4/pktN2im+zVFJhriD8OIBatKcKuFO2n1zGiU8U1kISh
YCLUeWCzWV7LznjdUbo4ZJ7s6ewRcHbufu8RLg20zWWmAFlfgdf5uJeJipJXQ59P0/NDjsBLGvsN
Jx2zWbFeqy/gVrurf2JjQiDYdc/H1+zzyUYI8xDZOKRh7lQU1wrxGgUCAKuhK7qh7+D7q4xFPGNM
HPs82E1XWM51UFOza09Ymx8a9qBh/r4HOL1voByegpqu69HpxmB92d/IA9Zx8zFIHNze5nwuzc9k
d7MzNiURaj1T1QndzdKd+t8l67rwp01MZTCwfZyNNd9HXE4uJUNT9Zvy7bnpeMgPI2rx8T3Cm5r2
XYLSZd1HeUu7wfKQ50IxdX0TLnLipR8l8/AZqCdyOkcrDGpa/g3LUrYjhJs0ds2cRxWtH9yitTpi
PnGp7PwDPYiebAt+DKUkOHPJbLcM48avwJlNkYpP/PpfObMLwP+Z016DM5Xwb6boPxz/3mq8MYkO
UybviVnRkIlMZeh1Vm9arYYJvCaRos7O8o+3NMxpZKURXzyTyCVQt54p0BmM9mmbA5efI35Hd5T8
off0WbLyYRYliGSqNCIaqE2qlSZEX1kCQlNQRbVi7aUiZ68povP7EQSEagWWqkT0Xio1Yrk8Rrme
xuVZ4eJzbUBspT86J8e5xKlkcmHwNfg5mO9RaBm5Zu1lq5cD2nGIehdkqfGoXCSP84CPlyH/xy/u
NEUvQJ0DGZMuOVUFpgWPrTJLlAOJKACkiMXldbDj2d3TpiteCNedqi2ABwx5uf5liB5KOLKVctmM
pthb9vom8Bs4R1TBiPMCSdDSTxNA5R68/Ea17H7pkZvfzAZq3rcLfLMjkIzQvFucxFHhruBH2IM9
rDDqqVHv5EnMf7XiLTD0O29LU0Q1kbwtzRnb76x2XXS7qTFTK1brBnnY5J/usFTNOwBke9G+RN0E
8UgBAqeZ6+f8LDNa2x21eMREHoOmX0ELikkO5euX0OByRgRsLMsDQ14K7E4wcK2tReeDs1H8JueT
JeYa8osj9HskWVrvrmnYKtkqG3n2Z7ERNsDR/VSigKLGCFAbId+Y8bCe6yaSYL1S/glsLyf8fv4o
6cluSchWvD9haW0qcdtzrmNLRaNHxp4GColLAzQJbuJZTD+vpL+1yhfa+LanbQFP8Xmank9OoWzf
EG7X3NThosF9wBkrxp9NNxm7ILKphf76k0bz6Pm10T4SEXS4r+M9i5rXw7+YErXshFU6BG/ypp1q
QmX/bS3vdkzFmU5JYTfWtL+AKj/VysWohPXUa732clw7hay3mxAPa2nsLs0kYEc8WZ70uD5EL6VD
HxDnA4GS3Xl21wAoWHpovw0MoX3prU/v+wmf02UIqksnKHiGav2PeroiY4RkLSN1k/XW0/h2quVd
r4cv2esEH3KZEvuobid3XISE8F+P3BZ0p9Nq4ldvtROpzB1B2yYR3ukadMPjkp+bPPtI4BEJ11lf
KgKW5ylfgB7hgJ20LqvtKhu7cYkzjChOF59F7QczBdGFHsCExa5qhzm20tjVE8NNvyeoz8CXD7+H
dzm3Hn78lFatc6bT3OUEnHo8PHmVBa4EBAnaeT1Y/EVDr+oUNpQbxpMu4Kp88wLrE21f9fuHcohk
n7wBB14Pn1i9RFpsbgZkzjB0n/Ew0sf22bSpoTMWWKeGUw75HrDxM1fIsQ80coQ8hSnKfPW/CMqz
5PexRNnvkc/klzzdRrlaE924A7aKYPmod8G/pg62W+4RfggphVjI1K45iW6VyXIdw6XuZaucuQI9
PFZ5lkhCWYJRfWQLYW3rRJvETHaqmxiz8gAB4UjnQr89a1Iwk1MJHtO7/3FG7i0itBE5yktzmNQ1
gM2DE2xQtdZekyaVCkLI/9z5LcdQFv5icsbH8lOobyubO29MliK6Kw0OTh2XsPse0J+H4beDXNDB
khqFVlH7VJNsyyirWOczg/UAqf/ueUvONDL4jjZzHHaIdxaHuxBIVOukPTR51SuzeaVIVLJthjwW
54uLwKjzZpdMSKMZKluD2e3OtsEO9LUbqvKTy1CVzDYnsLO1X1Wr42et/CDES+u71PkhiQDNYINy
W6Boemw/YJmGSjaXwTmeN13yhynPw54xlsw1FyO59TONrQRv5gkYAtaa/UMHwDsfwo1nxZDZIP9u
kJm6zpAsClPvI8H9yHp+7/tzesfU870dOuA9aOOEan/txpmxaUbtLiNZuDoPrXIVw4Fyo327fKz2
nQbpHDGUMqRh/8hUfnMW+nYUlXN7S6K6MZc9rP+uDfuQctfedrnqD7ByZIfPDzDCPRSdv9BwWovU
HJVYWf1tJps0ydpIFyVOIjcOzjLfYIio7Jkgn/LsQ4ny1gVwhAPlLXkmM/HzGw4WRVESv6CWJAUS
KDrkEbndHNQT3UUVrvtSm2VG3U5KcufPvKvk8A0SDd+sjEPVZEYLr+8DqRhfTYVu6aPX45nWY3P8
yrDYCj2b7rRcxoBidw9oQTtovihcjAv9ZicnFgX/bmryVW+CwMwddiMSM0MrPD6Cx8xeyW5OJyTf
yJ94Vml9hW21al+fnfEmSoBmS6j/7ghGCVnS/+eqxyIC5fnQYo6q8VWBK/3qmqkJgW9Knkz1Ctmr
+SZlgEaWdI5HTKVSc2M0pZ+Jv7o05XGLyPRp87JicNLoLLetdP0bipklvIhPxqmTzLN1dwh6ihXQ
fig04F2NfEB3BMb0GKCHvs1bKYvHgaTA6ZoYt/7Mm0op+iJHS08QBP2m21TsrsXEp+v2Sada9yrF
oTje2shTyBdoLrITXff7tGETwADE4VDTFtl0fCsfnrx8Fe7YivdGwqB+6ShwCia2fN7AmVsDjYmy
qXCpVfO0Jkbw9+7GZKfDo/QQZjSdu/A60+0J+Tjp8PEABtY91TVAlISaTsq+OuLdXr37O87peD6Z
Jz7T8SkocIVqJHoq7doNg0ykgogii8oOEpl8TgokKWJZ8603g97OhVS+oora/xoNYpPpcoeUi5c7
IYLsgHSsqDHwbtymel7fOdzcwsZO8BN/ZDmsNndo6WHvxgsEnkZYYbsYQaqJvXU0Pa1s/XFHGKks
AYO7zb3O/VusJgkZuSns1ay9fl/S3MijHC5vKhH33FA/O/WGqTLb7Md2T391ggpD1ihOKFdMFe34
O8buqm9XkXU+gNfoJuuAqJaYVWPwDV1w63Q69YhZbaqlmk9aZ4bmQxAbabbNT0TR12rQ2bnGEWG7
ErAGdwIKCmwABBmJh+JrLjUrTiLmzJYHrsiyDnfjiBh5561uGutO6NUuM8Oi0V6X7tbwgUbQ2qAq
7GXEwOgmHVQpP3FvIyAxlZibN8fVdXtFCChK7UYcFp95BIvyhxOWVXKGrAkQGRmdh1parQjbGEBK
hTo9Tp50mLb8K6SeD4pzl9+l+Q+ocxI8XMUCYCm6fhinuU6JI8bSSdi90lt1zRyLQQ0bGxbQtSab
o/3GtjajzmgZ9EANSeD2vKPhObfHHRyDk+AL3/+pv8itbR3X70x9McJvd4r5Dpa/mKcukHK3F0Vt
J4jFgPE0Z4cC84tLjkhtMzFi4/CLRdryVi3Ltz0wHXwVfDvwT8DGCVVrqE7IoieFqMVRJAVpYSNI
gfpon2os73U03t/IhSp7+CBIbsJSk8AyjqKOP99pbdj44msamXJRKZZTouBjc1xnVTi+/Y2skRL6
QMshyLg21wCNL2XilEfJctf8ucz4V6+xOx8xZcJfWdzF0GqVZZuqY1icfi7BzIvVwu4UvyJREvlE
1VSRxDZzga04YhrH4Hipn64Q0wqPrsFAeokGGxveQPLS+7Hkaf1EOtIw2uWAJrhBib1Qx8GC/Kcs
PQ4vXNjq3rDItcBA6Z2D6qbjEB43HHV10dp+nCTFbuUvu5DMBfNo5u16nVufD8xDRPhtCVe9yaGd
eU1f6SKT0R+mx3PsDUGqkeU5TMDUFyHSoFXf7d1zXqehfPZkb6Pyk3D/JyNQUGZ3/gb+JIuEKtVP
TGluULpjeY2J+dZQfJJq4mMHLAuDL9EZyqjGXBTiJaSzwcevYVC+LS2XLWTpjERbLgo2U+4fzA3d
5a0aoUEnMthISIOe/Ja8l93g2T8EKeLZpXuVCCAgZgNNh7HGvQU2tODF8XHOH+bl76m7EtzcuVHD
SokKACq5GhGwkuAG+hDRLjVv+UOON1h7dtLwAQijBczInnxpbMY6q20kqTTL1pkols2msObosNEA
xvFUY+86i6gk9YmB8s+DoEzJ+97sOCaFnwBuG94oJuTqJb7++uZBiSWg9bnvJVz5EZEprDvHNqz2
KTwUM6CxBY3CiAv7UfrE8bZ3AIqf0x9HWRrHI9cC2yLNvpx/THqm7DU00Dwxhgd5mUyCL1t+YLtn
LpiT+dfUeQLUdhY0KU33Ecc8yEf7vMJMU3hRsVYeygU/Jq1oU2+vlJICFwMCDvraZ9zaYLbVFomj
FeeDsPSFCS5khqG6zR9+6xQraOolamonco8pEhL8D5McTtzTE6wLRs8+W5NmrewHk4xNiQzkoH6S
nOA9WykWC9D7j9ULWMIelYHB2I/n57OQYAkOpNlDm28V3r3g1crRo1XnLP4F6Gj99wnwwPc5ZOmU
Qp1cMb2qPRQiM3Ef5w/prEQH064d/+V6FoMDzhjevNscBJf9/eXf1+FtQdHZpyeBSV4QTpM8RAPu
H5r7m1jefEo+fHahMV3sfL+frus+ngLGwFpkihFtrUYq3zL50i/RAcvhx5/eTRvwdmiVURV191QW
sLAEP/bBQB0vRAYW+7UmJ9k9m8TRQuD8va8tuJYM3+mrPDpJ/WaM2wTuJCAQGvugJLAfeGWJFQKo
Zk/Gwl2Xej95YpClE2AxhYtWavOyskaYTg6Ic9i26XxJE6sXR186v28ihgXIUq8isOJjrstVxc+c
dM0k8YyWpN/6CgJ6ZaPbJTTKZK5yOjF6b2jhBjpHyCOpFHSDiSoklmoo0IwA6K6FwAGtXH4noy6w
SxNSjeH4W72g4MTYyVVO1wTf4fWYd9U4G/j38RtCFHjwBYWsAJJ3VHkYDQP1FiS4H/yVctjE7a7z
1Loth2V38iOTvThMX7qETcYHlv1FIP8VPJl2KTQuI5EeWjDUIz1rLuO1y6EIRPfTDipb/kaOinqQ
IfbQTOtT/ncgNgPVMSfUuB4xfG0uQXVWgnNFuIbvIzIBAt+1Gr1rFgPRsOY8DA49nf5WFxtl0HWw
KoBvJjHRIhYdCkZ+hoRGA/xcQhhmYlK00qChxNzmnDRv5tvbb4JUZKcgNZ6ApQPKMxZ/0Z/I5hF0
O6OLGkbGYgLDxlCLo3DDzqiBU+Q6FJkB8DYkWJqWxZjFcLah2tueZtkBgu5Ck1eF0LkfOFY7GBcS
nIccKIFN5zWGzb36Na+7JNDRfqVNIF0o6Hzbh7BZvfAaxeFRhPQzVbfB5tWM6+dRv0Fx38V3//KV
I6GK9JOuqt1ArpGLlXRj//O3kgI6fJNBTq3OpXwRzMIBfU4+16CaV1vebB800b1Fd/c9TPsvs5Zo
r0Rn43Oy6bj1I3gYhnMcpcB9e7C8C/7Lgkiqem7QeS7fl2oRjJh1wY2L+z/vJ1UB/xqmQ9JtOPEi
2MdvtSKRqmU7dvOJPBC4tiDwXuTTIJivmXRnPEBPzgoeNJObhhNE9XFT2px3Xqd0fNl2bebBgi6/
qBr5E7BwUAI2YFoq486940/JGFBNbvvjmkHQZZKqbO1qaf6jVCCDJWKKYD8wpEYdqsSvrjQFDqbB
nQ8Y4lWrOo8xN+X4sJSpgEi7TomcPyTvbKlLeTLoo4TN8XMZ834oyCKjnuAQYOYs/h4AGZhAimgp
MKFdwsjDim/CrWsv5R02WkFbVeLZUfJdsJKhhIsjTqDZagu/5Gx59SoIDTV/IaWjoLXh9uR68Tzy
TOUpi2RherZEeoYbO4uYctdE/aDxMALRBtudVTfrx/B4bE20adGthv/bnLNOgvjmFLNR+4zK+IXK
RZG2Gwu4bLuNwQUvdz/In6cBlAmnV1yn47LWjOSTAYjiALBAwD77BfBwc7GpZgyTjdEAOMpt6gLY
bWytQBgkt7KJR6pjsYY3/cgKkz3/MfvHwkpHeuLOQPgQtdXtjebCEoN8so+xa3YJbNshkArmua/D
N2yhzL3/iyBGfKxFAIIOhy0+ON56TPFvD5D1R0HaWtgeRqXYNwpDv2zDlKe8GT0be6o1gm6FmbLP
bUmcVJN8ryMl6VkKe2EKHkzAjUsSa/xyXybZ6dX823fyEbQaMFbHayxbV7wjKeBEGQmF61ZjLdiE
LfxBdE/qvmYT2aAG1rL244WNgjybaCGgP2fm8Q8iEspjorPtAfwgXtH5T7pArFQ/7d3JiiGrrEuM
NZpZ3Pp9U0Oz2yTflzW9dNupYOVQBCbI6CR9qUSVPeUC2ZKNNit3Fnm9MbUH9G9O2shRdlVWT5XU
Kzcelgm0nbT0ZLKbjZgTQIxboLFRYSE/qBKggKfnLueAL9IEdmvPxGx+UzpEbwoDpoNU/SrLc/f2
Zv4izLHtaG2iRIkyB7q1HAT0aACi6a8b86HQpdXk06/qe47Q1dCOTDJhOVkwl4n479FO9unRfgjF
CmNT2mhOXq31+0k1ex8cQdYVCrOy2Z4eAFstOjP4Z+oUFZFaS5QAG37e8yo27z3gennMKOUkeY9M
PYEquvVMRw8APPPySpDeeiytb8ZSbsXJ/6NKXfQql+jcqxWd469OUyAvk7dIHR58fC1ulj/Bn8Sa
Low5WS3p8iStDiAnAEJlGadea+Hnk/lRVwIf1b+voSD4yKmuZnc2diTQGZKSixq3UmY11yUmvQd+
6CaC3/PIXwYKGGSpxbap939MrAc7ywzS+U26XhgHUQKqb81VGwVeb/oLIueO0SuC816dBFLKptT7
FGUKxJjvfr8mQ2tzJEMopLBls/eyghHtkgOOCciFJafBuLFVlL8Er24JNwJbOvHGfISofShkKFjo
yExRXfPwRjBUiaulCqMBdIORtEaHiqEgL4P/39+g9d5S/2ZGmFrABqp4j3oCwQEPFUv4/uA3IQhI
a5pvSBk3IXmpOlBvKnN3vUMesBB3nehBxUzV4LmfiJZbkCGiRPAQHvAM9brCcefIX9CWjydl4BSw
my5iJan3Kwb+KXRxphB5rMJId/cMijTJ9Fk0x5qUctsEEeAIA1JVPG0XfTt0+ip/zxfkx1zNUhO1
exQCH8zcThZjqGRy+/3gWaFx2Ak5V5KfApKH1GoSRopEC90vUq97D+fLfSip0jP+7lEmuIOxiaAe
Um7jea5HblSBKuY8Bt3eTjBG8adn95wSW38tqbWEYnchh5Shwyrqll27MwtUTjYTWLPfxM/7PyLU
LzKqw5TjBk6Q79UBZ8UrhG/1GoGZ5zpNBK7ziB/q3QWquKGkEmxFcGh3RXjQjl+U30kI5k6Pvubj
akWWyh4qlSvWM56/fnaeonqNhuF1SK5dz1AWl5mrMTDNnk75KaAZOHaSUcfn6xXDc1GoyvGKwybh
TcU6LVpY6Gi98GyxbbLSrXa50zcA5AOto/kS2qIeZ3S8J96HWd5RPd1kq6d1mgyczN278xxMHa/f
IqkMhGyT0LyUy51R9SRbJ0gItzxfyGy6+DgMWQrM79CVnkFEpMWA43qnBGLkQ7pbfFsmj39lxh3X
Dqk2b0CAPykoOickd3XjEpl3APsr3m/pMkYsOAufMbvr0ANoknZZubTBKlLrzGWg5MpI5gnvtQiW
dRlN3+dbCcsuDF2b6aoaP66h8AIYtjwC9MQ0Q5zooxldFjhjl7tYqBQAha6mZJbvklLReopa6GCG
91kHOl60nxME6BNVid/MOwh2++GBUBzDFtYqW6giAT+xMmrpCqlIJTRbRyGfRR4ZzUqIxWx/ooaN
ALfwP5jbamxo8FuLsqssLau5m8gngmZ16xxmQcsNhanu4qMVg+fWR8jIgRqhUXI9EY6P5RlCvbrQ
PnI0mO8Y4jc5Qjm745QvhlXgEjRkMUVLbWE5ioIIh5jh/TVckN7She7JCvpXZnzH03q+PAQJKlJD
xIMUpfeqRX0vN/ZaFG5NalNfNECFyHS6VvWUrYbqwRAZWP0oM5XSbsJuEUNQihXVM0XoYxNZcAX+
TyzcT2u2CrJad3JAgZXXXEzmmuSNyIfvh4dTtq5ZDtyfT2ny/xfH+FVqRV9xC5hLKb3B6b9zNqYD
nP4D2Oks1c4QhcFXytpKTR1XR8RyRPLfaXVLuLFFavSEa4tkWgZ1+cC28OP3w+t9QiObP3NuNXOn
sWtd6rU4CBSGnVhvn/f1CkFCM/M0AJsPFKNRoX2tUwWKh4G04YUlnCB19vdnrX40+w08h/8kJ3+K
fsspz+oa0/G+k/Vv5yikORqH5YzyINS+CZiX1MZ0FExNpntpMuscrXwGFPwULUH34S0x4N0nW4Wj
JdPrAtuI4U9ezlSy/3hA1eLNup3bUv/tsjCT2LNKWy27aV0F2fc9tnEgngdsbsMVLjdpvQk9udkX
g6aS9YC9M27GzaJGVlBkMG1AzTXagZRGE8ogzz9NZyCQ7uwEIfBqwh8Cb0rICfJ93f6MEfVuwkYY
ILP0XqnnxA8QiEWun3pyzfl/VfNCih+6rdRzWlp70LNUnF39eQhzqdHhm1YwUQN7/ium5QwV31so
KPvD4MAO2c5ToyXKqKWuK9r/nryYECXQGR2LaUhrdStfi82dVoP9UKSSdw0e6Z3UTiLeLTTm7GrO
JG9giXCwVGGC2rknwXc0IvGR83uqjfVQJOHuMBPSDyWjWZshXUV5L3GLitrNAteEnPnWan3TgpFw
ZKPUD49jqojF9NHl+Y+ycBGPYh+OM7nkTYzI7a167Z9ioTDJ0LF1mpPGZ/PNO9eYLiGVROB5pugp
xahUoo15KwpeBjEjek4TxughbfpZQOftIap57XiYBsLRKIikM6vWP/waH26jaEHaJxB1G/rpr+p/
sKhsZm5EmlgXc67waXYYtj2mHAHx1YpKUus60VmlQE7pbk4F7GB5NhXMexJ+N3sWQsTQmc7+f/rY
mQXqg6vGndJpOOsVU2Vs1GRl9Cw/UESe6oWGilOPk9F1iwp+ncSg2pUXGW6x3LEwzjmavxmCptgu
AmalvlUlHWQcqCzCJMpB0ruhHKbXsgO64XCXWay/WS+huCTlYLmVHNBZIxrkqiAMHl2grMXb3/f3
SLM2ldzz8mIRx7QO0NPboUuushtxQN7T3JkhpuMwIQOy0WyFSRi8bPsvqGwdF/XzgAEEsGARIkAR
Y2gZhglIuwvHNLwmgeLpjZQiP6KaEFMhal625bGb23r0Lp5Y3Uf+TwDerePr2kBU/b7LNyvuc3FL
cl6GBTcEcITgSoe3zarrQ7XE4se+Ooc7iQZJPGVRygIVeyF3fjf1LLLupvyyvFGgWdm1O519CpOW
5MtjDKDt0nF1jEr/z41pE8ZwKcSwB66+i4MCbKes9yJWUNTfqTT4FbP9y1WmXeKQnOMIEV+S0YjI
OL2X98r5lY+zhqPB9ko9fol624JMjX1T6165GSSodHbPbF/MvQ2AKL+Ko/Gt7buS4pCxexfEUPpg
mei4FgNu65W4GgAKubn8Mkt+blL/XQXRDWCO8+N+Zd8lEbfN+gru63qZlNSL1E1LYupmihBxy43O
1y2276uLW4wVpD6WPUnu6bFY/W1Y7xfAeBGOohFKytvXRnlLNTWifYzTmtTQ9wpyXL6CSlMpezXM
HtapKF67DSfyfoeOyMw86/a2WL8PXJ+WPxVMX+lXgD+WGTLjfmWgO4Ieu1z1pi4NvDlKmVE2HLCH
3k9iCDHQA79KtnWKk3iZ+kkl8KEGnuCT0uX/KRt85th9A42QFgi0C5UvDxQ24ovYz3YtyXgXQ+UI
++fQpqzpZz1sDvc33r7kcEQvdfKeE2FzcusUsmWFd/bS80v/+5NOYhiMq6wOlgqakmSAOrSlbsW1
tjH3PQI+ODrHUPhZ51WIWFMH3LVdRqqlEQlms3OoTWZaStx12i4h2tC+ioxLlRK2B+mviHMF4H6M
boZ0GvPEKjBDnGUoOodI4CObOY7qHOSLmZvhJvHOJf48i2YTMsNrtBs1JEyyTSKhJqhvaVq+l5Z7
TuW0SOTYit3MGy/gjc69TMaWA9F7zRpqxMOXrcDKPmYI1GCVJzkA1c1+rhbp/hUPNzfNwClJOqeg
+pE1zQ06u/fN9d9kqpKffKLrdtH1L+4ijBn6Pkf6Y9X3FwwjpgOabfBwFKvGASvsuhOGhtcV9if/
NPaae+/ELsHl2Ptk94e4kdVtHgyeHWLaOfgoxYnDf/c6B6uyUR6LtbBCem41E8agq8WpqJlt0KSu
vG04z60ffXKt9LOtHHMKJU6vE3XyOJ80GKSTD8JG8SudPwx8dnrPthrigljYacFCrVvCPYp3LLbh
+aiZwZsyrqdn87nKw17MQNQeV/DelG1mp1SyEMSLIhKOu+bhtC6xsj5KD8sV7m5WLZh3BNOBXas6
o2OwIYVWti86BNeoLu71X6mc+0UdV4LolUco6qUVq/tPM3wWKOv+uApSli/4go8QWVO+L6qbxglh
6XPcLpLH20UwvKZjP6pFg0XbiIf3UlcNfPBRhQqFkdme2xGdUULQNkQuVk734n6CDi6y2clSCH0K
m/Qai51AK/lgI04ivi9it2J5r5oo37bVQdeXtOeecLe8TNAAyblhFDfDhrUt9TcJdO8Plk/t89yJ
vZpv0CrM9qD4e6teZIeYb8dSeKz5MwJEo0iCnmnQwFC+HEVdsfuHBWXHhf7BjnPOubfez9Tj0RGs
3mQufY16oO1WhGf9nxBVYz8BKsTP4+lKJhwZyvZS+dCpkwheWsTVxF1fK4RIS6IIMVpqd/3NDLoR
btdLk4kbWthj6utNUzjnsKHkUCeh/Fe+3Y1/gPbY1X8iOo+qGAFnqMLIM40FBFtfi7C0ykI0nvSN
zv2hwRsYiXv/L01ca3uF5lrhXq/194KKHEf7J1ls0KfQwIE1ewDsw+ouf0KwdhuO/2oepu9lOZC2
k2ONDRPlsNk82Rvd/dmpNC+kd15UHrmR2/Ra9nKlsQGuT6Jjz+9QO2cuWiHFP2DyB4Bxx9+xcaIN
LGBUsHTsuBgr0sof1UX9lDkmkjMuLcsGQwQs6i9BHVSqxt9Xtq4rv/MjsNigIXeRa+cEheUFXZXt
CWVMIKQZIJB+1CFGeR8ZkF7WCx7h/2qZRgTCnPTWiXHwS3s+TSvIGUzhhEHNDOb4P0SuQ9AUsbn4
XUXN9+Cryhdr/iS8PFsJBs0WYqerov+2PF2mTCjEF7s8XIY/F+9NzlHvy7xYyax4E4Fxj7qrMoNj
XCuIWuJr9Xct27Y7RKN7U1+b0cqh/233MnRXbkH0w5c0jzj0+N7F4HGrtcNuN7vZ5iViuaLrvCY5
QqXgjp3a/JqVE65zxNouPKuApeFh3eow/CH2hm3BKsrbdjLYLehKcOjrtBH9p9WEsZUWgbY1dIQc
fM4bNDzrHFSpgVN0Pnwu5IzdICQb7lvIzkDWOOHskr7clrNMQu72eEN6LfeSwzNoPoACZGwn9vVe
LLTCTj4q0jysR5DVGqJCtNu8AEwq5apWilst7iVsQhNOYEKgMOTit9Tvac2QbOB3E2tbZIltxpYB
95ncsfjevb5zwc/iFk7KGOX1lk8e6luChMgJ6uhnFjcpSqYIlxZ1W+mwV8AgAZ/TcmHO5KBzKREA
WJCQyzxOBi0mVzWtQSy+sBXP5N8aTLGNPbqEm/9xLgPGN/XXwnu/fI6QIknv03xUuhG27faCSLPJ
coWEYpAducSTZoFNMkbC6ByMi/DLahSqqF/c+giNPVolHOwDKXai1bGsipnD/Cq0i6j5BtRvljZt
5GOT6/CYt73QuhUpb7ytg0f8mbzfrZZmnPdt+FFZpDsNQbPmDchED7HkkkOVNhkt5kVRK0ROPk/P
mZ4pUyWRjkvpps9MEYt5sgNhS3rVKhJzL5Q9w0Dwh1jFXoOj5x5D3hJU0e1/yURD0b16DXRa8Yax
1hYtBwuV/C1u139tIjg7cCE8dWJ6iGWC2pIwBmP4tNX06dqAOpNnlzrR3VjYxE2Ir00F9fJQaUsS
RIUOwLUbvn+VKUfFGfjO7lAHCfynTtTLkdKPd74QE9mhjKnaplwycsTu2OAKB7Lqb2Ymlfu7uMxh
uXLYYEnbiCixGGEpv94LrDm+8AcgjEUhfJX2AhIdT8240gMuvkrGKjwYZrZuBlrcCIjp46dwjkEo
X1YjGsfKfT+PHT00x6Gv8oKcgwkiNlBH0KfJoWR6cJ2MSYGjOt5Ca+96a8hywpWfEwvkHwUYEsfl
xaACot9bhzsceItYt61EzjoJuRegBaShUJS6WRanlKwcdKCQMIr/HSupIfHiMHPQQn+lErud5k1L
B0IDL8L9BP+MAflf6mpG4iLBbGxV/LUIiHp58PxP4OwQqkDYOK7C3EjeY32oo75fsnefcsBxEalj
ssRrLLVgpWdLRLE2InKG9vMhPZp6nMibLXeHcBsgS/3uG8Wq/BZt7xFskRrGMy/XJ9uWwg87FwCk
YNDYCJTInyke1IFo2JmEscLDNHfKoJ3q2L4yZP+qMjLWl1zW1xOpEYsS1BdB7Zv3TqTEk1vrLo7v
1h7o7EMw4uAed/sOCSkYaxVkVsPEvXkgf5vJcMLiZ6esgn24nSul+o4Er4qxn3gtye0GmPXlaKpv
K8O4+c2MpAZv9QRIVX3L+3V9XodXxQWts83oOOZIZJeBB7vI9TvqRCzcKqLmmLwwrHI0r8EjivGC
97nNwQDNqiJnTM3O/ap1AYSVYB5b2a4yH9X5bKUvIBux7hkrycx++kddeGmn1ZnWavlin83eX5Um
HxZn9BXZhsyGhqqNaHskxlWpVTdwLkD/+7tGadQtcQJvYg/HwI43/8b097bPNi2Jr8PRpfp1tPqq
4U/6GbWAgU7fQF46XYBWLkbWlnR7gCknmBfhkaxh1pz9pVwr0nhDW7P7j99P9EirVvxGO8rWzzIo
PYmk/SJCkamBloTARsxcDDLQOM48nM8O+WcYlSHjpLDOvT4N3JF381aX4XrZ955b9s0MKR6nehAb
fa7qv1AHmS9AMcSou26pEj9Mj68VAR5pEJH20fy8f414TNe6HNAIDusInDUnJ0DDK2LKj+PFi+IA
yqoZis+Ews6l+dpIEZKrvn6hDYNdkPglpluy5R8bo4vpbTeEWpcrEXG5CQ+w3HQvIZFBv1G9bhqW
k8W/NowNbJqRj7QFhXOd62tOwS720G0AdgB6X/dJ3Mye0oXAMcDqiQXRURtUGC04F1SMYoMxWOcC
KZbfidb1t5BrnGuvCmcFvv805QjWGfkwMxiOWnPZgUTcy7I80Oqpb09LY7I8Sn5h26r+XYlqEgQS
UiijMPtovAam2J4HQV1vQg3hK4foxPi1+l+a1OwBxXUwcmMPecsWwB6h4BcsiP+ZS3U6u/aMzO9I
C8H3ocnrqeZIAzMtiSot9WdQJDlhT2sA04A2cGh5fi3jNkHki+iK+aKG3X1yMKQgR6kF9C40KycR
kaim89P2wdngeUo8e8Et3TGsg+SHmVZZ0eyLi/TFEX4osXAVPKpYxwHJZR7DHQWMzW+xHRVnkkWN
tC/jJJCSs2bCV/5xcp98uU2MOxdlKuxI1Ro5ZWl0JOnlZkxuD5KZe7lDpJyoufXzh4F0Z4sF1aPe
zaL8xB0ectq/RlxEbFcrG9wKt9Tc11zciC3X16ioo5QJDfOJwfuAOOSh+V+cch7CNnBoWaz3qYSi
x5e8h6m8gxNStrFSkGaWtPF90wFVTJ+EOlGopqRATzLKnuBuKOhMH/QhtEomciGwg9BvjDPTiIu2
Sobsu54lYz6avK2sUxW/ZM+sG8gjtNfJIRWH+u1bAo//AEu8rstSvFGxH0cvgdJRGo4PtJnGZY7v
BolJ92N8iZsvb97P5JRDMdDO+Dj9hzvxpe/252Tqod6bD+6EwOMjt+X8xeINQu+jiF531yihQw4g
ts0Lg8W0ErPGbgqdQX9G6e1TadTqtWpAuZ4WtbYm1Rclzx8B9OAmp039wR7XUYxQ+oFppmjQxUKA
Odf7R2tnQw+hPuGsk5qHAPJc3uIk10anTnHrfSRRef05v2PPuPFf7W7HWVgV68xz5PhuJUI0SVZ0
V/Y5fbDy9SW57yOyiuu7boUaTlavWKJarZZHSSNtnAqWni0OmyR0L+N1seC+RkOCFwYMw8D+Ak/V
6pqz5y0+kKy9tqQ1ykaCl5kn7+hfRlHwXgpZipaS5hBZqP89nspvJOQKS47KD1jUFiWYA3YG0Y2R
L1lDrJPyKQQ/oKLNEpTyRkyKgx/48fYxg3c9lilmDGchzc/4g+R8XMRZIs3nco9ZwqGZJXyR5ceg
w5u9D1Etn2INCx9X3cHXwtXheAIj28rtuxA+DZ9gZ0VbYD/Ws/WwDSZ1RAl5So/Ay/vpttjYc1Ss
yGwWvbvDEqyOBBLEOXdcunms22hpHlQWvyZuyvo/coAEmimqErXzJXeQXYAMFUGcB1sizfJJJlfQ
mWcFWuw1aKS6xt/ncnwdS1/98go8Zc8At5UXevKjCfgDVjSFBre2bBqnWaw1WJ8VtPazLF8zJ3SA
U+ANr4LjoJP6K4SUw9Wq7Xe40c7s3DSRG3zMpyjuQtKzhI8qGFJFFewxepimhLshtV84sfWVACmU
ACU+BbFomyGHgji7SumtKWl+HpBJITzG1hUYLT9gc1Ow4sUJ60ijfEcNTP8auViiSV45dVQq1E2C
QwDIE6IPi2ms8gp1PkYepsNm0+R3rjJ+ex2Gc8GJrutGNe+v3oXNNKASxD4H1RzfOdqU6eScxHdA
9g8RWrAAW3+xjR5qpFYqIjvwH8g0SNMeOJI+4d7FkpqgWBNf9AM2GO4b+dKjxypudUPpO7eSqvZL
3oSqpY9jQeT4MCVqAkwE6p52zvZY7Vke24/hgxgirNk0JTCUGFMjKQYxiRzKeziLu+Ddz15a2Y2B
uRQ0xz6gwtcd9ZM+MGL2JAqNVKI2XidXWVmr8eB/FkDbth9i9Z0uy+xAx9iiS357r3GSLM69arTP
S8w8eiG+7zZifAmVg/qpYW6C7zrDrcJPw82afaukf6/GdGdiBCufXOCp666VoSX/tdl3H7rcd7Lr
bjgakTmlae7rtjKmm80U5MFSCcijJcdL+HpbuFH7L0U6FTto0ey01aMncgspE+a16q8JyrqeuPD4
bgHfFgjn/29zQyeolRhP3L7LsRXSJzodCn4k/PJ8oFixdhi+oB3lcsEVbeGbCYjCPJ/6FnJRVck/
uo0nRrMtDaT5uCTHUebO9coltoJOwCsMdYoL8UoVW4xlS5tQtVYN7/dKFLKmrAPn3sU0RF7i4lsn
DTt+7VV4zzXuYsm7OQdA8538UYAXy7JpoxkGJ4PTgwRCBqXFNnlvsOdzQV3eUYEZeczdubXYGeQi
NKAzSDK1x22r+mQqF3GO4p3wLBo2efOvbRFgmDLHOYIiHOl7R7NIyAGSYrGJr6czKsHs1g1ViR4A
BbI6jxKMvuWgpaefLLxKtiM8zT9hZl61+HFxzXTS1fOdkC4ms7EAkwuaYTlNpP7w530nUqUx6vur
umxcUnwYMRkXgV/jQAJoRQu9rGmoHmRlu8Xv6/6kVquBleHW0QjH7Xme/r872PfHdw8ZxMTkaj99
13IM62yLZ/5+rhyhAgoFPrdFZXTlxG/L/3JfilT7lRO0ltIJfT227eOGBbUrxTco0Zx+9W6/0oD2
Mcw26uksxpwNCcsW1HZ4jQ91cnL487JNfm7KXMryKLz67gnBjA6CEcZJsFnMOOyDTmJ6E9TS4CJq
HrpXRWiBFoyPpU5Y/Eu7oirqDMg6UGYeOWOTZIu4ndB1gPGxObID3Ri+sCc2iR0eSe3/rLWELgaQ
xz+tiSNN5PhR9x5rxM7EQ+xzWDgSfHpwvC7ezdTb3CM2KKtLAtr1YbBmGDAPX8HQ76Cs//a7zl0h
XtqK6rNiFSB7aBykXBXy7Iz3gU96sQaJqy0x2Hn2kgB02nC6SBPXORG6djojlO8zITL4Q5pep5DS
1Myn7jg1z54Wyxtp8HdPdJby0r+vfqyV9V+YtuT3l65YcVDSWeho9woNKZTZYERHtD0rU1HANk5x
qBhliV4RA0hCg3LftE8FigNvrzpp3gIOWyeBgAGvPUWgtOe69N/je7v3yYfXAuegYjWvfJHPS4Ks
TyZJLakepVM2XwozsjvrBGsiEoWPYOSn1NmXrODvYIKispPOTPICl6uOo77H4crducna2oZS8fQ7
TgigKjWTmRhb/On/FWb0UnqBF5oSDDy+kidLL0QlnEzrFIqRsTS3C4T/ZyjVvhcZfmJl0srQ86oV
If9Vkxr1F2IUXzdxOHKXr3OF0h5oX2YMrWT0hDAbC4tVRxTt12wMOQSiBSD3K6hfepmS7+6eB1A8
72Ijzz3CzcMbpQQhUwVRHBwocfVKQmwbr194NowenCpF6a11rB5UT7QCWwDIEo3zv7wg2PWttUJS
WJQkXNHerkXTOPHPCbuVSIbL2MVFicC0gNJ/a5eRkTQeHIAPxee439dnv/gumIENxLXbysryT/wC
IUjmb2+reeiMkQ1wdD12n/UyAmWOUdHhRblqdrwOj111qK3B9JFltU97pJQm+cEWCEUSbVgqp268
hP76HfV1IVxWkFV3OMUSN7Cm8kq49mAfzQ37EzP6K0xN0r4G56dVtYtaBpSCNaQQaoCtSqgSaoJv
/nZID9zb9BZBYUc5WHgMGi7GSu1ZKnIrRHOZYAQnDFL2FNUQuVjzICWecCobF0sbmEMRkaZ6xDfM
lRTYQxk6Y0zoMZu6bzS/vjrbCmrV677FqSkeel14aAt9J7DhrxVVpe43SKlv+/upxXHyTPNKcpe7
cqcBWCv1UAOL47gNAIC+GITd5z6qz90fRp1vFlK/Ch7nlNmo/L+zVps0Vooa2gW1Q9GxvELGpnOS
hiifqASBLw7bqzZy0zkTAmqNYVB2Ma3Rw/MbcSw2sVaXmTaEyAtd3xRxEIvjborduGkTUT4r0N2l
GGHhIXSVYOIME+TxwFBWzo1uYJWyzkNm0iwfK0E6eIRzUukU0GblA+rTpwwG85TZA8kOp3nCKsj2
MG3+kMnfHKzai1i7SM4Suf/Mr3ObkXTqnrkLPBE3KEJCBshgr8pP8wtS3DXltawTYYHyJ2sZCvtG
J/0Jy/h9zMg9cLmGxEeDSpZm64AFya995D93eOGcB4Mgg5L5wc3icqdAoAkr8R9Cy1zedZGMkSxX
bwrOlfO0sLeJpcT2XVIbfNvmpHSWFmqF9f+nnzZ/bhytca/+NCbnimQkkBuwgtr0eNi0EFM4pHOx
19SVG8DGOs316rl6PhudRQPoTzRP20ofcw77n6wMJCNbB+Y5Ty05gq23YULhVp0hNOXqwNUPxRo9
IzddJt7bXdlHA+lkqXm6QQGrQd8pQsrabi0kMnXHPvc6wa7JbS656mhzYlz1q0EdBrSCHm5ZjmGM
TBY8Vjp6gg1RKBUoCFAiiiXCUHxB2l7yKA564SvITniC6PPrhIWJNIp1JHE93ozSvMIP2fHNdWci
U+uqxthnMAJ3SJbDRY1mbiHBizJGIoaB+iQQg0GzK4w6pg33GInT93jOVgT6ygBBY6BjiDDV/3Hp
DOU7EYZSZouPCC7Rwoo8jcj4C0aLrEiCJqURXjSUggol4+co/fWuCFBTvwDQ2nSppzhGmxot26qn
K4BE+SfURsLSDZvCz+JcIT1un3TCHBfHrQ/rTUjLWIO+8j9iQQoc2Fwe3BZ4qgilh3kUVQbmMCWM
eG/8j5UqxzjolYPNqAEKXo49Cvj9OjL7hmFnrrZFgKzk3BETLNAU99Bm5Vg/0D10aFqJrer1Jsf/
rn5LC9jyLq6VGPYjeTZzdDCAMXUuAdVsyi7YmcRwNw6Chg5L2HK3ZER1zCqw0O/ZnRMhLHqRjaXh
34nBwWhHMFMnjIifspBfLGz7z9I7fgFixwE+iSWrXBq/+vk7JBZvElzNfJ7HjUP/AvwA29d9o9xj
huKnays9RObfLUPfTeBRWi/7FCYDpZ37g+l4Cbs/TC4F6KAvWcofvBtpvUdiVwrlDU9bu13h60ni
1t0jjPUrXb0VfwsFSYG7Rv3NA5oauG5iawyyQ7U4128cqCpSOkeCZQ7jgg/FhCHQR5LCd2gyS/rh
sSua0l5bISaj/y/2Q8kA5Kfa9pn9hFHQrSwYn3V9KnSCwU6lox35X2kzEP5Iq1V9xI1OvWKpOdT1
Qn6FoijTTMDJE2Iaontgib+FWuS9F7yUe0T2JBJj/2rRJz3waQ+61b3Q6uKWnv+9VzHa79hXy46g
Xasfa2uV9Y1nonv1YAAm4D50z6TulxQ6/rYZFqRFWDbF7QqyW8Vny0QT1Cfb67tisQ7b9N1+/G4D
E8m3u8LxEy2ppI176SyneepkRGtPL+Qkmb7Sw2S/28CyijW245pxtnLXKirb3K1HcZcUIk2RWGGl
xs4z+Tw0s8LosFcGJgfYy+xgjsD0C0K0apaAdDpcQnspYG99UE5Pqq2HmhIzvFFIjjtN7thtKnZ9
JgpQrf/PhaZouSD8kQvo2kNdTF6SHgJb0l9Df0U5SbCKKoKg+KYKXrfTVagtvut2CF4/K075q3df
ChjOoWhpF3OUeJb/BUIv4faVIHyN3fLIq6GniO0y/QLSPKAB8upfAZ7dxrcdy1TTThzw0I9K1FJh
38++0tE98zaOwXBRtXY8KRprydaFO5AaXOIyLFAqWcoqFGRWJzN7zlYYkL/YVuICjaf/nJ0/e6w6
zKkdVkGi+U4K6JiTMPviPHzhtCpxuEZmWxrcH7liQ1a0FyrIndiRYJVVbMznwWRhbpjZguCZuakP
mcQo6qaJIHbs3bWtyVqC2ZdyqJs48qGJ1EUtEblIiFO539t1aWsec0QElDtWxptvn7mzKq7OF22z
xurL8FMV5bqZVA+rljFxQLfxBZsl4KxlLoE0qfOmnEJ7QJBIDSoHECd7G+Wa0LMZtDD1GxKvKuFw
Nit2Ednbi5o5bUEDB2uFAYfHTP8x+fCA3mIUx3fmqLemwWBHix0B2mifv1bjxEwVk+Zq5mhFXAo4
/LHqelkufcR9JMVl6CYXn3G910C3d37ZRgKMJE2Q1AKWW9Zxtp8I8n7X0mKC1btlgUGbTGoY4hOG
8TB4yuQIMLEA0V79hPPkrH/of+rny02DZh0XHX8jC9JVpt4027ygBL/pXZ6v8vAFE398s7m3sJq1
7yQzXY8fMNyyOlN1ObDZpo5AldHI4Zm4DWhq/nqYcCWEB+9v3Ei8QP/XuLz4Oyd7E99YC7NCcw1w
CTDaWTjQ1HHTRl25/RWgaGECEc3k8k3nrZyBe8yRu1XAGESNGOMDD6/qEVAa9xOoMPjtq9a8yHTC
XUEakoHIgfY1speiP5L7TZv+eEyTqUTzoO2Mi4kfmkAQC57NWEBwRCJTBrJ9p/XcnT/eDnyMYkJF
Njm+6bnwBlXk36JPA+l3zlDi+46VtvfvV84gu8DBu9bIi66IEh/tifLaKj4EFSMGL5lm1gwhssvb
7onJCc1ZlAfkiUCU3bKgxlsV+za9YeyJjIssoxx0RI2GCOWCcsOBoO2/JBoPAKbXdlkjpGHPQEKX
sc8cumw4yRnJQ5UZrTqHl7j5MXTEORCZu3nP6+rvfti0rYRFkZqT1vaBQ96/q5RYmXkq7f1MYmUV
WgufM9BJdTuRee6eaq7TfhRvYDkkqfhlSKAL7XsL+Hp6apSYIYl8BAxMl55La/56sbj35qvVPgGU
/J3CPRD3buGROr629gW2ZQagu/U1JiYcqBKRuOHFJ20FScb/mefiTUqF/AMeTBf5BGkzRMKX7DCP
/lrmzVMvloPZGV5g66fBmCnmw/e0+7/bF5zV8GGHmHXS7FtfSBkIrK2hD1eXqiZhXGDxQKeFoRDP
w5CRSJqDEp42HvfiD55Xp0CwHgTxmp7wJazeoIGzjIrzGOypcEzMfawXsV9e8sC6xVaa5GJc5dw1
m5CAsVt6IZR0bMTUYLw0v2VlIrFtkgycrzFq4eitLf5fH4wC5/VnFRKtDx6kMsS8ABtqpMJZEddA
dPrhL/lIZvuuhyQVB2rD67uDaQSP/eO0CWwnptl04GpQysmUWiw5+aYtUUfUHd3znOEnt+dAJWwi
Yd8Yb7bnUW4xGq54GfUZgSrVMrqikOdMnsXR0+ksE6g7mZ0txNXGJxH8t2C6msGZUOabFeIVaQjA
BrffniHSDXVvEp+CFHRBLfY7XkqsO/DA8rrSXtvpqjyfK88mLXqtzI4ijk8OD1Wxb1d19eir4w2z
dbYin/srdG/HazAtCZ/p7ydmBTXSpjSnVNQ+bTZAMVK7HGh4jtXzudC+MXqXvi80GwzVuFLWOCoN
gSl4RkTsgD1Y/H5j8RPEje/Worow3OMr8bDbG/rw9QKZAVf0fmbQ71eAqfB+9njVQnOLYePKWZHK
btcP02voARZNfEaHmz3ls2l28Krs6zF58LF6rqiVyuiAW11LiZSLZpDZ54YMlK5l+Qg51Pt0KDNS
9q0A9AZcH+/qXVOheMh1A7yHlYt3KjijODajlRHyIwoIwVbUvlVmjN6A1IXOXdn4g15GNL5be392
xo2m5oua/Jf8vemib3dnKKqnmnMNHMtHs2QShnIIzGl6cp0dnZA/3yM0CvJiXm7Hi+x1nM3w1oJB
bD5Zah43e3wB2C1ejIYVANYIpnFmL3YT6lDDVD7mw/dgShGDtE6YRcp3DqLBAV/Utc80KUGmKDuO
ZYAqoqiBjnW775dm2+JFSKO9aae4tDFkC16HZtbKbFm31lRf/51jGyHAQcJckLhFZ/FAjcldDR7/
+CCyH/hiqqIphYQaYw5PKy6/0faKGhKG2aZlZXlsmR0vDTwC0GBEI4iAuBr0i8E9rpMwoDlPeCtc
yjix2EGxe0SbI75STtecG09YiBsGuLtjSZPzlY0071etm8tBRxscUTSqt8bD56Kpf8+KfQs0dyYE
CaJ6i1uL/DKNHj1NfyaKj5ZTih7M8e9SSl65dRujSZCz/flrsN60AcH8HjyHmqepVFiBABX60sG7
33S0wOEDeDWqRXqKqel+AqnTsOdoe7jlqtHkVe2cv4bcVHVmlLp4CTd4DJhCPgJ4jOWeJFj0ocu/
wk1qHjxUQ2D+fVjKMRDv7cEEcG9lWZamySYVpTaA+5dxNWya4PxOMZh9xMuVp/CB6VFAl96rMsQz
O1xZgPuApdF1pyPMb05F7q3eCXlwMYQbGGKVQ2FF4pNiycQEYVUj/8TuuBZ6bDyYwWESP9GV7nmg
aT+oeiODOeqoycAjyGPUST40D7JWlFyFbeiMtcLfzYvHtSVecvve3ltjR7MuzkqV4x0uairs+kwT
w4DDMsEKi6VJPx/VDL10UIhIyJR+W8lVqTYm9XDrOJBnvfZzPArlNxos+5SRRXwJVC8C3PY89C/4
ZbxysDXeO4ILuBiXkR1i4t0tucWzu3h+QOjSFgzplVpA8kwtP76tXNyKvOuCMMg9i7u9hVodsa0m
30rVfMMr9DsR+WQxZdh4/b2qZ8O1h0MQOuXg6XevH9434ZU+heX/S4WlnpVLSAYa8E7T/o/vuv+b
RTKEBqBFGF5d4gFS+mEyg9kVt2BqdGEJmL31Og4Eosgn4klK8bLj6tVRCFS0ALhELoM6AXW6HH8f
t4S9NZRGWnZqEHumVqclQpOyJstcs5KSQQFgmoY3sGIHTGPy/fFFUadddZyTR/l4GhDPeLjp/V6K
a94zJGlG2jP3lhZM2TmI9gWmlPj9Q8GEtHjqI1jAa2ss5pRyJtzRJpM6RFu33/qNPe57WzcnUPoe
9L8IKFActxEs6WIj4YE43NQHzlzCfY6QocIJPPAhj0/KY+OsLoONKp/UdLSexpC2Ct51aqisuOV6
FpE1i8g1SnYYkaSbe12/Lbv4sx6IJBuFR4Nw7PfheglT/P+uHbPScU8AP6/ORbJT7SpguNjUr+q2
08aOYyYoZxijtnYsUmlyDlKPUfvxvsTL17DaFyRWwPfG7Y8hc0BcjvGzwhkXCp/iqyZtl6g7cy0S
n3SKvEyEM9GjNQ2N6k9rXT4vbyUjNfAUbl5kG9d5P28KJyGJ/gjzHs6pd3j7yC1q9qN3VQS6X5Mj
1DwuW76ynKpOxtkQFcrH1mSDgxlK9yQPT3Po9t2uBwDjlpzvoCCgHCqwkhwuZ6xR6KRz9ccJhIep
D80QOerHDJVJafcBlONuewESk1o4S0255PXsav35dXCRFql4LeQos+mP5OxLD9V6EHXLRiCfbX0a
Xr2lnmUw6w9SDakWweRshOI6K5JWxQnOA8G5galMObUwpjemj6rbbg3VQ4F9lkM1M+LqojibugEn
bjjDKYQ/CU3MKeuQyS+m1UuBOhi14UTcL666xVM8eaZDTmT3ErPt5r2Z36Tgrj/odBo7HwOz4g+v
MyZeJ3hv0UvB9k0TBPpAzUpBzIjuB/4NLS2iPcm2YWnKhxHKNxbsj0+Do14O02yLlMURqY+QOK4v
vjUOh6RG0rAUN9VgWAkj8yPXStih4OW0rgTNQctlhTnnXp1aM2bjxuva7nE+PmVXm8SH4AE6YmjW
awmZijqO19VvJ7MyI4hddP+wMu5tnTDBmYXVqR1wpWv8CdzBsrcXLpb/ka+9Sy+txLm8X9v9depo
U2xmrjSrSRnONRCSSLqft1oA4D13RboeGNo24SSZaTh2s7NSo2DogrevUcUALjdIcYc6RF105nGd
0KReMEz7s3ahNo4gZM7UWdVg2T24iHwDzONAnW+xoDLLf/rCIvg8vfcMGtaZ4/AXwbTifSY/vbAq
zgaC+/F54f2XwnrtDL1xcJa3o8XWJqyLsVreLXcvVrF/8IWvOH5qp2UMPmD5+QqsW+trPOHF4Oh6
N5Cd8Ya7nqNLSFJ0G6O9OoAMHmvbokvNGMXHItYXgdGRz9xblBTrKr59Bi1BET0aMNvc/o5UvZGo
4aGN7nJXQ4PbRIjTmxUcGJPe1PJkvLMiScnlebaGjxvq9oeX8aZaph4S9H/tmr7GlsNr6sCmRK46
ygaOAJDitLxLuEG04zn0XaT6/f0zlW7l77Vnzhz5XvoU7tEiMlObEfwes3JH30aZErRuQxshNkyw
0KgPRT5FAuazBQk7p63uY2Z08z8kZCTiZfZxEQ+SVYrXn41ylCXjH6csJsM+0y3EokhtIDCB8Hhr
TCPcdvG+JIs4uTCBKcPnyrx3ZJ6LW+gh+jUifZzUE8pw4F0UlC0RO9zMQZMO/9AYBxL3jMpXXvIB
8Qk3L8cpIR4JmxNjq2jhqytPY1rTD3voeIXft/yoH0pTYb48sYZb9Ciy3RMWhq13SbT7Q69FdHRQ
jPhNwxAyj6CRhMi837GFkfaRFyk8zmRZwx5RCzUhay1mX6aajEW7Uq8zS7IVVVOM6wQ6V8nP9FUb
vCNOXRMbjjaw3+YEjryYwKTBG96G4UvG9CMaIaE9iw+g+VWBvx2vVlxZZXQHJBTTuHTrS7xZ/nAN
7H/4q7jK8Fiso4dNuYWzTK5yShaDpSoKUkuEWV+X1t24rLCaPxWMfOpa80inf5QneYRqJcSjpv7W
nAfwTy5l6aDa2pNG5XrZLpUPFoz4OUrddYTFqmClvsemHbi+WKFDnFybfdI6+9IiolGUMnaa+ZTF
zGriovQdhIWnEE2D+71/R00mFSL6TJYq++Fsx6n2QShSFkW7O1f6HLKQ7n/LN+0/uQWh0olYXhTm
a3/XRUtPrUiTYBpvoFeXDQUrIiX5aeDrllEVx8oUFbk7zXGQftTEoUY1LwBghsQGvP0v80kK5Sq/
r44kIrxFVLexnKpv0rgQu/ggduW9XqHne4jjAnXfiGHVrunXLyv/k81SqDWAqNSIujLziswrKWe2
Esque8DRlMDg8ZSYo/Ragn+vmZbCNobtstgy7bUrAR++ZJdQouSCJvoe7o4u+u+I46Efx9kBxa9V
SpwXJfYedSgi+O2ZVzoaMPiYG7EfM3BJKF0E/zVHN+D5dIVWHCCRsHBu2PFMy+9Ruvp8XMckrhqc
2+/4fFYBtguMpZFc1R8s1GW7OT84enN7ds/sTF0pVjyeFirGauMNnZAqMu01qqI5iwJcMnMkgZSH
gUzNRDZaeufxMEpe6JwQ5uRdaajLroQHY3HXUTydWq93BldPuCa5ld/PdzFsL4i71qx9Nve5jCj2
qy3nkiNS0fm/rz6LJS75a+CxN68L0x/yb2Ir928lZZQ8d142kGx2fChvtexE36QFOLn6SE3UE3WW
w7Sv2sQ3TAA1mkAQcF4W41vA5mRFKC38pC/WC1UYC8NDqF3BsJyl+WVsVK93Nb+wVT/jgZclZmuw
EJY4dI6FxQ2FrYmjSyC6rDDWEzsUDyK3GH39EKP9RVuEatOCwO30HP1FfFtw0wrmnbpPvo82uHRK
nOLPbm7pcdPgACU1c73hOzQEs8ta46FuUe6BkW93nz2o2kEaJvDsm+COgZu7m+9V5vb7mG6BHifS
UvVFtopqQIRV4ut8uY1aPO6O2YVlwnhQHNqiO37+0Mv0gLmay4jP+SGAK0GIkBy72eGqeNnf0S8G
mbn3u/7r/ozNadC2iMQ2vSBeObAM82S1+zST7QVFZpit2uqdiYHJx5VlOy67C/EZHDdlylWkHgVH
Bfcq3xeaq9OY7CYwiRmFUttYjf37RH8vhHpF+6+PhQkxziEWxEJS9aQ4cDFh0Wd/+JaWx5txZ024
H7EAzZaAIy7D7rgCd6CcutnTdwUdpJGVWKvQGZX036nh583ERNvog+ihdhB+Wabu80pzlEFG+Fxo
vy4MkhG39o6MYlg8iO9nZq2BYwD3cVLd4kux4vsP9ZGuOVT3rV2Yi9nkvvDcYPkspzmRL8cOq6v/
ihkYPkkLqhB4EiEUA65UyaIWFdVmKidwCiFqmK6qgtAyCwv8m2OgYoPIVWDaoMtxuyv1PJmPn8oh
Zfyp/owbR5I/XTs1jDBiMoNY+6QEkDt5mO7WEoUY2E+MgrfAVGvqYsH0IA7t1dcwwumI3F1F1L7v
UwaSVkDHG8ab+wQHDnLxbhcEjOFngs3IZ9JRaaAWKmEpW8EWLOoiX2yn4+krkc7HaUOdeMH7Iv5w
e4ANTDspKShDo7WecZMt0AnRgaQ7ucsGtWcAgXanMa75YB9D+S1p8szbEdtdGlV5tWIjlOcbBICj
Wh6bi2VqKyeX+Pk5UBs8Ufsta3ui6gTgOesURYy8ghvCb3pHR6n3bF/SeAteU25EV2U9E8bmNaGb
txPBAcs39NE1abXx3aytFyz5VXebVOH1HblE2ymKY+kCG8MxMyRHEYzGVk6D38l7vU4942CSowFR
qoq4VPNwYpEKEL4Wx6tIb4tXXWv5b/Np0hDYabop+8xRMaXcuT2njXNiTWx5wjp+QbvZ492FZHUX
cAQ0zF4lqvdRJ71bWuktaClU/k7U0a681aZRD7PV/4fac2Q+0MNFXUim71SMZ3+9LplPDjX4uofq
KtlYqkjLSfuS8Xccpmwado+sFzG3WyUGhCuYmH2+MiJw/bp0ZwsLTMiw6GQaeDY+jPx8HTeAG1k6
G8ECOsQHU0kBBkZ/rGwtSawgFeQkkDPw1WxfsHO36uWh9zP9mVu+N5yp2UCgIkQWnsx9VkEBbidV
mH5+qhvecNajIIrcsTI4o5YNsJiXfBlWCXkeAYap9320zJ4HpSf2IajtKcMT2EpdOp+DqekcNWrk
LhoeGQGnWLH9TycjYXJsRYkm1LJcKeeEWRg+BL9GuNaZDRLXfpihhwfYZNXXQAiSw8GAnWSzaqwP
ULQJENc9gOmj8z6RWVGLGZ4nn+xz+XRi9m8uzRU1w0ZcST8XEbRQ+kWWUTZteBHC+0sH5PWhlkBv
W4zzOAfyvaYjcm+wD/Ktmq76fDl0xGbJo+hZU2O00bHv1wLQ/c2WiG7rdpt0g43ppO+vJokK1f+a
PKWmDt8/voeWdS/EYdupnq9oKMQj8a7ZjPXn/wRknOetYxGp0YK/vFDO4ijCJInOEWqiYjauaFXb
S5bTART3GrjGW1fGTVD8mR9sd/v2PdfK2NegCRpfRWLdpboioAVeysMHHYJT5xdYP0PS7OFUMctX
a7VTDxbWaFyJuJULNPE0/yBD2lRh3YY1PNfRApW2avRwLSt0zoW7AowA/O6F3sWFwV/EpnHbavPz
XVUXml/SY/lwYS20safNYDQ/aIw0ZpDbRmajCUci9ur/XaQFSHcwn3rHXywGVSPZ7KJFxLIK5T3d
b6p5WqP8v6ZJmnfS/mn2RyhmzOT8L6zq5y5VHsEEuhDHS3jKfhSj8sJFL5x4f6BQtmdTXJmb8Xx8
zPc0rCCWgh2Pz6grtDyKbevWUoc2CZ1Q1W8VH66ZgOAiiqWaTN1+R9r9p4inPXJu7wEu6Wp+mJ2K
1seUc/PvJRRQi18kfEYRhQykG81w/09vRYOHhJ4zG8Z2oDPd3aLa1NxrEkyIPm71JsRB/Xu8snlB
c7BPmCcFY3WhNCqpHoQOFg2M/ESIgsoNsM8iD/06/0Cbi2rdxmU3j56mrGaXp1q3uLQclssEducP
WAgfsxZrDtnx+iNaODelbnhiquJGD/eODGPiWTP1giZ6tsZ5Xh62j6RFVeu81kjBv2s4EnI1nvVV
kQLoDCfwS+QKhLgiBUgX2on+SEc/mksAv5Z4dFB3ZH80axCJSNa5N3oBSJfty7rIhOs2tFuG2VCd
tcY9HKEyjwKXdVuiQ3RhINjlui29zpKqWO05B1/itJwYi5tSMaqx/0XLIN/4QL2mxtBcttwYqzRo
2uIosM0xmjEKsyo8xU0PLg0HEQaG70FPI2oDvAOfNPpYCd43BI6X3aTmk5uQkya/yBoUet50uS7i
cNMp6u4AecE7cN29fIEashCmVcF1BqJ5h7tIwF5muqa2OzhJEsxqCI6tdtBvkrG8XQUURATEaN0N
97x/bSCw6gEkCjdrOwWlbB4EsIUbf1r5NU5H4IalN5UxGoabS1EU74xT6Od4DiXHLQYIi74UgshO
GTumia890XluMJBE1pN8YuQZ7y689fGzKijcirYXUdwkZ9aT7De9e7US238axxtYYkpyxGSF6y2G
haCCoqpv4vuxPg6E7hvN70s/xOk3s8ZlWzlU1s76VuSyQV+nC/0XdsHQVD1E1Ey2mTBfHdRoJ9PU
qMtFEP0K9Z/7lVwhjJ9R+a2JnSXIKpL7NALcIjOVpmo3mtAuUsgqDNJrbbE3vyp91HKSfnpZmObG
ZkPfMOtB7RYiI2XFrks3y8lCtF8oizFf3KpoT/VatiKVWuom4JEgsbFKHlBEvKklLLMUI+Jy4CZ7
H1HA12jAKQFKyHbUwzsaCyQ8W2D3g2Xf07dFD60EQMWbTpDvULupVuigLb/ssOWRvxvVwhDelpip
e6RUUHV1b5bHKvmz+Zsk8s3LLtD7LOhEkUlzW5iucsNh1gMiKE6CA5bKgftLAgHcgtAXKhzI8KRq
O7KkifLzXUJPSG7xcgpe5ooOrufyNOB51f8+RBx1wNjdpycFso/pUxQPzLlFXPXzaxbG2pYxRmhW
pUMxy/ogvFMe5AFLiuZdDtdcZ4F0EskG7FaatsFJKNTkBR+IjPrvzKjGZcdfbi5KKQwZRQyf4uCf
zz2uOkn4bm99COePxW2VoQQ4u4ZS/NcPMHTD7SkUnFeP41PXuChxkPs+boFFimLQPlKq530B1W3V
ua09E90ySM6bI2av3LHD0AYegrKkER9pRLOAc/n56VBj69KYAri8OGjtDGKz5bgk9JZ4GIH84V1t
BTSls1jBOtj+aif6lV6qIzPfmHBSU349xKrWysmTy9ecrN/NrGePVlCS/8jE7eXifwBG02TwQzQS
Xu0zY3Ue3x4T7CC/XBr0MjKh3ywDJI4latvD1JwDBHlz+lIOh+hLEYCp2ImA6sS3dXYLF5OHvhNX
6V53pFqE3OzoN+TmES5BnEQYNujQ9Kc2VNuwImC4MpJRVWUl5ojeKvItG7c5tevUYDIu9zQkvbu5
u0ipEyaf/erM9onpjO7F84WgbOk7fBEPhW6AzyB0iVTclqMH1M1ojxlmPxCKRAwtK80ibymr4WFB
XIZd5P+PHfncVM3pMUjM130gZsYd9uO2kAnpmqzEU7bDyY3TguHuY0ZUDqZe4Dbl4Xjd9Hc21rkD
SDCANJpCTSwarjyqxO/QTBcJnC8ccpGunMzNBbmKmYlWJFvC1ELb5DZc9brQwN4x7swkDUMWHk3b
OKri7Rm3JeGe4d8aoFRVQ3lCSOx3jAfBx7KlpVshF3s3QWz/F42JwlKUi1VooFz7i8o31a+p/WLx
qPvqinSOHdpHaPUrqWFU9t20+ZgfZWK+DQ9YCl7Phr5tb986JItI+40s/mHl8UMUn6zniEahBRyP
vRjyBl3StowTUxrx8eafsZr9cp+koreAK9t/XFdgV7eEjl/Y2lXrzvJuwzElXfnEjINBgh/wBgC9
355crQhU7Q3OQo3/3C0pNRsPdiG8HvaGNyudGfphuZv+MB0DGV9X4jhyPv3eBmDbVkTBXTPk42yU
qUrfXhNPCIYvGsDtdrJ6e197ITdwoIQ6DwQ53+C0sY8R5Z7rkpe3l026a6CsbrDb9i6Mn9A94LlK
BviFo0RVwKDGOaOmoAPFjjLDeOAaaWXGOgRFf6nQcs2/QZuFgjnmX4OoQ6emTWbtCEiew8YmWHUh
/e2U+Q0tPDFfemywDv0/OU6H7yl4rfyIorpMyPY+B/YgHHsSFAY+1sFOdTrWaDD7D++o6qDlo47g
VIjAO+mW2jii2GfQbWvfEXHUWcn8xMRFt8caQ6z216j4WGAUyaSSiP/XIQF/Xg7NNmNrxjAlCSMq
8oETloBPo32eAhc6nhwRtsSDafcMviJ4rXAbSKO/1v7kqeKKO+KoaduKx2chuFyHi/83xBneZG59
hy9tBPIcAmmyRMo5i3mLS1YGSTV5zxtBIjiCbg/pjufXslqaPvB5jr1wBKSBl+dns0eFlUn9PuHj
OonGePFZlkAC8CJdOseEFH/pmUvQXPE3IwtNoZqU/KJDIThm9YL7ATYy+wG4TveSClBl/Cuw8Loe
jNizERFDs9CMopsSJFq+iu1dvS/+uFOlQjJgCGrx3o4MztGu/AWNrFJT4HaOVbKWXBM2BJKx6PkS
SrawWcb1mJvKSOFvtuiXimY5UI52cyrIhAA4zzsJQ3N8eWC6RBzVETt+nvGVk7qwb1loNyzPSJdd
e2Qy5PS45jEA+tSpyiBUOOxsHBVKho3Na1+PFm8J4w1Qg+vMnSiN5NZ+uVHnKr5PGZAmizdaXWH9
u+RXdG4GHndTwFh3mRL/6Bki3Kq6GXysTTJWMLvmuC3+dxxvL/iN+tBe3gNshIPh5KEULsjHFxRo
GEd4YJux45/KmoM6zMnxLgMsfT8/VHXRjiEXh1B9Qn3RfSoixQfMn+9EUm2aD0Y5e9xWiDwEQgCc
EKUuG9TPXOaT9ZQXLXvK+fqOYgE1zv6cx8dWzGvnbetPWkHVdu44PR56jumG7/KidDeqi0Bp8RJF
Z0We212oPd1uF0YKNCpB4jvfZ5Biml0c6m1axjZMu85DvVZQlBTiwzufZOKyT7LiDzCAzEQ299Av
gxh7v7djAB9Oiu2w3HxeGlTcWdP9UBn3HqVDimFn19USjbwUHptI7efAJMr6N7R1PHM27wXknzeR
j04v/1eEEbXHU2iOZhmBBffewhyjvGtg7GTq7BDnaSWW9UwmE023QjaptJk95EbxMaga3txHdni4
EL4OK05FmqUaPr4rguZ/v3YfrkNQS+ECg2wBkWQS52qB+V0tQVTCJ0JejqfGq6io2ibLVyg3LP6w
Ves4ziPJqe2pkD6R8d5ylA3GY6MUv/r01mJqfRlPi9aZP1Uvr+516qgz2Lai+VU8C028WejowcQB
aLYG3j0Bth3OmKi8oA+9B/uR++kcLoTrdmpATEZTtj0cjsBL95F19rIZP/9CrPJT7sGbLwGmooG9
+9Jd3zcnpwvHbKMmqen8q/zzkDkDKRCzG/Yb2yWnpl/JoUU2ACdEPmDpQKZvwoXFbh3XHdd8dXdz
/F5f49UOZh5oWwWdZeUGSar+SGjmgK+ZNZiw/kexCpYlYJNgz8RyUxCKyaSou46zrlP1O6QeEvje
+TVvhK9ZvKVDeLg3avZySQsst2fk9GHvyyBNsgGhA2B0JNizrNYBvYYuuUhbnqlWVzjcEG6HR72g
w6yuDwdktXUbwhOLl9p7Ety43FEjMme9rtstnsuDNp5Gk9BnPJ6D3iBGHSd8VzrqyQ4MsvpBwZBE
MQsQYZVjBsXECZwhRJH1yNRggqMnP9SdW5/febNZwpKw4rb4Rj07WSRzrmX9GGK3/VtcAaXxkzTY
EliJEFIRs56TCY6FRXJhCLUas6D4GvqfhPYDnwa4K8AEy3k/6WrpdCeMwelG/xobtjaufEzuIMAn
gSzv1R+V0LwEGY5y8zyeUKWghs7QJzLgy8ac56vUMnrwZfzeD8i5nysSNy79L1w9+mxd3fhdorki
Jzw0EzLjBL2s1/Hb1IIJP1/sL6rdzZUSytG7WKah/k1glEl3W79dTHiR4dWctjHdoWQV16n3GiX7
AKX6425PdABOmtmm7Rr526u/z4So1l297Eb+WSi0iIUniwY+AC5s6AUyvM8xAk41w4mr9jJnogrj
Hfz2AlfFZlfl2Xt6RS4GIijaJP66BYGCN8ET37MtqGxz2Eo9rcvCS3jOGcb/b27RS6BSTnpbVTSO
VtSxetQlIcEmLSyvMsC0KCVSr4lEaQEBvDznEXIphwTHO4S1HIbn7NO9kTJx1TJUs57t7RNQoSCy
icGM1wLdHVLDBGSsbatoY985BR3JGg9mhQ4ygDupY7RyALiPBUOCaILKIcAZqKBeVLDg09d1+Sjt
PkH7mcXw8NQnNfR3vX5PDfJwRJUuvjyhEmketlkBWhSKLFpQuoIQHtNsTcyKMbjTDjTUGXffPgpH
bjOyC/KMp5GMjLAHZcJsbdvKjBqi9x0jCknAoKlV1oeOXedvO3sRyy2FJE/lEJxMtRQoqhFVHAgb
KnMtG8ZbLQGwM4AwjjvtVCD2LuH2pFCtIl8ks6tzXS471pfnA5Uf5JEhKhc5Itn2VCvb9DFq1VbW
RSmyNHpRQ47qNpFmWy2XYV8nd3Vazw/nYZy/D4qH/vBnePdUM2ALdMMEwEaIKMJ7CgyfsA6slws7
yq/aGaRuVn6KSS2U30oRYWyrDmqjGVox0BFPhxWzsc2Z4o1iqXDTCAxiej37TgLPIKQ8SzVwbR66
LrtxIMdpjaxRP6iQvg85OFCpRbQYzs/DmNzeEdl83HopTFc3ZSYnTZSOZOy0gcY5gt0XKd0uMXsR
0USNbtV4OGaLdkno67flDYQC/LTZEYQvzshfOZzVAGqTE5ZeBSP4XgzlhanmAHG8khVgaVR2iSs2
uhcGtnxMX7BsubCEEm0G7glGw+kXOadLpxMeV2C7zDkux8MScCt/8DHQaOBKIQhllga9Z0mj1+CH
oAjVIxzQ15Pumzuw6gDlPfZkDw2EGt83WIyKaEGeHvbQYbfDd3FiT1LILa0kaiiYg76R9FVQaJKx
o3oOe6UAoM/ctngXhLkvUAyWxKMvSZDnMumOMDTxTmnyjyYtq8uxSuiMmFNd7JiS9xCW1XdrX9s8
35KUecaETgM7OAQ2rxocb7dIEu7lZuJ1t3DAX2Sr0px/ai1pSg6Vj10xwJ8IiuLdIRkD1VAciE4x
VZMU1tkX2PWobsBfGEy2NGZnYVd95TTMMrH+/wf1HpKjAn8ZJ0I6NtEC+P9CWv9/DRoMxA911NLr
5vcRaQPDqLTe+Nkmb+Sl9Akw5Ay/72S6AT5eGAlsWIbNR2xuOy7JHgVaVu8yrN69hP39DngUNsqA
kGjNiS7+mQjIN22sfxX7cZCUZXz/dC4Dqi9pH4KzpdsGwT89t22ui3gGJSIdVpTMRxYaZ4+7hDYV
dIVZFEi3R5TZUDfk2rTeWadlEbjfx30qdFMn10JBHdJtiMdTnHPEq9y8f4zJ6Ws8fU2sQg172obk
deVXJR6axo7gmQsMycTbf8cjairhMdDdoAP4rv3jZcc/x7PHl8IUg5yh0K0IuhgXSF9u2D4WXrud
kPblvo4quShESSR4LEU9JXMZ8VLhWeeG2QI1qC1TS2ar4sVHBdQQr8EkDcf6uk5Q91izgas6XPnn
JK9CE5hk9+WjPo4VMJMvXiQRfCt8ETv58w6YR86mCE3gpfCd5N9Z0GTM1EM7HSjPHDtlqbwnAJ3k
vdQ6PjPZApRM23x3F6hjIq+hBSv2mljn800khsJfRX9gYGxdQUbuH8nPfpbfqN8/OvWVHZYIwYHb
KgACVNXIFZRl/I5EHxPfAOJ7zSOe/E5Nef6z6lm62uOtZBRk0L3Lm727OXl/YU0BJDeM2gep4Jjm
wnNloC+gLRjjdH2ZbVB1naKE0BfLhg6/YEpZ6OHV9RSa4PyLP0l/FyNYt9YRfhwLtK5fJSS4o6dp
WQec63m06KsAI6r8YSgvIvaRti6TWWCalU5FowjmDCr4G2uFelOx+fEANs76i1YdOOuxYr3YgFna
eQxF4HOPohve9omnlVh1Tl5lll/xzgGb4SpBb2+tvxHk/csyBTMBLlYERfD7z48N2Kc95vv6hOx9
pF6/TkKIyvPbpp5HsA390dK1jDAgavUVQFFppqf260xrJNQeXbWQ64YjdB1QMqBPt3nht32qk9fM
3xMzXj2vtt3jr6oNm5wktZrKG/qRIpkxZsq8/goLdXawqIyoPJSroDxCvpdQiCLVf+ksUwIRUb60
n7Evc1cyS48ERPB1cJ0+gIHNrlKADd0azB4/bbEY0SLMkDAmDUO7NtJkI00izcOJpi7Rm1swImSl
zMY4D7VRUvmSFeBFruMPowszJCrOi0p52igsN85RM7/DNHpsdaWRgjnc9TWsXtNRZPgUrjq8rsWC
sD0qt2DPLiotZ8s9Zvmcus7azOztInu6SizMfcaiAUiYq1k+NzyieZnBSPDRRp5lORJDkG5bmls6
yD4f42Xt8nXjMs+Vralok4n+jZOuNaVQkLzHktxDj2MucNd1eJCWP5Z85tO47m1lSmQX6Y/SnrKO
jxedMcihamlhLktIdXVT732NkMzXb7+PZRWDulrlkEYRqqPWA2A8EH7kwzifJu2Y1U5q2zJBHqX6
MXK9MGey3RepxSX0ponazq43bpsQZHUCJ+jsJYnrAnt48HquEcVgjVZDtpHx3MSEcpU0NZlyzFDH
dTYra+OsGFDjm3plzRKhH32dj3IGHRZEAZQMlII7SpHkbYer6msIx/c8WtgUWtI1vuV2FQSmANvI
0+bRJ+vKx0dzagEkxZpD0803IW0UMaFJDj9XLZ5n6lpwIfX9YH0mxpgNEOloYibO9TxQvBWkmia7
En18O63wod1l0hlvvxhJscRfL4dILIQi4RM45ObGNYTSFgfX5r7pEtT5w7j7eSejIReupSRleP5q
pElvUSFK+zP5PBlSrihwITc/WDVvw0Fl2e2Cb3NV9sVExL4c8vUMaKoKGckFpwi9hEhDavV+5n8K
xvi+hKtOi2O9w8IqziZY1crQFAuhz5qmJZ4XAc/b5o4YjqPhRiisc6G4PnqtzGiBnOToUAuIjZb+
Byucmy04c6LrOO7ljItZfFzF/tM+VtygzHx047AG0LvQqIqK6ZYP3kQOnJX/92SfSlk31FnavjCC
tBRIXvcvo3rzwAVecclmfRUXQ06qlaqiBuExhkabooDDqCeBEPU4akYKY7XuOFvgnCwxMtOdOMfE
ci9Q62e4EEqldHsr5UYgzcjItouwqnxuLWEG9Fxt9PxlPUdL4OmCkx6NMIvFcr42Px60B3NmDUUj
QkNax9f8hUbxPCTcptUEv9JzkT8ndV2iT5MDi4GW3SVMtyNQ7jsAsGAftsEeyK+ffMbKHsOsT3gc
/Azgs1/fS0TtOqOiZicnj9jpgyPY3HzfnoM8Cz/Uaokrl3O1YGeV0BUoEnHalL4NsdeY/gUEFfgL
o2oUqMD0Kvj2lx+c/f4GcZqKxB41oonZHEkXS6pLNsFCrTyF0tF+abr4HOEJW6oixBc57IcypilU
IoWv5Yt+iXC+1y6kM3XuNRMCzYsrD9eVmRBFpJTxpQpADWM2hu2EHpFJIb6PGfVvwT/CzcGDb36n
nwHh0LchP/W/e2EqLM8Mn9tMil1CWo9/x6WQA4V2tgDbHi7Rj0HPAqDFhgl5aE6ttDJjt0kWNK3b
9r6azlcZ+LGnTZ79DXTjG9QEJhr/5c1OfklFPJ1shUmc/jtfhgTVhKJDNQbHMH6jAwcA9cKejwHD
itPdhrHuVwsoCiNfbMoeC6cYHrxEVH+yd7xauPcvTJ3wOQrr/3AmwwVaYyYylyT2cs5NJQE+TWay
T0GtftfnDWksNeh+psWeO+cBbIelu45ZfmbVPLjfrKjHQgtjXL4jvCqmOobAcKtrXEwQxc4xLscF
yuHpxOwY+wcx0NyIglqmUkKimdZL3V5jLNVOuH4SCD+T/Iwd+Ve715tOADqyB7523nXLUVokh4Md
ii1dG2PhM/lnQtuI9WkqSmcgmLI3KYrOQGPUT1PVitC0PxwjzpuTs/+sIsvYO8CWPrdfemdlV9Y4
Tx49pmb1QCgEc5E0PqqqoAgCOjFi2umcPB5POkigMyLxKmgtvGMptmM/vmpOmKx7wK50O+8GbjjE
RA3sSeeREmiHxlZArwe07adUo3+hoHXJs77YU8kxUWjXVtn3C/7WRuxhidUOEb2pN+wZTx3GA+lg
lq52kMsucxmZaGqEeA/RmDj4dcdHT+vDCHpifVGmzmfWgxBb56CliqSaaQpNkIk5LpyDuuFC4n/n
P+nBxaeGTWQgTisuMIAOuNSol07ucARJ3ImfKhHxOR2EkC8ots6Lz/OqyA3H7FSVJuPUN8tk6D4/
wgTFv4DTRMsw/9QqRZVojB/XauNZeTMqYzGDDfo7W1i5EcY+gqK06YdThqsNX8yRLsethoXHfPdp
4Sv2I7jXHNWAygCrJLPUdhtjak57b29hi0TbUa2cq3SnW3yQaek6MMMLIC4omR2y26F6YyT/FLUD
YQ6Bztx+Wy7ydqNuAZIvzHH5NYtlLWkpwWdF4jkX00mCWMYODpjjvRcWugHv4tQS3zzy/q1RXnJn
k6vyYJxvGxEk49Gx/w98z7K1nIRUviWDs9IonRujsAHiGhW0rAIw49pkysheMEV0GCkdwK1Yzl5Z
O2+KPjf5s8q2DUDSXRmqAjfFfy4F+5VD0ZZkyswfwBLpTmKwoYfBUN8H1N4CYj/GrAWJxLK+S06e
ZU2FsJRdQaqTMpky3WQFraCZKbkn/6hQb8TK3+Ov6/OerfK7dm9zE6Q6RJAOsPLmkdn0wqKWB5Yj
u6DxPg2yMZ+9sORHTwIGZx0Y4+JzP3LTuKDnAlzRUfCAAKyoICw3unrpV/4BmDGXtIXASTQiTRnq
FGWxCbn6qVd6pJAtxtCP5JPLoXiwm0WV0KK0GYc2AxoagE/kLxsGwBN6hAreHXRvQqpoKnA1jxuD
msmkivkp6Jwx39DHT917cpsr2YtOdL8AJdR0oLRnvhnIsI7/xL5CQHiB/V3CuIQLpXyXdCjR6Sf5
TwyUPfNEY73GL5kz+WF0Y+yNXeYhfbh3HBVJzVie+hwNDjaw2+gyQM4LTfjA8v0ZQDwTmvfTfCeD
xNhVUeaLh3LzXOJY81nqUUq/0TWL6n1X45gst5l6iHjlx1dorVGa/6w8JdiyCMjCk7nPO3MRoSx+
PO1nQm67Z/zmNLHsbfqp3BWdMfbdpjTJeuFnLkHCY6vTWJRNS6yzzmrCU/np8p+T49I8SI8SLjN/
6YXBInLe5H7rDBdSLw+1Q7+JheVItxnvratrRLPlFsvqiK+yeA7IGj3goFrtoaqOq9iRkkQVu1Iu
sjcIGoFWnMpj3PFYUmOOarOFwXdxp8Sg1I4DnJov2Uxk4a62Cx3f65CtpfweOOvF/cL0Aquz4DQm
Zjjn94MsMVZkrV/SUW89F8qQkQw37N5RC/S6Mv2oshDtSIZvLGv3rbIuOaOR7IlX8XPAAS9N6Uiq
TQozxM5y7VmwLnowEeCFABxtdJT2pmkFGB+oICi8vXO0HZEGVWuFZ7F3uKxnvGwZfZ1Exkc1rgqM
OjM/36qXvtPsFjfizXXc5IBE4eTQmHyqvDroJC6vH5mLz5kI1OJgJqwKz8lGvSNEvNwt6MY0fXJ2
AQTfnfhJ5y3vP3+D3Flh0V64iY7MYt0lQdGHFMwNpqxk2c+vZWRKLlY8sA0noUU/BXeBTiZ3TqRK
JYdk/TqUa+Yic6Gv1hOvkywdfMHkOb4VsJBDl2OOKZnzjsPwkVKgT4hVX1sNqR9q++upVOplsn+T
9rim1Ux8u5yKfP0x2uEDF5ro+nuRTPvBmpyqnof8+zZIUmZvzg2webEUWVyx//TiKn5PT2DY9urS
bHl1sslgsKBugWLWLa7d/kGkMCzsXzVTDhrQoEtsz/WNn6wJJLsKcYJrtSCwH0CXVqYk43c8SXey
4b9mAUY6DsjX0n3w17LAZHfrUiatUmgw3L6RSGhPibr7DCMvMh+x179h8hjYQCLhl2PetsJ1Kbrr
Q6TUZQ7onGnChg7xCQ/QI8vOXr1WVgeNG2Yd8sXkm0DY+LU5uNkdSgj1PTQCIWnoN2cjmNMUOcfX
uHHe0tN65u6wcUy/AtBUn3h20aFoRUY9YCiQixvpkKmYhbI2gI9kSSkgmvuMkQRQOBrX6XXx1RO4
9UqiYsVHa9xu2H7bI5SNZ+/bWBKhOp7Kva71OXDhf3os2efnb+mwrgEUjWCGqJoP0MPoO51lo4L1
A8ihWx2E9dkcE/5ovso4j1S7CFj2GZTlv/xMUAg7triJKKHgOPCPoSy230ZQXR7vRPQajJLVHd6/
OXQObAZweamLJgMkh47iQiUS6VKLgJNImYIRtipGUyqdUn+fYflWA+3oTGG/wO+Rnb+xZhsWhL0Y
4WIrjiu7Bfn1NHtNCR2vpUfp15q4Vxl2jAFdP8utl465oILYUli1MSNllIpLN8GyKZFKF/9wvNNp
QNKDPNGPSVhMd0YYcfev9ST1i1ZSetaMUAl2oxYnEFqte0CXl8i2K+Mqrd4eY37aRBIQ3MZeZIQX
J2ow2xqR04qSjPJ6LvFrassblWh14q/FqKux6ob6qVwn68SuzaiZyutIOqXuK9uTmcrOods12cuP
uDbTG0O0Vs0RyuntubPNS1vWhfLkSq9GWztlcvAxyA0oJduZw6diFWdthXJxB8Hl/LUiSdbZDVnH
B666lJti9L9cfB3yVdEZ16QzGMAAnzFc1xS832rdEQG+Dx/VBT0htxHV7zAtjP42LV7PueaYfIxc
JBNleGSMPgl4NGuKOAQ9Y9YgpSYY94R94GURj5It9kxhXb8KYWlcZrJ65NwCTCSkX3Bm8YLpoCyu
XflOjkyN+aDFU6FWqWO1liMeL0dpIrRyUyRMHm1sSTsF3SSN3tPoKlvr9NG/njmmuxTus22ns4/N
FHAV7sO/1GxaqMF4o3fKa5ViFq5RUEo6BvoOGMxde3uEAKK/LOk+owVxpUcD9QLSyZJeoD5XDKm7
GWf9+jEVnONUYVCgc5byDC5BaglaC7YX/+7ti3qbE/sB/6hdOzJ8QWp09nHW4y3floeRDJ4jI4AW
VhdSKEHJ0ylO9uXzMWPg7rYUYlLjI1CWubZ1pY/rSEPEB46SgdoLzoL5rmSCEr8eiQqW7+6SDWdA
3ehiCjiVfZ4Gnvz9215GTf0FLfTDC0rWJ9VuFctwqydE6AecT9wxiNRu6BSPe+m2ED8ZsyMDomUh
45ECHGLeEb4rV89hA3rlcUfcc7Gqn9+GNNk0Pbgswsabbxw2dljuDXaDvLSQmFlV3AHHfr0gBwRi
4GuTNsKnSEcumJoCEkjqY0qSg3LtvVaVizPiKDrMWk23ODFbpYug2Mr64Lvn9TQc/9uMYQL1uBs5
fqYXfL5WzYWTY483/ybEiPe67kHPvIG+DDtMGlH3gNhdOMwVaMU1rJ9gzC7PIdnCC5XflTPxlBw0
bSZf2qC3IxG7guc5UlLFyEn5PnDfa3jvJ1ou21gElfEaTx4S56zFNq1y8ac7V6tWp2OPwOI91yVC
J9cq2ClswGn1ohi65cLOtGa1LmujJmEfykl2DfFCWw3c69eEBZSuCFm4JMeIvTZWNKBFJhtQmxYi
Og4sMIRpQVlortDgfab2SZKKYOSbOIlfyldOOaAHtoegR+H0usVAEdLraCOXMnIMcOOD4FSbPo6v
H6ZsfWg2ryTLBIdFFyxd9qCLYka67OFjU7mPV+xO9uhmjzixiu6Ul86X91s0pxOZYk08z1H7fioY
NUtuacwtFCyHBZi+zXhJNA1DQyjG5v7kBgZZGLGIm+2SsDF8O6TeDFw3gIpsRVixsVLISHhpG3on
HmjEoEk3rVIxKX5WOcD88WBi8qkKZCc8CpExE5HZvhdm8/ZZe6XSgYn9qzYtwIxxc8gKd5Upr3F9
KfXpoO6DeDuPgmVvrbsH3usrautGQQJWjNKGqSBpAw15yu2u5ssFutPJCbzUQ3l6eCBNPnp/9ZKg
fZuFkzg0fEb5SqSgd6mDDs7CcvGJQKiMt1v4kqKTGzwAMvEk9vOH7RtgKB9SZnUdgeTb33paCHzL
U8fv569nExcWF6xylz1P3bj31Ad8rSp+5O8ixvqWgFRqFaYN49tMvIWfp/W/fJ9NF7wUiID72x/z
+8Rvs5j/4KAk60dV3hP4z7LlYWylmSVLlbnEnHbMAFxKniPPp37gjO6U+Xin966i+uKHs9WY70Al
a0sSX6lqk7AtUwnTmNkBI1haaYDG0eN8/PJJrvcFq2M7srUHfj/4oEf3Ikce7G/kNZbkeUNL5hCu
Ace0Qhm3GMAG2xIaTFafPl2K7Qunh1dWMlCbzcP5dYvYcoFwuwwqDoNHOutYWrbTv6cEV0vRabn1
UjuqvALXC7d2eXslsMnufMQTIimqnvt3G45ocJC+I2iw4lWxQ2l6Fz4nscJxdyIl6OMpA72unLIA
j0/cl7yF2gUZYEmP+cgbVkeAplBEXrNeNy4RuRk6O4jmQ3bCQn+9pUQJOglAg9GP45vnUHvZzth7
jIDdJBLaduc+b2h+bno48mK40a6CbkbWks+j0hd3LiuQKOYRRQulg5jeh6Juqyga/VeN906D5sie
Yon5UIZFHDyjq4Nqj/9Sg6T0weqmmliB8pG9PS/9vtOs9Uws7foZm6BHXk7PIrF4D1r5hRc8j2Bj
lpNxFkOxoWxG4GJnmxajakuH6jIfoBIL7hPvx0bPKgdacdA2hl8obAx3VTnXyvuXJB8gzOhN2Fr1
ta0HN8tYwTL9YwNwqfkbX9ZSg0fkH3VIevb0XHfrkq5ugu68fKSRFIq+8491vCx5kUXYKi7gHFC+
cLWoXVcZ/dM47Bw0Cehug5effnJAoHJMECRjRzVpLN0vy8qgJSNxqkWLKwMWAQmvf1+sUgyGtwbq
KmFkmDjCR/rl3Eb+7oPN+ksTqgMh4lBeq+An1Xb8iKBkX02vJ3Wsks6lSGaG4dJ6QzTAaRuVQ4Y0
oFSRNHwgtj44D9hVVlaB5nzxEide/jz9mGaCAVqRUZ6Xj4qdA34mQ4yd6uALXmEdUNL8EdNO950d
6bkS2uHCl0TKQqIi3EpKtc0aS1VVEN6MVtBCdB9uTlbh6XL2+7p4iAH0PbHa4SX9HoQkBNSlBNeY
nQbQjZz4koSWjoJ42J94xY3MqC5ozw/E96RDz85LZXBeIM6Q9aHtsEp1cSo0AcI/QU6eFBxLjYAf
vMKvDmJo3442kX1+de5Fui11aNKvZd3LehfDiO4xRJimI8Cu2VutKEvjuMuKHHKZyXoqAlg4ya+F
Kgcy9txMXljriyKINOLvwCktXkKztd3hsseiFt+e5EaaO6DxUL8EOdpRzqLs9dhGcRLOWowSkyW9
o1DUrg81cRUBLuH7NSEDP+aYmeHpREP2yEr606baRsfyC+d4pRN4aWwO9w0lTMOFdyTI85CXqQ7M
VcMNWWS60FHFevlwsqLafG7Ub3DLp/reaEcNthOKSeKFrFXQ8EP40k8b9QPRCzYotTuYPJyo6f8V
Zc3yctvDzavO9uMWTO5aJU7euX4Z97+vom9UKBIuFXDgx1zg/oc/LcYSjdQi4dUjWfye1W1w1esa
AAGvSv4uhp3I7D3+svP1WGvdUwSfA5JxG3QBaJKXYkl64/VconbeabWBQ+sLZ8XCR+IsltnZFuNB
HzgnriuGWYkTpzuir4RZPla1BLpZB2MVFWttEaOujwMiMaqSGear5VYAPB9+VFUxl6bptG9DrGUD
HA5aw8UVq0NbeLpK6w0x8StyyVYf0MTI7SxnOwq/luRneC4bTvZpTKMdg1jruRFJvwKsgAHeo7rX
TzFD0D6DcuUsAnDh9SYHaFk2Tw9dadOMesbgDvOl9+V7r7HQbAqPkFRnKz2MlBvc1n4hAwRwpxtI
1S++15Bw1eeKpzgp7fDlVIqLMEwCoFT9AicipO1bczIHEQMwoTJhhyDqAcvdBSno7Xy+nBIJn4el
gkIAI6Mdub+Xuis7B5xOZV7JYQL+m7oz+V0XQVTXb24OIhDZCEMRmyB3vDEwtbOzkbAMTwuBAiIk
t8EHjG4zFb1vkJizQQLQejt9zPKcGQegnJHyKNCV9+1g/773XG2zAV/otM2biyDSpIsnDGg9CBwL
LEUsV9hpwF8E9cXbEYEqnLi0orH6KNcMLXl7wja9mLTsfl8Fk9tppARwg8O3pfww51AKcxO7xjV3
ZWFQx9VOCfpdlj6MeLiXG0xlezrOMNb0Jo/mApJyXn9nHuglpDMP/MTkpIThEDyNjoWTtmO2oebz
kgxZd9ZWIwAJI5KHwC1wXPJgIAwgAAWzJJyueFdrT/tTVqZ4/LiEy9lnZTkPca93Re8mrZD/Gt4p
5xHO0Qf3O2T58j8h/HTHQX1q/I9Ml7Y2mS9n4wY6f3FzdLJjpQbd49PmpJkZZtZhjiAFMSAfQJiR
4mBoIyHa9zDh9MHmUB3b4cwgG2WQwziGJq7tDiw1dMxR8SNefSMh0TWT0LX3g+OSRrWjFbpIKKJM
lI7ZBYRJom3wTCdNxDkNnsaqNwpUQ2DmUYXACJA7RwiVgl6TR3UP04OG14kWFyrZpx5ZVTwEeKMl
Tk3N5nMHzEKEa3pdMaLMvx+aFo+/4O+b0xQvNkPCVod30w3GnUJHh509w+Lb9/eN8gV1cU5Kel/l
MQ33yUYCtOyedHntrvuZER/oAzQfTVJeSur9qABGTnWcIShaS/tKbcnGylDW3wfAIfNx9aYXXwLJ
QvZ4CtFehjyO3s6h47/RhmRx5ilY6/Aa3DUoIwKMATMZ6zMgnlhaAaso8tKDdXm15XUVVKsZ5aTB
GZoAqu9khUuryL8/xmxDxjPnB7GaKiKGotKjfK7bgKZNe5vajA88/DiC/bRG2cNvnvhxdfDNw8nn
zG1ho+2PC7RyfUlQ22+m5jdDUziy8jUYfSG39wlU8e/O7x6KVKlDzt9X+bknb/SRrMkUAQvhVCSD
vniLGUigS6TzdOe9RlRx/xBM3f5nhLgn6Zx9kVltQbuOELCVNJG6gACINzKxwLtqlvrbLBdLOyN9
WIpl6qadzwrtKu7/86cE0pgcn3h4TROnZbuhC2KcKPJ7847FMjmFHXFBI2s2Z5CvPMXEgV0T7swx
SO2fsGyA/A0oChnVcSrD+0JSWgKIMqEIFA98ueZ2UouIJmkgm488Yu/25o2UwMrk3stdtnRlVh1J
AbQDrAKumkfLkU5azs/hOuweCVn3T54DPk8DqWVDJnsr8YYDanKUqx3TPyQay5tGJRtupQq5pSWf
Djt9aZJBEFLtLuC7v27sSHRkcZpfXUnKLtR9jaqgN1ivNPuTkW6ihGLZXzYbkZLRwaBZQ3ePFtm8
tBFsAHuOMz/YWpFl1bMYnyvG2o3hiy6WMWNBSfhC2MhsUosH/KZ4vAv6T+GUi9RFo6mWfpfQorbo
bcGU42z7Dn0zikZOeYKmzoMrYdZQvHnL9g95HcNcJc/Z2vPnckfFek7JfEdboXeyf1Au6HCn1GYt
kpuiJnzk/81qmnfkaqMncGycEzJgqeM+nRtHbN30hrA9n/gGDrT31rkW9zOtib4RxQny/RY6MDaF
WzozN40uWdVL2SIvObVYsoecgVPuJG4i3AdzSBwoy56hQibxW95frohX+WCjPRxOQstgOYAm+RKB
bNTybhSMd24LvrSJEZwUyRvdQ9tUGHkDqC5j2U0NY60J6137oc5Z0Y+dgf+FXv8v3Aw2gMgmWmHp
TuXdQng5jRjUQBkkMybn//CfCaHAz5zIiCPiNR78iaUc17xex+qRpjinNWA5iIhdbz9FhH2P4xYV
WzsRdJ8ZN4bcerJpRK7keHdQ59Y47jcgEzEA/D6ps7vkZvq2/wz77cMpKd/9SQ9Vgfhlw5GTcgdd
6+f71ELcyB/18Kwwq1ZoqUcgmhES9NbQkcZUn/5VBmaW/KHF3QzJMyjhjRCfItv79fTk9HdbLElK
B+u4wW+mYdsw0TPApQOLZv+O+XSpv1IgoRmVlN4rfbspGXtfXNViuDKW7v4Ek0XcF5tboxka+cY8
t6JQc1/pXJ18sLOebcHeaABRpTNb52hX6vezFznGsmliMUJ6vMho/s8ENxM6J61oGxaaYJasJIhi
IXnF8xFcuWq178iCXRVEeRhHh0ovyQHMXnMElS+k3bFBlWSGzMSnCXT6ytwPZmbX0oHs7RSQU6Vo
xcwR60p0kZR7t3TqXZZbv30N2Sq8o5b0HKPfV/pooYrnoVS6qw/3M87Y3OqHQoosrVtFpwNtaegA
jyHXS6c7OOznnYGv0aslR2lRpk3Ugk8le3gurcMu78Dx/bvHTyWo8Gy2mQhKHM8q8jxhS32rjLxA
Jx5xAnpqA/2koGHJNJ2pp0/9d+5Z2q37Gb62yaovvonOBhnpqF1N+8mIiJbLXqHD4Ca+mRNPjyP/
ClfUZF6HGScEf6lw+kJigI+7VrNbUm2Sh7HgilcpWPmVfoq5MfN6tVWSA12Al1m4fm0BSFbuiJQ5
/m3ZmpefAWKOpsuFGqDwIDAtOSyXkIvc5RCNlHAH6cdMu2au3K+9Z9bOjdSOaOjurSMbLEqkiKQe
dcOrsXWNONXBm5ntBp5ased5Fc2S5fN4MXLg0h1bji9sUq6EuruGmE7FBqjXenQTFaJhluJE7YHM
6tH7+IGxL1IV9JjxVM05PN9dV5OwEENCIODu9Qid4xJBG7phZCEEQQBPYBYKpy/ozEHzTEssvRPb
W2yZuN8OBz+n7f8WqzG7jsswq4xnD+wB+9+HmhAy9MiEF0lFoO51H11aJrIwyW2/Txud32YY1Zgc
+67gejurkJEXWljZjdfPtZaFfhZL/8KUmvV96oxb6edG9luCuRykY1cx1wWeneFseGvxQBmkVA5g
tEvI2F+tigWz3hhdhCMWzoe+xLfIVdey1PHnlR8kkUg6AZ9Z5uxIbHM5SwMRKpZSuQfyiCkXdRF4
H1Z9/oo6z3YnMSCNGr4j0AlVqALRA1VMJCg11AYpADCmY1SWzH9qXAf3tlLtDqwyu3rYoGQmw5I7
vWSgXH1902RrAMVDmfp+zc7vJVde7w03pJQOa62dWXOZtsrQCYehGOpCx8IQRbmgc8yPBvzfOTxc
Mv58eXGRe6TRaPlUML4Q5G0HOsjYnpaXxZd2IK4NE9DXkflSINucrieqiRFFp1rdquGk2XepbFdO
nyOBpO4kdeeKBzIsWFc9+NVkyiqp70+6JaohO8zhwDnW7sG6Ih7gfgzfJu4ks4qb2/OnqDKvWRjw
JEQAfZAnhW5VJv3pygMCQTdVNdX+RIodY/ajrSz2NYFxv4A7MibwlJ7QylNP9MfkFCxxMRh7zhqC
xAAk6h4oUpWS5IYmKL40vVh9CCfKbFGFP9tjM5tjcTpydh3moo3/QK8PFm7XrwFD7tG7oFZXV2e2
V3SB00pBm8JhyWeJLgDlrgAgh1Ld8MFJkeTg1JiRBdiTurjF54U2j2ibBlSa1xYVFjVB6iVQ5HcM
WKSw84LHSljRTEq0JHogvhqIVB7Pj1X3jxrHORbqhnQ9B4j128rluh9p6GKjxr2tWlg4iXJ+i44G
nKb9/nZQccyBH4U6BdGshtHxydNTT5ESQw3LXJYrj9mALt3nPjluVTp/dKauZXHwqypfB7SoUZUU
lAoFPWJ41jKHLqBasOVLv2w3c+XgTmgw3jn9kWV4APK4G40rI6icbmPnKdFFflaxCm6rGAgPibKD
RdXUi8O3ZVJhTigMsI/rPwsaCTyT1sdn8eUiVQGnSRKvOom+Vq/m1mT4Z1YkyE3rhm/asrYqVgUa
podOY1TVf1FBWuS5QEMqPH2OrOeDP1GbJ+jwT5Pz5DyAxpe/ICSFzaAAUmKa1aWpHazCAS4KOHcw
UAHsMesQqV182gHBk9QAlDYFgNjT31NqtjJG0h+vjFGSrkvNzXV83GTLg6Egzf/hRBWOsy444AN8
m5FWssK9pNCSUdDLEOq765FHwXhd1Pwey+sKcfwRg0VWXj4p6tH6CXPu+sgjt+Um1WSFOjl6cdVX
cdBz4kyQvOE0dQtYNkIpeTqHgiGvRUe+CINuQ375q8Nt914bD7Sr/Z2xp5RtlQZvw4aIuTWUI00i
LnTqcYW2Ei1DTm2NF/HSLCwdEKpnMz2zgJww96JSe+hF1mNN5dJEog0cPBM7FfTu8aneyJ/5IGaK
KX+J3ffV2K5hWPeTC3mgPE7M5n7UzrE0lvaEKEQR1lzpx6Ve7CyrGuqKrhnuT8etnJoXywiXOjQW
kij5VPITlToD1EMQ5PpZmAGV5bCTFKEY8Vxkcgw08o/9YC6NWQNpmeaDxZF7pQClQ4VrY/s1Bi6y
s2/4X/xHLgXvsVMKMQ/pCi5LbnAQ8Gjm2hImqKyrYr4/SKeyxE7op6pmW5CRfKe9mUxev8JSkkc0
mUvn1h71y+f/UyK+CNm2uICaj2+ZDpcqDGQPGF5iClaxc7nRiHW+bqWppGjph2l588h/RfD0PTVd
4kfvpJpY4MvRzkgXPmf4AkMoDtZQeDhBugURLQO+LQJcN/S51kadGV32dQ4gFlShcBdkwiUKWBLG
9VSkU/jzayNbUgv1jELQTSD66mnv0M6XbZ2hg5ST6fggONbpY4nNO02ByhQwzGaFYOBdmypUyUhj
gnQfIK110+y/NYSZp1HmKeSBo2sDt5TGpLllAy4eoboBaGkFAuZ8ag4tDVq83hv+RAeSZJ64VLjy
nmbf+vgQhG5qntIMBXkLEnur5AF5Jw4eIYcHS5QRJpuOfFnE5I73VX8q5KvxHe0G0+0nuTKM0NpE
Td9xbXWqbHgIBa/xIkDNY5C5zU+Y8TFjBpsD90MU2cvohiMzVkZZdcEY2Nsd07OZKxMcogh7qZGa
dG+kc925hrVdOFVzeKfgFxZ8iIAxYXr4GeHrLN6+LBEOEwXZeNJoxjJpHyv/WhmgUH1x7XERfTNM
cNXRvqdBfK8MwmPxCumBK3IuvfAs1OdLDRU47z9iZnl43VBGdnPdxwLTNh1pyJ8g1cQZn1EA6glC
wofI67zrfs4HAwu1GEA2KP6brnw+0CbUcRkkmoJ075C1Q1kHxiEiwLVwy8P1HXjvzZ2V83HaKTj8
6ymBDgnNv9cCvGslNQVCic7HL/nlZdozzEbkM3NBryiVJKOVh3jErXFpAcj2VvjLZCX7J5iC1U3Q
xIW3Y+FeZl+X6gNYXgFD2RhZY4YmrUH78i6R8FlaBj2Nb4sRQ56xyOw1K4yj+f0eVVxPQzfS4jVE
ExxQ9qWSADd/mVEfSKdevcEgEyDJzdKgD3x4o4OkcTvcBC7a1FVZeZG2/YQHR8NpFPYjFLLKiEQx
I720YfW+V5FLquwzBKTfGulGeWewPOHDUjBdHE1aalslKYrAq5PHBCMbj2WGd3BYX3wVWXStAowp
yHcEuOcWDkhLs9rIjWJDaVgbC4LdqeXurW15uKtG2Se7OPXNrs/ihtx2XmmvaZ6unndWOkCar2SN
RoUZU6dLxVi4G53SIRQ+BI4Z62ol/9MOIfvd5o6cZih8pcOI6BqyKKtJdiUID79wKgdpMnyMHxRO
TYeFGAykTTBhx/ez+lTMC0lNDSPuQqKa0Z73TFEFNaBNdhZeMUCxBrlShUJlB0vFwjqEV8ZuAxwn
fixwm3DndMdD8IxX6Ze9YcPAhW6WO7OzrRzmiBvd2yrk6UclceMOdPBcR4P4xuvTnFooQLjO7RXA
PmyzVbQjoX91aaP4OKAaSbd27vMoJkGKhXBsmXFMd2UllzvXoQ09gEsW9mr0uVY4hkhJYGJMH8fb
IrK2qWfJLUQlCeiqDNZUMbSKRRJSsgIqWo3VY3bFMzwOZydL8X6a9m+u1xSaf5QoncyMHFhPtFCv
qdzhEyKI1fYjzdsAL4v50qqWT0gcb554C8Qy512WohGBkJoBYP4Ty8X2+1UaBBQ2JQciawgYDMgN
pIhn+pT+yPO9iHl58Tj8Rkg7JKRvG0oHEqUH2ugUULsLiKYR76Chm7FzX4fElB0LFt4UeAD52zH3
PqV/LD0faGhiGDEe4IkOlqDcepVqk03F9aisGw4J7dt8nZ+xtnb39b5c7K7OA0t3YLkGpz0XaBZF
mx9C8QAILngvkF/6GKLYj3BsvS7jbLldHddD1M29BKx1lCW7+oJiHvFJ2QiiCJwHnGW3l9DseSN0
2xvDMBZWa/hmiD4FAbeaLoVRmQGD7vfWvSvrGuTHgsSfmM1ht0G6wStfS8ijhDlSY3JDdJaNgMtJ
BsYCGg6oIWIXSgtkcl/+7OvWmi2GJLNHkxlRMVzbIm5opqz+xkOF6Ess+2xEjwECysqo4HvVEgxz
9G5SorZ0qAnIRqV7CDXXIe8xs8VJbF5jDrLz3LKiUnQp12KC9YQrrIQD9f4bML8DQ9HVH2bQGCrx
SJnTlatIBcfZ90cGnatf7W4Y7Is6ygmkENgW5tHhNqbqVU7DHS0W3rRC7OqIp0i0qIpVlnJVW9Of
Djw4u5gMF0QdHfKnv+3ix32nKyfv6B+CPssAz13ZvRq3GA+ObtexasnFj6juPZp6Lf5Chuot0mKX
K5PZDjuC+oCSj1CgwRVX/ZEwqn40pGGkmSNCA0ToHbe3+UN5e7hoRkXcaUFPwjW2UJExwdyxVm6f
lAlxRvO8wpFT59+eDfvavZjy3QyPD34b/ifOtA1ftoFOV5gU2hxB6CW7wYrcYswV0YT08HJboOBr
nth50XRQ9xtAT/pGd/BeL+/YRZMvUW3Io04dUn3zobxypV6STyNI7ZukyfIw2b3HMIwxjuDhEa2b
hh6ECvi3DbApSZ4GpnJ1IE8SxTqffaVneVn5+jaVL2DQsVTwcXXhABMGQ9sMLQI7phFfHNNy6gZ7
pBuIZcaVtDrjI0yK5xeU6q2H5IRyiIL2/kG50qrnPNlzLLEpsohaj9hv8LTrymfgyyzcHWVKEN89
z9FaMXG4sTPyR9v1HjgQn2hab34FABqzzPzCDl1U9lNI2BOAQ44KTjKnU8XbQlOdasEDGwBQHodx
gEkMUk6+gSUJv8D4zpb/yeFTRA02G48UnMDjy84fFKjnNNA7KXzDHleXZM3EL2dbdSS3ugBnIxZw
HOGJ705mYFeh9sIHmWWnRKMju8ELdj0QfbNOHOio/q6a4XHgdaEDVISHtYP31SKpPn6TpwppM2eh
MMNNrWJw64i3aP9ajpkw4yPfRDVOHx25/w55VFP7xRpf2JH7F844+ii+03LeCsV68uGRI+FtwvFw
CthiueC/1v1SQQTOvzF2C6SdjyJ5u4ahQK8CW6aqwhM0Tv5wOHp+XolCRW4iIgblbuJ7mNf61odn
b3jnWRzrQEhjJ0trSVzOWJOONZy2/CeqMekAZqXt0i5qotZEaPKYt89/Gf7tQ/BUFvdFpQVQk4c8
7D1EDx+qpkpbYs3sClINsALugVR6FXbBbOcC/29mACpzdekGs1KmgAWL+2swEevb0WoHFIgv145w
hLqJfSGPznb2zvnNdPf8oBVHAlL7oSsEekuZC/hHd+lhDm5DoxIX7rNFfe+GcJeQuf3isSYLX/Q7
ihr7SYJS4Fk2hDWloaqMlWwTr0JQXoIUqSDsonvevZYUbzo+ZShiMqXogL6t8du48wUrK2Y1QAf2
royeIoSW/1QnaYYv1Yj/UUzuTV0FGY6aS7woPgD5vWyAKmFXk0y074tof6z51UjQbOWBuIVlldVM
e05jPEopmAUu53Cle6FFUMSeGzS4fDVb1AWGhdVRT0vy+shwYkHN3g98xmVgr1dx7tatmbAlq4uO
OEX6vScqyMF+aR6CA4/M58ml7vH6pKo/eDYIGle2yV7lgdn2KMKl+Ocjr3W2nIlW1xwfVVJ9llB8
6U9vCXQ866ka7aZKbETIhw1iBG2kIXjZ5w2NsQgF1CB444b5xLUkfAsn8rjpDf3zP3q4QUJxGZnL
YClAOkK0eFIdxt/Yul+88jquI9zm+Yj5q9vQWeQ6FkUMd8S8SXtQzyu7pozQzezbu+lRkweCDIaZ
Ov+kM2slqnH7QXIqRTkD94gjh7LXKCnjWb8awF2NdtCGkUCkcocT2ZzIuj42uRnAeEOi/xs3vlID
OnqVUh805wBrRgJIUpbX7HVX7Otrsin1qxZ859G66rKck0B8bT5uP0Z/+h81bIfQ6mS01Va4HEc1
EmxU1VyGYbMkr/GByXN8LMCVlDVLI5U06gk+1IRwY4lbqvGtEzmIzP7stWm+7/CBHvRD97Zy9UVq
e7XjWYP3Yfpehr5+7lz0ivG0rYD3SPAzJByebOAHkTdeWqU/yORx1ilqpSF0PzN+qhMRU3PPE3ej
3eijerhVl4I08Wm2fbroarfDqm5oeyBoQo6pUm3WEGhbBkozExqU5u3nOccOCIOLKcB0hNEXLvcp
FUZBKCdKuupLdxsnLv40AlXvkvpSFHdhV4CPH4w+uKXcPxG+8LYhGKsFsDxmfWcTkYAVmC7ZTNRP
ns/44d7Y9Io4UQ+/iPD6zWBfExwxyyP0spAkKZ0E5eYp5EB7pv5mtXtVLHJ9/UeiD5yc+aYuQjZu
a/AUcUK3RrYozULmJzxdjr2DUu3YJJbAToyiMzVouMIF584wIYRRtAwpC0TAXTUBbEcbv9IrHIXM
esSPjzTfakV5Z9ZzdHbcjWyWpn497YWz3fFq3GPoI34sUcGBKsHpejBwbU5tPrRNXyLFlM7SSpa8
hlukDQMnKIszej8QwlZZB4f4LGFDUQbt6stxWNJLrHf9n+nZA3ul7GdXp4aE+M1nEnNymN654kw2
vFvCgPjsBRbjED8z2s5UziC0l3j7u/L1bTIs1yck5ZJzyvF1QvpOK6MQRpte+T0SVg488u+Bzl1H
m8SGypkb58wfZaFg6orStvs+2sD7DUDhokLmR+mjc0R/r7i7zg7j7y2URE9IJTzfDID3tBcyuO8o
bHMawCVFTY8lrETbPJfczMbX5im3Q7y8q4Wa3RCeq9hbnbtmE64FGg4Vn1L0vNNYce8Qsa2VynTA
xrJ1u24zKips1G4mQHRFsqJyK0j9WwYQsWQfdst6sw/vVIeRSHZMux8Mp27DAC3dGg2BDSVvnmCt
bUvcOMIMneY+tTTjIdkFVVYt7RMoRMIdS0IWsAu1Sd9AwtM3VM1S2SfnErNniUmbuW1ydplcQYpj
YcKeA7fS9QAEFTjesrt4Eu08ediZqe1I5g6GEpCLR2cT/IW4hx85Mu9ms5OWBLUfAlOjRLecLhOG
cuEA+XfDQXvV4OAdUcYAoP8iHIqEtDjJmb0NRv14t/07fVLqmSyUXhUWqddG18ndeyxvP25Q7Hru
CRAIOHCf4bUe/IpRftZIVBj7EdqW11wmqByWJwudyQcc2EQ24VOqe5A10+V+AMRMK4dVVicmM2jZ
z0twHRSMzexDWhgoVw7bJIZcIU4KJL4r4/VVNFom0c8GBlof20p4poql2KGQbAlzb3gzJ0xzjaTO
Gsp9Sfx3v/wHDQ6uXZA2hNgeIiol4VARX2w9k3WmnjQ1nrEIKSv0TtmLxW6ELHSNhP+AJKtZt3L3
rK7Cmn3VbxQkGSaMc1iwaaY2+UuEUoVffFyjUBoTpTn4icVLxQ7J5CmatMvve28yQJwc5T3sXZBf
my99joApDrGBUR1oogyu/zFd9MNL8BQG3PwNm03zDrsIbJqG7xg9XYttEuPHEqpdXR1M6H/Fbu1R
Uo5n/VJC/i9C3VmQ46SkctrupKj8wtW6p5Ud30DTKSxGq0sneqsj1ISoxaR02E1fXeKLb3+F10jr
LRHPdFQxbeOBNVM+kyupQZRqAxHQt64N7QRlnCDR9tyywfGzUryYY5dEewkMM1nzr8yywvDwW4r3
9FxaUaTLPmvfKUFc//nLyrpSIBr7ESktIL7gF8kV+fLK187MA6i/9ouoo75VlCmMQz9eXXh5S7PN
s2KUNFpKekqOafaFQdLuEGCiRk3X2nVLYVtb/I8JnYk9ovXqN58i5yL4zEkLa5qklYzwEz+WMb/I
TfSbXIc/h2G4EfaGMHDKpGTX5AbiGSncTw9SQ4D4meeP3ezelayB9OTgJojbb7ehT/2rbQ7ZyDpv
Bq1XbRNiQP1CaBDt6DydV4aogv+ry2frgkn0zxBouwKAW/kxTMxNU7OvENAtVJfNuPoOhd+8Vngz
gq008a/5aoERaQQUJAvqImYKTu8xtbKjwrZuaH1+8VbMkFJw7lDKNgtzXMqOZ/JiBfnQ/Bm4+C+w
ECzBMP8Wadbnx0ST2Jp5OTP5crNHKbESnbxCBEH5L5hLTAKRxLGrM9cbn2PPmfmqn9VMOgXGKLlg
j69bganmWOQNuWhpzid4BRgGW/Tsvty8heW8hj2NiRG75aY0cU4+aVa3WFZHEuWAVj4kloa0gPaQ
NWdniZENIoAezgcq/u+2XFFOeS8i0d0S6Y0X7yvu50v7FKx08FZ2bqnCSrvb5AFrFc2J9FYpZrdB
+I988mPiT0Orxw5GsmIR1fR9L8nK4PSBRmNLsLnvdllQnO2pJCEnjmUIOcn8ZzsRnaRD9K1pIT3j
jcN7g102ScL8q3EH+4ZrRQE1snDVxRfNpvgIE7RmcfT3FusqTi2LSAVTNXuyXHtHzFgkSB58/m8o
l6LdoZg1Cz1VvGPouuW/v26EDfsm3HnE65GWjbwFMmpO1po03MxmnoyEXj135445asZUqy7/FehT
BMVjTgJ7OOytcif0DJl1YpsFLTb2AajNTJwn7Jy3p0kij2D1aD6ImYd5hh341EpvFZhfGSyHpqqn
WZaIO+6uTkay4H8ML77ZmAt1NWmgZd5uSUDWA8vCwe3Cf5PV4V9r0eciY8y9QJtypgCNzGz0jCYV
FkimGRP31+faEHHds7/9fAZJ5HDT2wJ1nfvOrsjZ/q6RiBjjWfPPNy1e6hZlzt5TH2SjT0DLTMCF
FDnnhsh2g+MI/DSHuB4S84NSYsGE4aNQcWTUBUoNlkyziX3CAjFwzP+rCHisT1074HS3oxG1yh6e
5MV0SJxWcipb53yrlCKUN5pCPcJnS2VLuc+D5HlhPfvV/tbOpocaoBZ3508g1ERtVJuH138dJniJ
+iAot9yODNYZwoK+iRh2tAjSEe5L+ImjXvlQ75dUlqT1Dufyv0FcACR/zBphU1qBVrPWoY6Vf3Fz
Zaa3SonORk9G2xvtvIZ6aGCulsVO4hHdLoAXLxWTI2iQwZSh5DOLP6EGSmCU4hcsLkpT/+cYVZBG
FeTdH6LoxkVOaE6pHYy0Qv58pn0jyIMWb0HJOo/k+VjrhnqV22FMKip+LRRxtbB6Gx5td5hzih/4
GisDGF6Hv8cOfFabMNRZYT+J7sVaezO8TTjODpMAkJRcshC9oXYrN68fVblABWK3ka8J9KE/jaaH
EfLslAUKb77UMPPlMOJ1mQeWq0jlJxYn4wSE7ItBavMoUYBUVcZBtaW0VL4KwHFd2AhfTDSz/5he
7d2930r05Hx+rdIEShmuTI1w5cmnih/Dud8XW72LMSYtUdI3rTGIEz8I65Q0Hlq+gyVx4SlQutvx
VbQ/11490BFkchozg2RKXDque7wwDknBdd6CK+rfrQ+q9ORPFLDSD/hLnXEXeHhPeLrXjTUs9Vs+
STvkbjUXG1Gf4LfDVsEkPYPGi+UwFSOx885Q364wd9S7FMh1l5U4rkVPBG9qVq5Ph9CbO66bvRVF
CZkK4gyZurMfIK6sfa/cmFTLkWrrYCshv4Fe+OkUMnGH6MJIjt89LbOCaXOAwn82Alq35UR/admQ
Oojv4XhQgvYUqiDix3tr+nfJq7HKggkYVswxCGOqGObEldDFTHieQP5YjkTJ9T/izClqQFHwMep7
4r9Dk1DxFgyFIw88wfHQ7e2TrB4jsh8cWSKgcfoNgpr4Sah10KDWa5xoHPkDbiCJSn9hGdUrRJWo
r4LBtPPVTek8rHtnGS9FUXoWmKh64sd0mSWLsVQnY3PURudYq5NFbP0LDlBwPan6+nXK00KPESLR
XMhvJ9XM+D/KEF1y6F2G4zQWMggzBi7DuQWDZDTyXT0vfuXgyZkN7JXHgRtQsiEYjkdduFCTmIzg
pQ1ssKdGFzuZOwxEs82wsmgfrip9paUMGbw3Xavn+d32cthe2VtbFXgf/xBc9a82AhRrmjmkvvx5
oM7kJ7MMjhh/OC09DFpBE5EMi+0LAEC6KdNxNHL0vqv8OWhIJ7+a4zV84jz8HFiyMfTesMvE+aPT
2H1CnuFSuDCM/lKSjyw9admNRKwgXiUZwYbqyGBkq/jI44MAeehjWNcx3+vtBxElMfNCSkEIBqxe
xkRRnkBiVKp7caixS5N6HVlvEfYfp8AHvr7+hIEqrp9+rvuehTbFxPgQxakXXNUaKCXeulcf9Zj1
cT978Q+o5CeSJDvGOMBIrNNpVtiL/V5q0A5r8s9DwiazF4kkx8EKhDgq27Z+N5r6V9i7CFtc694a
gC9j/pdsrkQXXDwDyhNWH80/Pxkj5ryWgXfoplo52QlZShRU8X/WrYfl1ohiJyCLS3cSUAXiF9EL
nyTuH9FcF+I/06T37iDqp7d9Rfc0Z6+AFxhKMqB9d+t9uBRTKhZIYXzLxsPyaOKkWuUX5e3awJS2
JZFzEwknQTnQA134G282HnK/E+TnvOyyb5IHF4j3+kNL5WHDE0MpmTARRIyrekFleOEKz1yTuEYy
HCM3M/9BYhH0W7tkTiYtInB/1GqdqZwPtdkS2s08yIWwflCX7Jnto+X7kayi5/2/Ke5ptq4Gwljo
BjOrQojxfUzFe9Gz1qsJP4UiG3NMwa4PzMaOO6BzqAVxmwsKrRYdjQy96McOk88k2CvuxXHekjYS
9BU7n0DJPdH3H53N1d0VUpNNqD3EBC2mQVg46gTt6L0BXwZtrVUsbwj9/cMVx220DZvuNHTrAUJH
7FP4ujKS57oVsyKBIT/qvGJVhiNqO8YuKl/Z2/rRbxofjS7z4ADc50q6O5s/ekNUvreRKMb1DlFZ
2q0UQKF7P99mgmdUTzqEBgMGzwTjyMwPIORUYvLp6bMAWt94MxmCdiCz1xpibYaH8BZkGM9xnhyA
r0bwnkEZGDKvghcFoOgGvkPUosEb+B5sNEfMKLEYFn/Hri4br4Q8UZGoPiIl2vlC88uOcYZHyL6x
a4TXZyGkZDcvAqKg73r0qX9i53jj17h0wE0UNmOC5brdt+ikMLi1LNU6BtikpD/t1abBs+uVfdwu
BlCooJqX3iD5OKFVNn6d9IF+6lKg3NBsdcAWsqlDMHpKdfkUDhx8aV3vSTULuLXx5miYWcQWy7Yc
ETRamYJ9anP39xflDGTN2E6I0OgmTmnH2x3Te6wpN25kj3pEyIBrwKk0FzGjiKsXpjIuxoV6LKFd
crFbp+KFngUM9gmEZ+z+SCBVgCsZT677cATI+24kaHk9cfAPVSSy9lBSCvo4b7zn3lVZTtBnmZv/
2u30i5LpbGy80dm2af38gbUQapsvgnoaFqWdmSSJsiUvYIksZXgsTa1XALykmG2EEMMG/H7gboBI
SNG5oL0lWkGLIUYfClfWogQJoeghKQJ/GO1ZT/Xz3aF0lH67mOAquh5atLK1Hv822O+8biE9FdZL
7Ywo5XzYtlbpr+oE8IKOQ0geus/ISBHmUtT7pqq9gsxdi1Pb+4EfhVOyXbGvpUZbMDKrfHeROx4q
oQda1SSGe9pY4jRhG3vOKvG2GM9siooKHKEYdErnZVsax1R0Mb6g0IjR0tp3+ucSqzyZMmKylf+U
oMwnjv7TKcFTqsC5Xqwd3PBC1YE3liroid2MgyG9lwt4mMg3XnbJua9IS9cSD9fDyIb14Hq4dPBU
/ALFFP6MWNPo0kQEqI7qg6P2eV7X8jHcIEdSrRA1gnkGqTt7gl6rKM/fEaCEQcO1hnl3CbMCeCaS
dzZ8izKpg2driahLL7ym/ITn8yluMCpyqZXJf5M1l4VPA4ZcLPv1JMvuSqOFIYWlxqoXM22Gh6Bd
qWomeralb3P8gyqLQVxSPJWB/IaqF1LwTa8KQx0jU2OfxI5sXxtogJp2Ig6HQs9koptPJrqXrzJf
fV+b57WNMkbYkMSIp3etV7CuDOvqrRjS1P07cZ2l0PtcatGJSorI0dn0QxBrdu0s+IYgfj2ZQA1u
5pgoMIiKOE7NpOJwtRgeBPfDjfNlDpTLtY0CLS1+gpI03kTlexY92zU1/dJUE4m6sWBsavxt/upL
XMCVhq7pgXZZ37zOIEo1boADqhgQsGjW+mb1rymuVIN23lHwADapt9TAydOnDQfbYZuWPUUXzL6f
6lHdcVwiQ9tHWW9WRWwvBFYfEe4gHBb2EFbWWI01TWYNlEGOH+hVGPlzbTyF4vFSB9MZC+FYciVj
vYfNEfqmKHUkP7w+iryhR1WO8CR/M1MCqtiGRqGUcBxpRQvrbhIAVE9pLBV+p4wgA58ZsVUQkazd
WgR6OeQyTfcIbWKWTDDGphBflFi4ASyg6Vwg3xkhZLR7EA5dUKnVnkhIIiXPgMH86jESOciRbHro
c8r4RJ3tPDPZLL1oT4hmFa/T8KrCpTXtytLhiDgR6UswWWwEhdg1os5i35A3dzdWe71mVz5PLl4Z
KpRKZnh+OjOv4qZCT4gAPEBUrKtjLZCAcraOmVZzFaDUL+oCr560KnRNxbwWUlQrRLG4Ch3UxiTv
14UOj5+MPSouSnn/Hh3LhMpdfeEsWqVn2YW0apWwvM+PzEfXKcFBEDanxTSdECwtibn6c5Pg7t2c
P67nMhlyEw9cMYI/o+YxGaUhlRzsePgWSQIA0OT5XEr38/9vMUy8f8w/inxbRZnkracbH9hJ9ELl
Rk3f2sZAy4UWKQaHIqArelexuwVEJmg06RGNTSlukijemqDvO94AVJEVCa2Ts8ziHyPgqBs44UWo
HlNQG4FXDm37o5yyLXmUXVvfLSM2m6Xz7OuL9N+kpHIbXeb/iGQef6wUwUgEVFMdEjGwg0y1O49M
dDRz/z6XZXxMlcOhMCfMhI+hWj4jy4+abL3hkOF5WfwRJ1mzN+O6t57OQDN1YSpUfV1CnYfPB8qp
Vp/oGvDzzJZlii6CoWyB2A7RZ5hBWZrRCFwNgicM+2f+TbMHmqFBdeBxfBN7M7F8XBi0FfjwVo0n
2Mb1+NRZAhJnC7SkV72iwrLYm8G70G39Np2536WFK7On81ceFjmSBnw06nj9szb1mE6gb3oOdRK7
DriSZrCIW3MHgGvAFOQ9PiuAg1iT63VR/4vgbE5f3ANFQabMNNG6+EhOfhD56vtcDrglZjFxwowd
B7125m/H2BBl/yMrPcFT4KEM8P/+UVBSwRVcJYtGu5aoAP2/J7BpP/3ogHPwuMjZ/Fnb2wrKNSgo
wRJex10sVB1UT/WP3laJ4/sVwDO6RK+GF4PgBzRChSyYxao4W4Wz8M0DMunhvlRc51+xH8/5GYcy
WVAWwgn4DuYRea2wMzHb3TEyx/N/75r/ZQyTRBFr+USAaOoIy9xqK8O+v+po6VrCtDBZ4z38IpHI
M0v6tcOkyo7qaT7RevNXFcjqIDjjEMbM3yD9p1EbIBQO/V/N4UixpN9waB7zxw5pqYbUMXi3HFOT
exd8D+Ha9x9Y578u0wU9A2J+4H0klh0PLuGo7aZNXZV31v6exbnNDwCH7OKcBRxJ712x2nVh38RJ
r2EsyQOiEYWAfgRSnFGpJws9qGvRMhSothWhKa/wgk8Y+I6zmO+DKszET0gon43UT9R6/gKl3ypO
fi3VuaBLktxxTc59smvJWkcxn7Xwu4wTHrYeI02A4zKIfs2JA0aKol8bQdAgi45mgPz/UeES3GRx
bmjwDGneIXv3cG1kY/ZQkTp/rgDASu8aYXrmNOqeanJY2jyvjCNHI7m3Ys4dNJi+utJt9luh6oUW
vuBvf/+jHTWK7CXXKcF9bNHW7D0i3BYZB4bpzUQ4IRx0VDZSIOhYYpDx3K5Q/YDHdKaN70i2Odjx
QUuHAC4BblRDqHmvr/74bgzVBzUdWc2+6sKm+Kk867zHj6qC0NN0kCs6gJffIxMyaJu2YGRHqJkS
LN8J9wbT3e7VszLBwomC8lXLg+TF9sFr8gKJ6oocMuH5KVnWuARpZaCf3TFdUJd+4sY1ApB/BevH
/o/unn9bzlQfoePmDBM36sFEo7uMWtYGswlNa9krp2NdZx3JwDKT3iEzme6iWB7yKnID+EfrPSCV
JmdwM5nV7aXvuXj5xzTqI5kFTja41yQRTXzCKJfbvbIEFVFBFIOcKR374JDVJ7eIc0hfmvUAIoK+
9xFGD4fAToWWbejcHzUnZbetfW9PTkSRz/09JjSklTOg5ccII/PbSbdUqBDVx3w2H0lVyg0DcUug
xpT7h7nfDDXSQiPMK0g3oGV8vO2ggufI/XOldng50gADJOiy33e7GO+IRZd6Kg2hNQSdw78mzen1
XXX38/wKw2tLE7lQeLG4bLV6ALUYe11luv8KVXG55lk2BJY6zM3vs7pMAtrEEyUX7D3unS2nCx/y
HnRVilqZLfj4zqlq/lljWG7ERbImUEnXVedHyPcnZhqwjibyR2vf+HOw7jhJMAAJWWT/qNbV7Pb3
tGwdDYFyL99ifZgZjioStQMwRoLRHBqxY0flUlAf8GLblluMZtA4boMjbwKi8C1jHGdagQLPGLVw
D6Jo6Wy3t1sKN8L5DwBHATjhegEhCiGvFUpjxg4Thek7s9AQItOlHcDG/282yCssTLSfejxNVnga
jnDeSAKMUlv+F9OUH95W6u08SiljML7EIyECQE7spyJ7nO9QNFtzcuMmLHBx/q07o6NsfACRYopr
uKN5u06gdO3WS/KZ4uGEZRh2HC/qSUH/vZsHpdonquq6qvGQODjINiLZP3An5R/pBDrCOXpQ0eTv
UuzRPPxMGprdEe3UPfTQpRTcrHIdlmdHBXG1nIJrMB1+79vDj9EQy9sSXUEv7CbBHF5H0iZ/nGKH
HkA5SfAZb1MDKCxExoE++yHJIeegLmSa1o+YNk9KVP8BOyGHi75u7twG6Gz4WCk3ra66LHMWVKGs
8WkE1X6DC4QHVvD/hMg0uY9ttkByCWev/nwFY31Xf4ktPzavmvBKbKvAcPRGzKIkKguW+cxdoaNZ
UzN2ZjRwuXRuoxmWFhA/0fTfv6o45kwy2BsK5LHmdhhQPCVmxpJZP+5ruVHFxNTZB31s24u0olBL
PtUr2aiypTjvZO5cviLb8IRdOo7f1uBEy51y/UWmRSeUalYqET07aGQClYzDjfTE627GVYJXl4Hl
n9bjVeSFAGRtM8gUfxbZa+HduX3Vzd8DfR0lAACnYTEdoFYyzF+DQmE91Rh1lADaE0Q4Yw1o2Lvn
gpUCjC1+AUt5JxK3TZrIAd0+zQSH9a54rV0revMDUBFeHDSy92JD6nYNKvQwVJPeTb+qpxu2L+z7
5NtZT3DPwqJjoSpv2dZUu5iPApfGzDqCn1GcV9JlULeOpfE3M6mLZVku2HtoFG13ZtX1LQ9Bcg4R
Z+Kk9d9S/ZGBUi115nJiA3py4wuRxNEfw+SOVEiYEYOlbBKQrhZf4sStsWZWcqUX/w9358pZmcZ2
97Gcgi/0PvocPzsmGDUNxZXv0zX3UF2vaVe+WWrPeIHj+4RvK/JfzJQvn6FXny/BcTmLTjHyIZBB
eIqsZm0Y0NVnEVxSUbJp6FrfvwdPzf0xmGM7Z98fvoCjYuUY6ABzfVVlEsW+SolE3KskXXRqlsIG
oVLkY7/jDF8Ut6XaRs2y1LTRtcwDeBn5sj0PuFmME8Jo6p1VOAtMoIHfGbF5poiiKu4ZfIgnxdtG
oAZ/4UWoaooGBf0/ZCZWk3y3V+4QxQgyS0YWSi0RFLPxnrmVJetRXPzqTTA5s9CB290bG/KfWKHk
M3FMmc2eGmTNCJSSW65Cpff5/pQeeBdDw7Fc9cYdGyOc0yYMSn2CKNq7fnA2Ly38vtk4ydvIX0um
qWM+Efo6fdPrfxRTZrE3JDRnJ1tLV+/ihLowKfPjaVwKmZcvkToWZmR1n0blKNO2fqW6Ni5eM2XQ
lC5JzYGDIh4Cc5rBASxLBUhLog/EtVxLFEpEA231EPdDSy2vx2y2bifpzcoZ5YA5sM4Jmwv52Ebl
cP47RE6cXo+Q/Boh0DS4cdpjGCGtCcBhlyE4LzQe0PvYDrJ/QO786ejefDegIoWgFtJGUdZBBnc9
sTpbX8WuQJqr+FwUI5cvb0VQYvUSx+Umj24Mc45Olyszmj5hnOlpXo0q+LrT9U8SK3fO0QGy40XG
DJquv+QmcyRgUJvgr75sx0PVSL2LKkvy3vvhxExMDzu2nY/gQ6y9uqDVsjkkkywAlUwGyWuE4SOE
9iTrJFS0/+KSrT7LthhsfE+wY1yFm1mM0Ry0LOZuFYCwmIBzY/Gd6+8FMx9Paxda21equKXeFM/p
qJlxM60W9xrKjl7MulvgnYe8Kf7LEd8OYfQBdNY9mUZECaFkhRp7NMRAbAep0NjwMwpZLKmwDloI
+WcHOczuvvG+T7q3bbN/DjaCuk9Xkh5cQHy/wiLLxdfCj28vJTxk8RtkkbGOkRwwj2bqnIFAfMG5
wxMrkDuaXuWEGUiQI341pXeMo6jtZzLeGbndgbJJpRa17o3GepnLgMc8EnlUGyaUdSv2inO/Ppoh
cG7DG/AutdmeXtibT5znkXLxrmlX9I8SpVO8hEf6BNwEql3+pT3wn2X5OqB/B90Izaufi8Wrww6N
ATxuCoSc6OIp/m7DMRcWoWHoaXp3hoqPODsw4OCzK9l/LXbppct9lum0wQgTu5jZpYWr6Fbpqa+O
LnTidvqoQPXJN7ddEM92NdGmw/2qrTdi6Z1rMmqw0jf1dfu3cQdrHK99VvNasj2e6JUip1o/GAko
5ssD+pIaXtqSJZBCedhXnYQKqF4AeklThjVj1np29i6U4vDjxQGjozPgLaz5qNvnU9wPe+GY3sIS
HFSkW+AoWKiW0wZhIx3EvpDwhX49JsaNnteL4Exo5wbQPXv+nN41upNAB44mLo89RVceLGyqk9xH
24eornKfWO3uR7b7LHbi4X99aAAwmnLG6/yLNMrE3qpKxnDjyFfOR5HJLB25mVplfdzAyyP/uzO2
3L5fUUsOoNpr+/BHrRVhsCVYJ43j4OfkxCgwBi3PklN63PzGvN3Gj5USJvxBeoPz50s/jdGYGAHW
GR2ZAP1shNs+BrdfvoknghSN8GCt+LpyZD/MSB0eG7UBJ5XqCzPygPd0wo79uKQGpCHudhNJFRqr
o+IOIE9vOMeMv8t2NAEX48fhhdEuj6ZMy7PcIgZYfsChomdJw7PK+ALs6v3GLsDAXSdAe4ZQGu2i
szh2hMGRWsNVRvG+L+8mjM/y6DSB99p8VKWIYP7hlFx/J+NMwHUfLCxFbgUhDM8rxVrmRRTXwoRy
1QPlgIqnyGNndHfsBDz0gEhV1zAuhGL5vpv2mHDZzyiJuWXW0EA8dv7UGfBM46Ynh5rMO5fwjTWb
g0myZmRfa6B/K/7HAtKSNgX7hblLqqdz/bcK3lKQ5DsboPnZaSvs8/SRZIRoyXwVNQqQ+UO3D8ph
q5M2oI/7WKZIcLG6qRuRhpVs4OS2AE7PCgDYxn8O7gEOuyBRVMe3GcCYpNjR3d1zUsHImMwEz2wV
Zl0eOdfFGR/mVBvN4MVMy/uvpJRVKYZp29HLJ9FzEJV3rHQ1CvVD/795z11p1kNF55Ibiv1Mx0PR
kfk9sQxsOaNzhDbfOi1+uKe2f17QimW8vQXfkl/6t4bDZlE1/uK89kxvfNpVauz8G2M15FRbTZvS
5rWY12ngrggabPwI9PNfXsgv2BGKl/cpLT9er72FmGjSui1IbRf4fT8nWbNqz7p5p72yLTUt+zG+
wm/umDtAlGSB09AR39G/di5mPKj9cUWKmuns0SACat3mOOPH5rPbqmN5IqL9CPv4SdgUTocndU9q
d06QSwNpfjffmgkMI58HWggCt105QzUet6seYgUlm9tK0Nfx2eFJefgdFh++LfyV1fmydR8Zfzax
91v+szOpWASofaDvHmUiHGSKyePybKLWBFYhMaatZiTiK5YkjC/ZlnOKegOAmUbDmpkQ7qBqfTkt
gBLmuVmIxqPg2S19C3Z1Wn/4PIZU/w4TMxK8qCCmDLs0A2YLsawAazsC1e89dnB4SeMp8Sw9JiUx
xoJqiOwrnr+bJPca3Mo8AI+DAP5oTG+Sy+JCamdIQf/t7HhFLIm6/ONrIVHNj8z2gc9M6eYyra/j
Edy2rnTd9iCYWmJo9C7qKW1j44is1Q/YpvS9OQVeN1vG/fyGoGAR7XRAI37DaMn98QFvLuDsdxcE
V8CMjSB4AiybI7dwTDuap0J6wtl5r1/5oG88/QBmQn7R0QINcGulUCxyFFbcaFXydfqJrZT5YN62
UsKZaPJR1qk7Gb857SYK2rydJk4vDeI1ftL7+5T0rLNhykaG0C01mn7ocPaSNJG4th3QElqpoLln
z8LWhgBfxLAsC+evi15/SzfPQn+AIn5WKUCR+h5Dynt9+j0UOFmyfAvWSUweMIpmsPtMwd3Y2BfI
xEo9bcXNwQzhvnpd2Hh0WVSheGyL78UOuMrrKBe1sNnPD+SB06o/X9Srsnmz4TNvA9JfLZWV2tCL
2QdPl9VJLtgUT+BWR0GUHwVz8dCPxhSCF1UF3D4UDoSCrZMf33D+w+JWztQNJ0pRmKv/T8a51slW
t8oWwJzIXsW2/WGW38m1cw8Vb+eJVKGGk0SHJqdwY+PmJilBQ8HCGMwVnElIMez2UcpeCEcaxUD3
K6gls3KRwpM6kSx6MFrw9VrJ7/W0K1R+VrtdT+J3BvzvAwaxl1jrpZ6UrILOswKXS1exIQvOenpn
5AThmp3GQUf17aDUeN95QXBaDoKS5na20MGBJLHY+2TT3SCvMTqpiup9kVUUieVWjDIuTrXRY8Hb
P09JxudmyLHAULWgGByvxKh7ogJ+AHu270CQ8kyVlj/u3ThDs7dv2gCXYW0YrkUOd0ylGMqyObaj
s5uhwNxHmcVVQ/VaaBarDJldbK6vP+7GKhibZmhBOfTboasEGWPKKDb+j7QVah+Os4oouFdeyShH
ev78xDZnrnlGj8Np9sTHrC0fzuP0xSpBZerjN07auyMJgA/y4QsbjC53v7w51G9O4H0148LAmhY2
LAXTCHf/y7OhQmAwU5NqMaOAxPITlz5pKlsBICNVj49Uj7Mse4fr7IIDqpGCJW1CMqGDhn3l8PsQ
QT2/PEzEZZ0yR77nrjvrSKfxqDAwkDz+4ak5qPpkU1/3rV8AfLPdWrtTzbX4HeYBC1ldMnTp4/O3
S0rk5y6Gfy++ueMdp44Hc7dWIh8ZsgYIUIkKrdgrvrcpgSKViptb8zOTWsNp/M5rcFRc5mGT8JHb
bsexDRXgNHTQtxfNL/8PSUxQRn5E3MfYmKim9hOW86FRZ8EbqaJnyMnjgCMFBAHKy6ynoyL4G01d
0OZgHWcpb6LqLv8UQKwoAklo4nQfyq1unBsPAH0TuOA5+89CqhQNxGwGCF9emIWLFh9QtUiizpiD
PGjB73VEImNshDU1TR+OgDgLSmkhU0ECl0qRceCARzhd1omZqfgSRP3hgSnyYORn/48Xagear9fb
qxy9h/onsaUDzp664NLZR5ydCrRZNyyFLPkoTuundyUIE6VAteURsLnXt0lyrnjAlmIdJWXicqmd
eAwJKr03hC5lSxshbJg3rG0Xr1FTTf5nqCIDU2N7mBFn2J239z0KkVLicBRyhBgw1CDfpEkioy0/
1xoQLQdTASFbzIOeFYxVGHZ/ZKETcjXC75pmWIhbWNEcrqxkwPxeQz3zej7MXZT3wmd/yH/AnGcj
w+Fe1nRmC6XfgloJIr4/0fxR1yAwl6KmTL/5HqqkZNRHOr6LYU68DP7mfP7bJpUCAm5ZOMzxFwBE
OG6cXbhYKGwL9bU/PQ82r/JpsDAei4KgKBqq7Oa+0qKcwpDccAaQuE/7vPcngRqj8GG2SX0HuKm6
MSbGqhFZ+zeyEAxvUnuDYiHmABQFdqcAtdFMhVWqV5VhTDRjXwOak6ez4KU+VqKVEzwiL7UCVK2U
NR0Rb4bmU+WRyVjULjANWxYtQsBVX9o1Y9R3LvSf1d14S4CONcthlQCrfAlnaCNsoljk6n+o/NsU
bMj22oXHCFLoBxBLmPev/XJJvHuRevpYLa+AJMH9uucuS26bzyYmKm5QrOGpuCe0NZLDJqRN3abC
5myqqiCd3BLlV/YvtWr357MLls9Xk48nlAQygUptlcrNt2Plhl5rmPdSP18uD0Ed25Ymq+kVxPsO
SBj65RielnRYGYK17BMBdJZwBIpEOQ/IECkfkEhNi4m3LVlviZ2IjgkfqyW+oa26fEfsEiCgkUtE
fuDykrWrmlaZyjoW3VpvMTnQiCMMFTQTOJQBmIeDfd7sVhIiCaVtCNYW84iB9b4wItHdQlvAo0Hj
537MxELa1/Yz/xxG0HLI1+buBT+3MbxmjGgcy8A3b7GXxwtnIRApPnUxS+YlFDkO+opgWQC5/tHg
z+oEK1oRRKg+iSuNmZe48bmnziHK9wt/EGbGD5NNC6Ia0bhrYZotDGEMzszc/sFE/grDfoEhvdXv
aKnufPllwF9z4ptOGtqFRoFOuHI4z4mujpu49yVCkC5bV7hnHXBAQFqh1FzegTNR2KxBIhXBbn66
FR/jNO0GyKvnk41Y56gYofI/0ivfvg0EDZjqA6K6/pD1DJRPJ74swDy3fjhdI/LN5d3ZKezeNiIj
zBOPsxmUXXC2CJYiDJ1BRvMmVGcenyoPHvbgZYlTakBmv02AkBrdhq+ii2TsBNalThQ/PUkYWgsh
0eWRUgIRPEGpHiQp/DbzBl9/v4S+E8En9tj1A3Q1Z0dwOtRlHT+GMSr9ly1cjwf/C/7uNjkuLLoh
6ftlPqnlVxzk8pZMjmX9+XAmdzKQ3m1Cbtu8UFY+gRP8VJd/1J2HjUyvKFeMHa3fnbL2HopKgRSf
awALFxv1dny93BTm8mv9UFbxv8BLi/BXayY4TuvDjpmQJsb2a9UgM3IOt/1YppcXOoDcmc6SnfGK
a3HZjQi6KzpjZUyLVhD+aSKU1mWpcSDBRxsUKsD5sauU+bxKP73n9JUg74uRnxtTf/Z7lLUUpv27
VmoDZJIIRUfhS6RMlLcwddv5oyZLhDAQ18K61av/zDL1WT7IGDtm3ILsgNWJQwmqF03b9wPCh8qr
H5HDNyI1+2cBGmDDghPPs0GhWijzoDUkunXl75ZdezChmMlJTEQZc1NgU8UVkB2EWUEkzmh/Zs8G
lWlnou0geQAaKZ318hIgHqpOe8i9GUb+rvPis4pgrUvyGTUrHfeGPo7yQVVzIGFreJ8q5BmRS+Is
K1gc81MceP4x/WP5Qm9ks8i+i88IS2j6noZdiPGy9msN7Qn7X0x7udSmNpEI1m9Dq68PnInp6vcm
W8ae3V2KCYfMiGFzRBvGEQqRIbAXE2V0zpJtbf2kZlkEtEkSdxsWyOTo3HNY+8psupOM+JdoEByj
OvTDaO9GZVEK0SDBSP5PjCuqtJMEfIFmdK4+q3Q5cFLfS0mf+19HpXeuu2fiyalbaAuwpavA5cp1
90XBLbhlSaXB/p0U9QP/9m1cXwF+8KvG9AlOUwZR2BORocdGigOkJQBv2Woi8BXU2dEKYRXvSwpe
H6h8kjfeju3TIBmomRTpKvcyPs4Y/JzKrUCD3j+KGKp2D4UjnQx6lmvspj6irSQS3du+wSjul/wJ
BA7WVIMixFF8DXPZVkWqkBnd+UQvpbIErTsGiiMC0P8iws78UNhPVm5S5TOs+Cuy93iJDpsyXChR
xShs7/HSJN1o0gC7P3chMZyEyIkjAqEQGEr4NLnG2N0W5UXLM2Z8k31XFVDdXjJCAQpRQp8Q5LqD
xCVSvGY0VrfuAPlFF2aRb30nar1k6+qK2nrKgSYqK6KLz7KCTevU3F0K8TLy5bi4X53GlivfyHJE
87q5u8pe+pZSWJGWwyKlIwPimDbZ53GScjwZPOwDu+F/Jh6NmHLUPJfsOSF5F7tHxu6Pfr5B08QQ
z6OmZzyH9rzlRcYSKJhHpxCbj0921Uf1XcXfu5hSDCdite5gDNhGOv9rD1FNy8b9wCHPKq6KiZJa
2vX/ezKRgqNpegQzFP+SnduEisHfXZlrV8wouLCKhGXIEeI8v35b0bdGvm7Oe51Y6U5ieK3b9REc
wKrXHNr52IvpXxhIemH7OCZrjiyzaxaSXAz1NrvXFFukB9zrj1qFdJISIDWYd4K1w07n7S3bjAfZ
VTR57HRbk+2yeGP5oGBJFhSSPuQ+ckx/fOLckWGO6i1xvSDPp2IfwdMVt2/vCtHA0JyigsHKU4on
cNwPN3yixN5ZxbOqM7VYhipxaZ6BXfV2sw2AbdJQ51VnvqKxxQPMxqwshYag3q+eCLBZ4CK6oTP/
10BsecaXEoZJmGMSKvoIDsiFCDkYPakVp773NnMNl+zLid4/HjpPEp1NvF1jASg4wbC8Vx0mqqQ5
w9WIaR+cauXSLoZ9xY8eTmL7mrqh4JSvZxdfvDNLkbhiXANwdXO0LqHzSJGyRV68g20kJ8nv02Qb
i5G0wG4jPg//f8pRLLF/PgdbJn7aqO8Y5SwZc6YAI7XEyLxjfWM+dGdW3dF8wslYDXO2DziqzlUc
nrmNpBGxeL7pdLa/0Ns4EIGY/g1tB3b8E+lvTcIH5P0U6Q8kCS2UNn+7Th6DCApRMW3+cll1tSNk
UDXU+vsJ6UsYlNYFqIM26SyvOQqybdzvn38SW2Ot5ge+0XOKtSJlYhc62dC7t4YzBp9y5Bv6qkqJ
bHpHFAM8mTicDBMa14HftlwNv1CFfFxzPyOJMJl3gRB0wMLmU4KZ/KOQvAzv0osts3dOu3DxsQSX
hPKw7vTCD+UGYDQU9tCOznM6g8laWPZCuLa0UQj4jEOqeWfx2x4hjuZOx4VcOTthwAar+7fOK7vD
MEC8H3YWv1FxD09VkPehkdRtJRKGgCmrtf2p+iJG6bgwrA8Z1D99H14s1nHuX+enS8RZ5Muoduge
mBleLZTyjpBsaUbZ/aD7/1jljB4TIbXhkut/QK7v2X0OWv6QgkfLf3puyJQ2sadQCHAiK+L0CQ0H
5zzx/fzSQXOITvZizVRebL3g/v3QC3PeUoxD+jCLdPNK2BrOZG7CFn67ftFtRa5A4xZBfE3HTFKp
lncsLkgL60MzvjSFkYRUctmQnpYaSp1B5nyiNT+aRUODbPL82/+bH2/aR0BrJSvlVTkCbt02DzYg
mKCOhYKI3kMHs9KmKqSCwiHpu/6FHBGT8kxNRiMp8nSujBempltSEha3DA+Eadr/HUB5KQGjrCbd
X6jFr4/rMc98AO/xcWRY7xFGf48i5ZMht16Ok6blvblGrPUacVYxQOw1PGnGfwCrr7NV8eXI9KiZ
OcmRDFrGitxtspGk/zPkQy/8iYr4WSv3Mm7TULOcuOpffawaQIESVG1LcZw9FPJtWK1m+O7K8gKY
Z5eh0eiPqMWB7tl2p46OZFbDi6QdyezW+ofL3yDbMS5j/k0lE9kdJfUnznyDZkz6se5TQZwz0pOG
KXkIX1vncuZL9Ayhwk/9qTt45WOuQH1wsPOpI5DBZwd3LgV50qsAtQA2YNRER7nNaZYpeHkLOY8y
8EisQjwL9N1msaYJedL9yPSCnHq3/pdmBbewiN9tufgPZPNCmHqcBhokOfn8+57d98jT0NGsUto1
kaUpg9HMzIEo5IPM9sAiY6iTH0mzM3Lmmykm1y7Kv6oc7c13YCwEAvG+4BnxB4SUZ1CiQZEt0kUA
Ku+OQSO/NwaaQWfCmMMAKOH5hUIcuT/Lstn2rR4Vojz5jHmFSU6TFIVYLAH8QOOipWF0yZqbr79Y
O0YjWMGyiuQ42ouSukt/kIU4JJojOz8IP7CzFQIco+rhzBgpRt1LEdc8evNHrg3J+J8nNwsyLNFk
RGf/2aZwMD5UtuooP7iaaWQRWDQ9Sujo9xVAxHOQvEoEYVYgBydmxqTBPbJW2A5pyNlMm+SLVpH2
rVBqRgtYeHe4p8CVAQ0zoFICZ/PZdgjYxl8t3Lfed+pro9MhFq/wUXqj/dh8n8e6Hbm8PdVmoMa3
yH9ijpEbFd1xLABTNsc7x60zGr9pA1UajhbtRjZG1i2JJbvL7YLkdhBEIZfw966pOdsmHriGeWkU
FJHLekNnnoNY6A2F5n1QtQvBCqHy/0uz8YKqv+Q419r4/jPrrZulRWkTq3ztkhdpyFLpf+7EYoJ0
AweiJ/N3Br2PPoi6ua7H5XF2jWJeDzr2JT+gKnhzMj3Ep4FywYdpwbLuACDiwB5j2qb26EIYeFRA
XkqSU+sAj9Y7oC8k09RKHEa0z3iD/khSzBT9Un+PhW8NOQQ3ajIBGkeo0O533PqftUc/f4dwQboj
xPFAeCAbVZ46j2TCNDp2K96i4tUgxtBWMjxjervNW4lbaASv8/vjzW413rGunQrjZNmibWjLQfY+
uzXNnVapBmEKfYE5G5xds+bX6jG5BpvO5M+u2gBfnAHTF9YscIJViqKJzgIKwm3oA6G9QDPuM7ja
PvBDe3IChBRfDuPZQ9l31mi1noQB9Z9NIFChnLZ+25AgtQRnHs5id1LGFxBUuh0OM1U/EUHJDEvE
/eDQe153wr/lyIW38dePDDhpM67f7i1tNlu3wRsPYNnp5WGG9unjWqFNNBNBOZtRGKgxOPrwRdlz
Hw4F4OmO/NV2PDzSz/nXECrg6PMDqDQC83saDWJwZWFU8GCa0MW5EMzfTMm7XgfPfIOdAD1s5z/y
di1kMKAWRiv7HFxHvtCEXCSWybMa3fjoLpZsSuzj2gJhyjmr+zQX+Clf5PcJT8QiXPS6jF0k6onB
2fam77eF0sCU5L9hkoSS9gM/FEUTJ+f3gaTMvaZ3mXJOFYdwZMTSQ3gG9ueZ0lE6HJJAfDMlifgo
n1e0WJ+LHLwXC2jB7z4W7Mv3i7wG5aAemO1h+wKlD44rYH029DELwj76FAdreHoQn0Y3GGWt6Lst
WVmzyNj/7Z8FUrlOpEfwTVjCE3vtjivF23SOsxbU8Gxl0Y1V1Ttvd5YzV/kYA3EMGnmBkMimQFrc
VS5UsLOcWzIkBPPpICsgO54Us0ZM06P2MZ9t/wu6K8VkmK9re3dSA9ejJn2WKGeSiqCmcN7AVvh6
9T7WmncQNLmBptzdVIzBBPJLSk28dCul3gmxFC/wgJmPTl2Q2TPb498IgqYz3FBwPwWa8KXFzUX7
g3CRfeyzDAY0J6ijU/ALkybofpC7Ug6P7UVxj9WIFwyfv/6V6qWsS9mNBpIzV8DFB+aRMvhmjqTM
/gusB7+PRxVZc6kHkzL6BAv2j0hXrAzt4UUz2BGoJNU1J/prp6TTpW75ZMfYgLopEDowaylwhXnR
jTeLnfBAkhDFXfUPeYE1csaWUz37HDnGOjOd0cwaGL6HvQRfJWZcuE00L3E2dTNieOnCQspoGTQH
fexagjlz186qnwAICqoN4vW+IZ06qlUKHwbCIeVlEVhvOK8bVs1sCVgNk0EXkrzRDisvhpo51s+O
Gpd5FqacCEjSgi1FdGXukrjpJvrevXEW+HdU1mXkDefB8WUEAds55m+rPAyRaO5UmfPYbAdGtq88
k7ri/VyQ7KjIkJrW8hwT2tXF8bcdDzd1WNPqGH9HJJcx5NK9q/9zHBR3m/KcWzOlGmtbbdq/fbjx
vBl8esyzStKzz7xf2WHCqMBzVgqYuCNqLocm7VXzq02kUqbjfNL2Ajovjh+aY4ZTMtEBKZZeMdQh
MS7geaiLZQjXvTojrLlZfgUhAlbFGjjf/5npq5UdGaP1Gq+RnTYTZc0/ulT2iEHnf/B6tSnzksAi
/slQuYyUnokNa//0eFoz+ViNIGVB7DY3AuXAyk2WuT2+Y8wzkgmRGogkMYjh8do1X9pqQwAODvV+
eT7F9GhPdD0+GtK53zWNTGeG++inq/0RIraRxlZyOKMMktdRZ0JMfulZ6XIsxhrlPCjRu8+lOPo4
dGXmif3zeyoBJqTHWGxltbJ2uaiRhxeJVz/95Zzw43FXhT3VHHBM103AEv31YFO6ltEdJlRF6tZ9
igiyDSLpfqV05oerwZ8XX4bRvJmAf/eEzhmHx6SDePHfiSnk5HYIqfl6QXHlkT+8pi+luVvLJeED
mG0XvZoDOSVh0S0ACgRCXMfWo5p6aWYQ3pYX5Oz0tyEMflLiOzMqFuqQKAWzAiBiVLYbun5PEQ22
DsULbGWcqL3bLzXMVV8p5BBETn7L3e18maj/UEXka7FXDSCeDZCluum9mmap+f0QK06esE5LK4nm
BADycNtxmGOuc8edlP0S3ISi4jW+83k175h5njFcVJjtFnV/hximt/EW1VJXm0aJ/lTHz3SgZ4nn
tWG10PpTEpmr1kk/mBRTU7taXeZl11/WcOPyTsywpYJONVN1ltf9ahP6gjZv6Maa58e5Q0IhGYES
qUS8CPZ82LNFLNseig1qZAuN19A8RBy0gQyAz0Nte881qlfv62eZhhErCMz+VlElk0A0bOHjR3Jz
WBt5EH0IJcCCSKEbed7/oa9teg/OaBXZ7TbkMFax39AofmRgmObmfPFZkyKlKR/KS8HpKw37gRu8
N25Jx0SzSnab9qCRClesNG8qmbEjlRz1h1WTsSqGJc/GdBZb5+qX6yJhVvgkcRxOPbgiof9U2tt+
hZNa7l+0/HBHuy53Qw/M76BwkiESxj6gTOVP+89ohVRLp18Y4O40qTJ7F4xMXQfC4MJWjaX5W+tX
ixz+b4LQCsEbW/oNDgC8qDl4i0eLdW78Rs1PyQYtoW9KeoLeE/f81XNCNaov8eQh0jTkkWFlX5EZ
X6S7H6r7MPTM+/gInGzxW7fpapfsSTmIZLDSjHGRBthQr2aWWigmakKis5wS1ZFglBnb1RABthm6
QRIJmqoKXlm1vw6VFCdj61tQ273AQ6cwJbYwYbouTnCGfaZE8i6Zn1Q8bptFZ64WxuslJCeyjc7R
81eXf0+soK1imQrbH4IfeIg5A7IawtG+RC8EAMKhnC5tzx2spBEz3TrqsV3mmgheujT7rIp7Tt7X
Y0MQ452HjmueEd9dxPWaMEJBXI+EMHvXQQ8PVdShw82sgnMpYWGENca2MDhVpICMs4kRFnrl7eaO
LB3mVPxMARGzQ9uvLIp0FzM873QvZZvxxxCSEppgY8xlimUI0SxW1oo+2t58tpVVC+ywOx2UkcmG
B+FXuehsfFGRmEBmskBlRzWS9dMVafeLrdrk7hxqJ0du7uk9zoHw3osIFFo8HXi5pOYGiwDXzyg5
sSzZYXTXxlE9OFzsze2D+RiVrxMwpaWU5PBF17q69hpIxi5OIUCn7hCXWjMQGEjK0KpKtZ15nwZt
o5l72IJcVNNbW+eYqwCVNBxD1XI64vPDFXAU0SzzpjaIjm+xKVm2zNYGSbt3aQocgxeKBpgMSQpk
Nitr17sPjBAhyqMckGFGRbBRaTm813gBv4SsyYBTIn0R1tyfCKsgRfacpRdv2ehdODLdK2bmIyfI
sFWXDsJl4VeasBMNwQ3dT5iLBjjgyuol9qScVcZw2TaYz1qQ6Q05RX70Q+kIy/SPwy+9ziP/F01x
BXZpV1o2E/ua59ED7quV0vVEwjexL33Rmy9x2/euKRMhykcQuFI2JU6/3rocSEMvyMnVj4LSKVHm
+oyqFBNWpU46mxWmvRyn3uNu7nbtwqeMHGJTVq3fpq74rGuCDXhLpFBMQwCLowXmqFcOLtcf7rgf
t7pl5Y3jdsFKME1Ca7gFNDabhepwbfLpzLMD5jGeVqkBfUafFbvZgNQWTG9UPrlMmFt6wi3D3w7p
WhBFT774LOmb/zDBSQ/s55P3IUGDTvNkaaBboeYIkkI40oai9lyi6UYQ0JoOFbKonIEruahS7E0w
82zBGASN0+OL72GEYORwBE/rj/qNjbDFF83xTm0kWxgq2j5olRF0mXetftfsdVxf4aNwxZapcb4n
01+iC+PLjJgsgO9RMm8GiCD5Hwv1Ikent+LyJ1hGjkPChyp6q8C1+YbG4SXYO5Eo/oDZ1/Sxuqwt
Z2ZSTriLYc++YwE5ujn5VO+sglRP2F1qCBBm51gfS8EzYznb2XJ29MpS4dIPYQU//GhnsOlUj6/Q
n3cRdj0zxFA6Hfhty+czLtSzACj8iLobf7UUrBef/qLiY5mpmgLlsel8zmyg97sin3OF+tyJrtet
v5JihwfNDKydDI3wQ3qVpQf7pEWcxb+wTmAH+xYYq70uAD5WRZ+jxDpNZPV0yMyYsIwEORtIV/0K
axS+6QEZot7d/BJeA2YrgDcCYCIIaFOkntV6q07TAb7mDZEpQuJq0Y7n0e9LMZo29S0vUZg4YSBl
OFxsARqSHgDt/MuVH1iQ37GFdIldhi/2PNC8WakY7ebT5zAT+f6KePjJkOB2p6wZuXsyg/TwuMNn
5oH08eCWXgVng/NeU7b0vrLS8paSUdDcx/5+EYFp4uh/+IZW/X+2Voc0S8uZ0SZod8VVWOX04zUn
yHYNExbkcYQ4uzKpJ/V1yxlLEAOMVjIMDiySBN0GCYT6qKmy59xe58k8FBqwGN6Zf3Yv64ZrLvER
Oaq+Ws7zXYe2YaV8YVlQXykuefbh6NwePY2twKWulzVBAy05IJJZ3uTfHKTfp5OF4TVTaQ1F+kI+
+1+rMTEQHsiLHQQ1L9SQ1NOv2/PT7evUvdn8dmg1lqbYf5Q2Dks6EmJX3M+QkrdJC7F/NDkyxeSB
4bS0uQZAdCyvc2bQOdG738dY3wmSeBhACN9i18IrXjQpQY9cVhUB4toDWzINIf0WzQqUxYSpY4Bq
yQQ5wVSe5paIqO89t/386CdLQTsCiV4o2Wg1AhZhYFZR6FyrFl7QEIohjC7Y81vvHMZQHuCS09kp
d5IpUqCml8XXgtkP7XWECveWcqnxSUYvzmp6uRyXnEjwia7aM4IRW9PZ7nW9tquihXhpaVa+/fzC
yszHZs27S3uf9g5U55pw1Od6/Z1KCwx7tEoSGViim/AmiE18i/++LEMBvjNA/E10ZSTFJ27dkXFS
Uf3/JRQ45gP0XGoW8r+FTz9QnzTM/10i8FiOcRRhKgisJ2nspYPiry+ggDO0zsO7anbw69VThRcy
/Kb8xzK/1zwtDo6cd283cWZXQkJtUYaA7oXmJTv4zEF6uJehNwJCegATuYGvvQ8BhuaX87BQipIb
1/Ps+AdBj4oUK8isSCBo8IapX3BuzXQD2XPXPHtSpna/xoUGee1LAErZ/SzHxIw/Z0vTmGxL+KVq
bzbSKJuCt8dNLTB8VPoh7tcuo6uyFl3qgghZqkf9mxTf0SXvcDGijrAVyWRshzrjG7TLYxqBmzYL
z7BQ+myUkJmYZ67urHpt93dQ+K4/uMZ7QukzdgEvoEk5A8sl+mnv6XgvsrZChcYFKGN0RdAMgFBw
UlKB7qJlz0P9MxT/gH2nDAoqCvdpTG9YoRv+eh2+pi3a3PR5klDzXjVxumEpJy+hW0huMEWQX80k
doKUROb6jb+es/PJyUIjE2J2kIUboR2mEei6jqXOvLbnE/03dLfNa41v5sAYCcIItCHEXcnQFyBn
uFqIyNH9n+wV4QQ0hMCqx2GJpPXrxslrKh4uOO/A3NzqI4tsqgDIxFC7Z1uYZ+h+KZ09s5yUN9Tw
7liZHnb/GsCMLtg1M3V+5nxY3Xl2TJZIyM2eI/4xqL5ph0L8zz0pgbSVTuWHaHYExieEEfhLgDIA
wpKjYuwv3P6WCgHL3cGeNZoSZ4V1iAjUoIa8eyqEU6HXb0Wy9PXPRzFoH7Ry55yr7mvb6/V/Qd6g
15eUPArfTTAkn9KgEmWGxmMQKbtrVz2LGmwsmGqVrZSTctdvA2ADxSNVgP99QjHgONTAtLHUCTaD
qPRponK+OtFS5BHA3348O464NEP+pIHwULIfu3MkQtNptF/ChkwhgGrCMjv+/DkPD3cQ/oJjiux1
d5/pzIKv+2k1FBecXTc5ftwFV7M52O66H+Y7rbYBsvAH9EfFpIveG1wAxLCmIgfWzCsONdcfyHHh
c6AIGvY6qbzCK00INo4aZt+L+5iK/669jFQQNhwFbihDCRZjDG7jhPLt3vEG3WSIrqTrPjJpn3WL
3Sla6JNe3PAhMjhlYei0dZTCfhchalzW0EJvd6hefCF+xlTmhEYKaxwSCjFDDx39sWERmILhTOoP
Pq+XIrhs2D3tpTVMmavDET0eewcpA/ed9U/cDggA8HlVdjHZapmtiLIWg3u7o0SPOiKNj8B+AUMy
aq41e0bXeYLpeNF+f6i831IabelZkaHR3FLXZfWZ5izLGwSKNlLJbj9SL7zo3qyxPo/fuj1nM6A4
Ncyt5UAoiNsSOwfyEsjlqgr37ouL8+S3Op5ONeLqd2/OVdR+OuShyCGcAgDZv64tjnY0fEnQ1NWU
lz641iRh0pYVweJu6Orpxd3xYeEDg1IbdgOAfCkjghNu+5fFQYQqHInHDRpp+AYKWbbrxZhoOrnC
DOJHEjNb+CyoMgM86Nl/87JojICdvALCvkwdx9CTj3rsaPOoM1GssfLTyLkx4hjU9WdusJUGBOK9
pTeZ4AwScamoHaOSjK/3t/sWv8wZbnqYIk+ZrLrWWVmYv+MBs/XHlyJ3u3uIYwpJpGSlXPbVmSjn
2bmUBvPANbKcnWcBIqP5vJX/nk765VNOMXKZBGUds2CFbG/gqOifRWl1Rfw5m+bPjpn5t80EImsc
MXqtCWy3DdzubO7y+o+GXX+S+zs+bg6wDSgqodRpOTOKJArd4bpsiBR7vt2KDnx0K33t9EeQS2sX
yjg+XpqAsj/Rh58WLGzi9wVXZTbnfYYnuOsqFoSAEiifw3UXKYowRcNwt4gw9xpcMHYPblWAMmmA
KJvRp8GfjfjMr4Dl3m4glQkNjEEAFKktU3CvztyvnULJe5ZQEoa62sC23zu1RMHAEbm49AQEDWjT
1vT2R7c6oSIB6E70u/Dz7dwMfWx6v0RdyN56z6l6sFzi6iadcnJ4K5fRj0YPCJmWO8q58quqTcCc
guOsXSsz2bQ49JYgQR7Fllkxc3tq+ZUHKLYsgBNDrSRdkcptN+uafecV4V/UUn5tIkcmDD0ReTQS
cvqWI2jDxngfBOpXKk7aO7BiEEQLUnIHIXRx/306fOJYXimuIVvF2xk+JP0+jH05JH7TRh/6SFxS
FFig9fo4K30eN0gESWJjokiiXAJjrFdebkCUxKn5u5TAh3k81s2941MSGetruUY2ob6fmxgWJbPA
oDwykr3WyLRDCTX+j3GCK4YWcOrgwPL5HgDo+GEQB+vS9lTfTtNJLj2BsMeuxGPtXwpSEvl6Aug1
gkth7XGsXCslI3EoIqC9m8Vib4qR/L+LKVQ2wNY+JOdkF0Zva0TqGbbwkIb0PKj/h2bvquWV3jXA
gk9u038+QTpxW4w54ZQj2xNA7JKWEPNDZJeWeHhjVWK8cyLL7iCWKZ/rucGr/4aS3WpHazw1pWiz
JFBIhkgPAab8QIOli5SLFWOjft/L1MqNk5eJEkG2/6zO9e0UUHq6acsfEBV4jImcIAS3q2SzTulc
0FSXdqlY9X/FLrNYlINlwBAPyd3qq4MwOQGjR0afzqIl+mbgIi1FhmTYgrbu8LfoOM50ZH4v5kWK
IjDvqtmaxpN9H3zsij7YrWuBrJGX+L77bJyKjESNwQKa1/7Vr9D+uZAp8e/EJkzkNzwe9AS2MXph
cc7EA5xlyTI+7ERFYxgpxsxm5yHckStGjXNYf0xijorys4FRh0Ej5Bqrji8vDIVsj3Z8XiyeUNdK
y94jZABnr23djDou5BTZFPsSH4uy8AZ84oGCHBMUQ4Ad5prMlC5d9wTskJzoHbteTQudmjvfpFZi
lV9e7BTqngUJKYDZmh45gHTjr0ADa6Ap5ctRfgLZe4jR2ABhRjdFb4c6UuA+zDs1Bs+R/zX9wG2s
ay34Yc5gzEyjQ8Fc4N/iwTBO1EUhn30uyVOVm0sfSIOln7mTzfhqxE4+Eb97B2ErGfgdOW28kMrH
Cz1pJCYtnzs1bD8Q4ESGKmJMs9zxPRLOz4y+Bko98i4YtuhFq3Svez/NGgfok8k/CDjOnYmpgnKd
vroLAHFsT4nYCDcaS74r260FY4IJS8c26Nmoxu7jmG8lOcpy6k/8D/VZtIiGhz//neF0KBE2D7Uk
MAq7wZxVKL4no57xKh1e/s6xER/lmWps99lcGNssrFuBtu1zz98h8HlIro0AEjulRaX5ElPhBc1q
XOxpF4XhyUgSmAq0hWOPPP0irrEbrqC4PqYyuHDL/cgKSyR2JXHafxtJWFR82dIoWAV6mfGDwdV7
DWJyT0KLg7kSnTIxgAE5tWtXVodL6OkD61NKwlx6Cq9FFhjAU3LF4aaFMxT5I2A7QKhpojoZeCfl
1whN/KvQfOcw9aykM9twqpbr9bHl514+IBhevKZCHHtwEFzZlnB4vXEBZFMVBtTrLcsyDmLKDdKC
YD65CB/1L++ocoswll8Cjjqj1qjsNldiWBl0lM9e9lzeynejbBHldJGwEOoJKEnK1F5aiZFScE2M
vmxdMriK7Dq+7DNiHoMasEXQTJcKFSDWaGpfVAR2CjcbIEcLGTiNXWxXGAXtynOx+4xrt2Pmuaaf
Za05TnR1NOx7CDbw+xeALixQPHm6l4DGtSFHUbuUTw7Qx13hTAtARklOxWxOg+qmgDn+s50XATBN
F3us0oKdVtCZDa19fykMdWg++D+lE0lKrW/EmueeUwWwzmWEjR++24I80IAdW5wZypz8pBdMGr3n
tndGugVGAh+Ivi5N4B0b3ZCmhIdcklhNaN+wh/D0Jfz4nI2CJ5fNGk1VuzlmPqTNduI4tGAtcXH/
ZaA14jEKuPwdX9GW4zHEp6Ps0l7BGG+KoqezYw4DvyHy1vrTovV92UVgAXvCgua4vwalJt42tL1w
uIWRFYjK7f1czqd344X3/2NGuCsEVxpjsi5r9iPF1xIftcLV2hmuVMf4irHt3vzNJ4ydhTRgFxD/
TSLIe7LtqV3bcCzdDPOzvWvpMwulegPeMEcmKavySSldZeZezCkOMIJgmDRbxS8mFSjbgHzIsx69
y2rDPQZoTFqnQ8xqMEBnVsukMDan2o5JqmYZTVMgHKTE+Fe+RxysStFLxHHACwGonkpRiUQZ4qn/
vVSemT3XVsnAyk4v9ijoCK+K/8E60cPZopo6OZrpOT2iZxHglQvINJctekBGO3G9Tyt+mJc7WwVh
Ce8z2KVvmP/X9qpMKyQF2uyX8i+EThEaE/mYya2LMAqBRHNGbac1RTuHlvmDmCqV1KZCSgiUxdyw
d/KJ0NW/LNquW1lNcZuu1yyA2PAcSlPj24v8aUqvJoobjqr//Sf9AEX8h+5r7lqknrENwe4ojBR0
QlanZXvkcozT/odV8q2cuJllvOM06wfAQWzutiJQBFveHFEjLwwJH1jUJvN7JaQpBlhhRLEE4N5O
zzOUUWL48jrMXNf9jeXmkC9Ts9bVf2tUgIT+qwX9O4n/XLlAvyf/jhAHnH3JZEcW1Qm0BWEw6ZRt
WKqSTTX2BbYC4O9j2S7/w9vsemItenIVVUYeEWbvnjnGPkFzEZwtvlbDXEJflxauTNtz8QWBKptX
wPScc2DKITQLxFyeQnjx3JFZXGk9x3hFDQER4Li+2I477/frehQZjPVA7brOSyhTi8dS+wu1Q6lf
dY8U3gpM9MupjqaZoeA2dEca9wp+i3DA1x5RLV0MMN9t/R5+VZ/rLu8vjvkpJZ2XpvWSprHcZWoz
C9rEADJy1shBmlqosSZycLr5sPy/fONoBkUkGY7FpXj21YCopHzWMAxa+z6Kvt8Vw19ZKZvJPtx6
1ekC1gU8skuHjuPj19eduO51UBWf7ug0G41YmK/j3eVp7WhYBilhh6EuuVOa05AuzNFkvVNENnsJ
d+bzQ3EmeDcfPuWNoLg9wt8v5paR3vgsqhguNMxBn1/NRQHgupOTlKXL3BqCFCvgjw9MFk1vjIcn
ySREI0jWKxYITZquECVN0+klvMBIeMfoE50RjzXrMUC0erhb7Nn/hkB/496BIh8D70N+OsOt/QWx
iYWw8aQXJ0Buh5+K9Grn7j6gGdJuBIby4I6VLZv7O6XDRvlCDmF65Ey8nCP+SgakUotIlm0cp80K
EI0vTHmUfPz2jTDpdfj5mNPphJ3TI8WAFslqapWYJY287NOf9QqMK2C+8bhCh0GEvkaawcekDopf
Rk/MF9DGLXqALbgnP4Poal/bv/AVjA1lgU3eamh+CVCHcNrhrUx6gu+kzGFLWnrt4xg1dffSb2JC
JgRq5FgLOntN8DWO5Qz5NzRAKgiCSsN+QmgpMz7Rb7jVOgmgFAWa8949SZTVaeVDfr7oIiz50uNv
cI005mCx4toR50+2Yey5bl1QGsoec1eAhx61LD5q1EEVEk9ZKDCmOgyEKPgWDiunLRUTvJd8a+DX
LpxfHdUA2VwwAh26SwBMaaQOpIiBij1fHSESMxcHhO2CKYMmaJTleykZWcT5MjuvcjnbZcZ9mG7n
DoJfv+BDcqNZOLg+lCmgPFJFAGJRDpT/58Oc4BVNFE2y0E+T4Ulxs9v2436DCY6bXdZjk6N7ASaJ
kqguspPZave2am16wyP1454KF48ZWrQtDJX2AQ3C+BwLbrW5GecEbrWoKG+HQsgR8b3gd/Wf8VU9
OMUIEcLzU09yveOuQGf38ZwTwfrBGIIQ9Gv7NLoG8fFx/2dyUs0DsojFPQaFvFyhSITrTi4Lw90Y
F3lyFLgnBMi5ugRVXLjr95Muh9COAGr0IVV1Q1yiYJZDMEA7lAjPNm2OIljde1jzBCkqCvJT++Se
uEMM7LHRqYElpJ1XKAQzz3jvoEJBq+GSGk15SWG/7UHffYDTjXGEfu/pIX18y20h96v+BJmbYCGz
MGRfVLABLQrgutsbdBuF9JVUJsZ7M48UutWMsy+Kk5hktLVjadjpY3NOc6AW+Qd4Af6zqSSqkk+T
Us7CnBTGd0oQXyUym/74sXRPupj0pEvuVO2x3LXN1Tc0/pWyuN1DYnXxtl/b7hkoBMnPe1Vu/NO6
CRliZlz7ABh+QflbzfNexC4cjf4j/COVuT3pGmrFwfmQklgC1T73HCqdG/Jdeoz6GCbjBVPt6dkF
9ipnbqfsy2ci1acws48UlUoT0i1YmnOsG5H/xr0foT4XyTfzW9oNhCudbN8UujfLwdXAibI4St0a
8g1xo3hvO6Dqn4GLTjRUbtVNPqlXW4n/Nn/kufMuOcvBa1gTYTdfERahsiZu1qKRgl8OBz/8Xq9f
NyN6pNo08L9CkuD7euOCjAhHmhGZ84FN/R+kY8UmT9gl8gsvggT34Vk9dv55ma6JSBdYMX26JDTF
KcKJwVMXpVHuW9FPLGCC18/eLJJZzsoH8TrYhfphURph3e9j849EpiX9lNooZeNtOwhFfUh9ex1l
nnlyMgmGxFPUXYY+EpmAE+TQnNfr9nTu/DngXCNGJl4rzTE6Pl/6pkCbqosod3YfkrLKPzOwTDnS
wHkpylKFxUqJTJ0AAy9YpuR+8Hfb8uVcFcdpxBJOB0VfXTUXaGqZ9DnB+AFwgFHy00OG8JHOIPpE
imCoBbchkFXKFxdD/Jza7cKLZpHb9NxHNSpLTBtVCGks6s0LoX5L6YVosWG1bnQnLvXOgQ05sTqH
wI/dqXlk7z57tPksOxkuFmKPqnlaszSNNYBh1oNKGF7b1H25pfJcUko4XPg7D5fCBWk4EYJOkMsr
ppU5q+p9UolEVFNQOgyrgAy8diz4Vb3QHRIZ9YV3B4pcdFgjjl2jcNv/U33qgvWJ1baXq/HFhhDo
4HIsWtKWgM0cFKE1VO9ONHAEPRnoZZ4L+5840avEmAaaFWei+/+Gh8wV2OvtmsLaskxNit/dsho8
dJ73blm/ax7sH/Ft8AFgNQlaj8cs/CEWpYWeqweo28kBGWQS+iBCRgyk6HSAZozOle47WqInMTTu
ie9W8ofI1MaI42Rmoc7M4057wmC+jNTOjCAWUDVSoWXjqR6gOW7JQUIM0CnSr1/1DdfzseCwEvM6
9VHkcSWAsdO+oNuu24vbr2/wEMWqACz2sdbmFffddkyLe51lqgJZsRsFnvGH5NAqjwirhLyu8vDB
BEwfZZ4k5gF3CsiotKwqG93b1P2euGhSIJE5Fu0ZppVOX7M9b/0gaMjfR96Eei3j0n1KQvqJ4h6y
DPwWrIVCUXRhmBfX8LWjDXiWtnheG2KmyfzgYFBv6tH89ZeBx/xX1SIYdz9i1kY1UaYDkcqTUI5U
c9Owc5eAPhVVv1bW0NCNbKaGttOKvhzXO7Vn9Cm0Gpbnq6mj5i3E5jGWM0l0t6N+kc5LUpjRNjgb
ogf/1zbgMa3CyMNu4ihYsSpEvVcwSJO0f2PSMV8RzIJ1V0S+N3b4Xkv6dCwChUh5yMxEMq7PY6uX
zdvB8pBJxZfSNPT3TZiQC14Zu5VWlEGZmPlsu87gjSfdQ/tauwIkVjFmJHnOPnwlkPh28LQXBONx
JggK6UvEOI7yFWETOz3rqOtSdoomLYWtL+OHT8sXayJc0vEMyG2j8mgCtq/Ojok2ueFcCJD9wwBa
Mt0nM2h5aDua3SkQ5stNO7iSEYEiibiw7cO3FbRc2PNaCd6Z1qWBwaUsODzddnMTVKActgNGdz69
cvi3lIlSScTG/bOcRxGIMSAmtADK064wt5+ltZRwGSady0YTMu6V9LhBMgPojIY2Pshgdx9O/0H9
1ui0jiZ+kaV3Q0/VkHecx2XfBDG1hh9XfN801BE0KRvdqk62XtcgEzSabs3VL3HqdfhEz3n6w8rW
4s7pWr4tmdJQzeFiN6Z7kwTZfeabq82ZoDRD89ajkMNCkEnWpM8D3+IfyMl0BWzMdjtEKnE6h7eU
fSZ5itdoi7J4vmhqDmTCjvM/B6If/qMUhg+BDvRAFnVN5DHdIZKJbCzHJyFD3cJZSw91jimtYCea
LviGibTkHPWEeQT1LjtL5O4zh8uqNMeRMWZWEi9ab2Lx8IoC1zYTTARfVrf0cxzGHYCSyacgTgQ7
kPxn8VxzHpvRqpOEAdewj/76AeblInXX/8B7/7RoVwfJOd4AkMjf8VjNnTqQnD52/iWpn2algCcl
Mjlp8v4UsFsGQ3x6VeYvc81Pb/t/vex+nY0o1AE4kgibN9J9IK/fWUnOOunSu6Dfzv6DzkCs5OIW
gEwBpxsAvM08q4TEt/lsYPfcyIB3KwqYeOusKvlWIZ8bVcLcln2MHnFjmqFHyUcN/KnAkzQ1ZNBK
OsXzOcc5LKDY9RJVUOb3DBHcCFTz7NtZ1qGZoKWld2o8beJmJbS2/9mXK7ITop50uKlI1Hm60GMO
AYOIS4nh3JIlY3SvkgftuTSpsQ/+9zV8EQWzxsuarl+yTqCf/Sb5FwA+FQq5UiMoxYU9UL1csB/V
NRdTvCeXpiYeKUFfBMBbDZnqmyfR2B+0A16iJF9zXb3ggLnK1xgpL+GXzgYv2WMcLRjOdltVVQyZ
kjOJR6iOTXqDorqPSBd1GpMOUOORc95gfNNGsInW+gM01Q9T6Jo8PeYbMgO9TF9ZrWnyu/ZW/t8K
CfgPInmRE8ogaPD6slTgljweWSMdVhQCSVyrbae50smbYuRjxwqPVT8FVW//grzCHJplcvFu/O+b
f3r6YJtWtqhEgU0G5fcRU+SfPZVOwU821O+o8rpWTjaB02E8Pop1QfuOHghjHEHQY4ipG+RAIey+
ow4yQZBlA+24vBh/ymtETIYXMgp8J+OUF3/0ADff918XJEQaYuyWEzCvccsv/jssMa7yQmyIFj9K
45/RYrY1uKYYt/iyY7gp66LJx1auuUBHJUslJ5Zh04wbRhmdl8CLYIx14t4WmZ5RvT/ZC9MNGm1V
s14xbe/DpKTX2gOak/nffXUOFRTYBlFiBhF9RrE69DnDET5MOWBJYRnE6JeBWgQtTrUKWs7fFOGA
eqlW9nx9Iw1vopu4bcILUwJCLkNdvkjtaWVln+InZQpxwaXsXKUAq1x00JvnawYtqQRaCaLUYalu
aw+aMED6ILHZBPXUvzSNIOmgesYUscV2hHSaRCQRCqpeiU3RXD/drnx/gGrjhkzh6MONIednnYRa
P5fEajV4/rewxQzkreezsAjbNmCYHMuSG7k+LiF43/W6Szj3vMxhehVqovqMUHc66mDqgQsTU5tX
qV+5TwvnR9SchKqcfbp/umay0OvWxiWbQ71HCOZN/yNLjfxW1vgbOa+9PVtHIAk+BwYB0k7IW3w4
Fivw8ogHAqZwRSO6QJXYTPt0+guga/VSoGnJ1Prwuri1rIK+Ss6apYqq5H8l0S62lmWPVd+nOl4U
VMLEMubgEK4nk4bpMd0tMDC0tVioNSwiG1Wys9G0uyNHN2pXYP5eHCGhd4sHwW3LxMQ0g4qgLgbg
r8xwj8HpS4Ft/U5g28db0Vg0JBxxd9WDzVnUNZDzRq9qWe7Sj4UXYE8klOATTufoRglXFwvu31b7
r3vbhGnz1kj0NTkQtf07eS23ywrft6rl81Dy8ug66I2V19zJkhVsHOm642VKkckGAxwktyD5UrEv
Agrq4uW2/lk5VLoH2n8bvyQOj6jdaBsAZXbdhyNhmpoGwgQPBm4W+8I6vF2pBMWFiwDWGuwo34Tm
NJa+JHlApsWGdhC/VbgLtD+bRtFcV4M3JcLLrb+Z8rmfMa+r13axPGzKXxaXsQm5ooaSActBDt21
+ExMd/TM+hYF2bXQ8hRsLID2m/53dpgz+3OmGDQbtiCKP8zxXBISSYOjNOju1cQpdAOW48zlzISJ
9r7hqhqE7ZjuWNhL2R1R4kGGE5LiVRUN/AFQWjZ4Jb3vN0ek+FF+Hb7un+k08Q6ORT8phChMtj4m
Eh5BP3FwsI9XimJF+/Yheg+MQvK1+kojvdNWtVdUa0Yt+KxTaaFakN7YSNDis+TIt5DNTaQUp8py
6ESRlX4XsNroJHSHbI+66sPms3uPK57qAcc954y6c84QM2fDQqy+ghNACg79fSxCLE/6Wrs/QJye
w5KAx8udS6iHhwyOOG6qVOI2ESDy3V3GoUEkjZmr41cpyCEqnv+n2//gYdAQ1vzgvfxkGgnoQuig
Dg5dC9s9if3ihmMiYafW0eXV1CJ9RqingzVsJfK9Vjfx01JuRw3Yv12zlkZr/QobNS3XZvZBC8vm
iUO/S/DVz37ZylvhhkBKHIJlXUg3CSYYrIvxbM0u2TACUSQKeDyPto5sgbmFL9Ny01uyFbde39AW
I6/YvYmKfbv7Zix/tIsxM6ijJRRmLy2sL7q96Qlz+E9HKaLwERxRHep1l96/egpcy6vCqNQxe7sZ
FSQi1lzt0E9/9Yt71EBcPArGmZfhozVGOe7Eo7s9U8H7TiEOJfU2g3v8GjlePiB5Kx53ALSkI0Fs
T1aAwk5HoBiMTMxLk6ITZN6j3w0SJRsgjqXiIb8t+vYuBM5H+Lxn/f8uritdD+Ru+j9xhVJaZdZk
UWWKs/yPqGk/ypPpxSRKcl8EsL8dSKoqmpHhqz+2KMTStN6iWFcucaGeVu5rPa0wt5cbKmBXmHpl
VWFufuc9VBizisxnJUyGSIPdyMe6YbLpPAXhg1vZUxUlGSfDQLph7zb3hzc8plluQk0U/tX54Q3n
DEYXX3UJ1EwoQzyLngGbCSTSizh1wUseyXLlJURtZvqzodspKaGoAmgyiUHTS3MmGDdfZ2VP0Mo/
ED/Z3xP/0GbSO+U0d4EYT5sh+JVKJfQ1WV94SCjMxo345ZdOnYwvyK4qtpLi3l6JzLSzW1+xTn5r
PEc41J9qtMpDM5Sos2qY5xTdpL8oSQntLRT4wXqqvhfL8fRYvrldT4muer3tb3hKTLW7bg2iOYYV
RiSbBvJ5hDDkGdRPIxd2CqtkD97yE4Gw85FLhlgcQ4Hz9B9rMkpQRJxLruE1vzn/pXRfKSwZ+564
0TNxklUMPL49UD7Z6N+uAJDtxE9zmKHkFLRDOUuH1mvmCz1pCaWSKmIK32rJvWlwnbTbKnoe6sHo
voCuNpzZypSzmVpH0bGkFa8dmrtBm7cz3hR4m932xDuHpLhoVp/7FzVzUutuWzSLZLxvzmmEwbZF
B9m/yowIsqvNjEgro8Lhu6OXl3hiJCD59FIRV+1Us5tPnNamK6ZNZP8t5YVFpy8z2xsnReTalUui
fYl5izx+Onq7dakO+HPx6o2t5p5jNPjRmEktqY3vU3mo2RMQlzNnxd6atU3A/1qzONTTQzBpb5iy
UQvYgwAVFvN18pacjI97GOEjGcWwQ1+B9L0XASLvRl8a9i+pHA8akGrl562369HzzxDbiw9iadZ1
rOIrSxFCAVpDRc69aTOL71kn5UOEkthLwGgeCYpBaPsbRMrM+4gbZA/lWHr0X9zukpbQH8l7oMT+
sR62YXFKS++Pj+ySdH0ngFJmpHlnwmTIb46Ouf1gJswuP0QFksxBHQT9aDEzkeFNnzDneKCmvYQ7
kwcTymJb02OavRUarul3smj8RjxCCU1U+bjRi6c+2V4nQmmzP8UOe8rJGYxUDsSFKuy01AY/3YeA
gOHVKkie9hA6yYfuW3Jr7fbDChQ5828DwgP+ywz3mKn79Sdg/J3WrfOGZAHJ+cuiNh+tMCLJTHo+
oQZC7zYikt6GqiQ4vYuDjre+Yxp1zbOm+OMEHCBYZzooaxkhPNnvVIvGRGTtXaLXK7596mAJXlYM
XDl8EpQog2us5Q5IU3OweIvx/b2aniXX4TQSITyF2goyOknwMznzEsHLY32y5v135nvN91lYAsr1
bqQab/WSiijIZZ5yxZ5hJ37fSfg6/m2Uzv/4H/lmXDhk6nmFhwS0zTkUxS75O9E5wgcbsAcDxvVr
SUhUHZf3Sxx79sTwOf4eSEyslhLKZyKYxy8BZsD8FLmM28SAsbuSPCLovvKJEZqYQDhrTI+nm1NE
O6/UNRHIOcPKpGUp0c/PFvzoxO07ld4TuCxE/HOA8wp3gyLpp4QlzUDHXwd1NzYZu97KsLIt7jyX
RH76lM17GiDQU5zn8O8okuaZ7XxXJFgFyS2C396uMvHIrXD2p3g4/xtWvSjp6pH1QiJRQWdnV3I7
MkPAgNJKWr3NNEEHCFnTvuMmmKZN8T+HocZrrIZwZ0ceoHiC+wWwxgXj8vlBrdL8hAMF19hBhmXV
nhDdCZP1JiwwfxydtdFxJYRQ1EWAl9G44RiRI4BmmnHodMxU1VFEKmqC3F0umaFexFbp+3o/qCUD
F/K6UU9zoqd1fIkwABUCOhiMzYcvaVWzsUdKLxvjG3FQBOBE1I6eGUcZoRFh+jSmRs6LPAwh6G8i
+FHmIWbwYw0WfQ0dxJ2oqyA1jiscb0Wo+WzSSNuk0B15YeHQI9QEc/EyI8foi0eG8IKyfG/aTsiV
FVBWtKaMfaFHaPTJjESd4ZGdcX6wEalmu0cftJVCxhGoqsNX1OhD68XfXtbY5vhzTQY5FYEGutMQ
X2yF9NiQzsnfMlcVAqxYb1pA3jVqE/5BmRshlnfW2QZwlsjwLqRh5CYjo2m5otuAVrY6MM6QuJyc
BelLGboZUYMnF11lI9DLC9BrRK5rEgyb2IqNndYIk0gG+O00yZWop7YHxwBDMhW8uBWc+ebSShwk
TYB5fSBKfMYEJ7Em+olyu4tKhHITLsFiUP9rraBbs3sRZUJZeZoNUC1g3SSIAf3O8lI4XtHFrrVT
Zid4e70jDK3n9DB0FI1zDyT+hXOoeOjTAtOKZ0uXXlfYkInN9ReDwzHwNBVLYn7s55Y0uOfmSbBg
327bCYEfAIUxfSBmjf6BBOq2Y0zUxt2CCGEzaMx5PFRG2zy1yxVJLqrS3erbkJDNbXK7zqhowpRx
us/CeSrtAPdyvKnlH1V5Ca/XNESXvxLV4c+wyrOrMZOdlnEz8qN05D7MaMK2zxFuhJ9PzYlt21Je
zsc4j+yUHhgDQLuaCI6sL+fn5DFB3pBCPaefRpFH0zKrO1KoOWEVPkAin/W0s6frO+w15Tt3bF7m
/cG5MNM1IXPbaEtdef5RsgViljyXC95ZggnzoacSxGXrFtf52yc1Uwh1QXYANBHwBsjP5FVY48LN
xvrmLCobcUsdeYik+SubGCY2hKjUw0mGHJRAziaVOavQS8PlNH34RMcT1jIVAfAtcUnH/EeoQ5k+
B0NxpqRW7cPv6pWLYh+BpW8BBzFIwVT7W6i2TT/CK7S6ptPV+VxncPjUAffvraRAI1hR5AuRF4Wk
aF/Vslstn9QeiHMr66AOiEdhKJ36m/LalNtBrTyXltPf4aLMaOXPX2R1nNtO+ZxdbLPSQXT9bY9n
jsTf2ej1OAxXUJhBeypl8DOFwPRNrvx7QqHeuPsIVi10WUSD+phq5uDtexjjOsYeb1cKcXYmp/Gx
klpIJew4E9YTP5/LoVfQGsJZIFQw8b48GP0T2QThaH8aXJUwYq9/sAmPiW+x1IDgLMfXQWjPkOEg
rM6OvzIJ2v4d7nOXlmU+d7S74biFWevQBKNAIE6C+J6LcB0gmP4cuuhH45CNXUJKK2q5/9jN8Jmq
iXg06Zub0Ri3KWXinjMQEAz5MgMiLy5oilu3nBWffQW4ZymB+bfcGnJtMzDVDkkGeLwR8HJMOfKO
nbXzbUhQIqUafEXVAXeQ4rsywb1MtcuWXjG4dr35F/9MkIG7CcQWmHKuRDXRb9Yudm31qZwz3sBs
eaYwvB30grsNagam6nz9s11nyNPTScnZNxIHJY7ilFPKQFzit7OSFtj3Gi/u0XIzMYzlmfpaqm4W
qtp4+X5PV/PL7oFR3ZDk5suthaZX/cl0f/ujkvgb3IlFduo5zrYtylokgKP8G6uuA8Co7BnUBIJ9
juqtagzsOxATLnoIZOc+Q4uecN9H1w5P1Fm0sn3op1OPO9b8YsSigXEkFbKFLVRHtfNMpnBGxeAf
jtdS8ZUD8pgewjsXqeejoko0ZCbVZL+TOzC3EImLufjFL1srOIq3iFpazH8203hgQyN6ykffOo/r
y9jeHIs4Lg81a4g9shsSwlCwEdh+e8fWEuOkTpoS8/xLFe5tQ3NUCIUPQ6RrDmiyA6TFh934kzSo
HVsmyQFuOhwRDX18B14jV/M+JWVd30jGvfiXbe4RQU/d+za2sfzBP0jpYpAjVE29MUibTVV4nhKq
RBehP1dqsMFcsLMvOMXDH/IKEDLRcZkXuMCw/D08dYKd9x5C2sf5Hlkq52nOYjKbxpLUnF/Cne67
YZRwQtCGhNopbi6XdfgGA03FJGvlhpV8/wF3+4v5YZzJef9gluMmNEXh8SkQJU1TZ+EaWQyAP9dT
VZ+fANmBtpQ5/iPbF30GZE65GjKiXxgoTrJSIQM1O41rRc3YE5KC2BPUTL/UnxMfmHxC8iZvzXuS
bIXyYxPba+9N6ghuYOpz0YMdVIb8ABfN01N1WWOrzRADSOTsNOAxsP2POZ8g9wU9gXmCd20XU4YC
kan6UYUHGim5XEAFJr4PSAMR9wCMQEtLRnvYy16o/6e6Z5xOTtPe8VWZMwW/k+EFPfSMrfd/rXzz
3Q9RiXtAGtHvmotKgXaqiIUvZZ89/EEJGyQCDQNgPXl1tKugOfERSrQrWgMSULD1xnQAv0huq7YP
xXMSaSaZZhNzGO89tnQ5VKe4Mf8j7NsilB+Tbr63j9caPqbEh7pgpT0QzbuGLvKcLQTpXhOQoM9T
KR53MaNi2GaINKGRpIXWTJi9eFN/VBCPkt+MUqvMWGoNvykrbb8NDhQ6eUmHxDbNyISOEInJK3qM
zzcn3Ye5downprNrCx/oOqmeghIZIGHojlj/mreUg1KfDvMb8p8k5B8R6CfKxJid/7d1Y91Qq5+D
yi0iSbbJC9c+5GW1nZv7LMORs2AT831+idKy7KaDjMfBOcWGPR/zrbpwQMnFT/u4Qu0ptK/ZyJb9
TQIv9glYOfXxXa9N+RuA2bOZBzfPTB/bwLLSipwfC1C20bUfntozzBdB01HJVpIfLVsd+B5phE5T
3pg3u8EjjlXMg7fYXrV+k6E+B+jy0wxlbv7RjLwH+oYvEvfWk1TrCCAQz4ijzzGsiKnTqJ2NJqJH
ybb2dL7aChU8+PRUY02DgZBUvYlNdJs2oBgV5nMbvMCrMwewKyPaHt2lEcnYYK7bKe6/BQ9/CObz
eAsasPNlu4HURW15SG6wFYuOIXvf3iaSmM1Aj4TLLmVAl3P0ZPiXAyyraMO59d6T0Gqjh2FmrrrR
jFAs2aBhzYcqyCIVzran1UrLsDiaxZJOmggi5AJpTrO+0oljA992vNpiRVZfSf8enhDsKGguSd94
4m11e2X0yl8VNrk5ciBi4/0GoHwUobRZq5YXz5QR3qkdx6Kk/GViHX0kE6IwkIHLi4qCh4PYc66D
9GcUspJhsAXYebbSsEGjefij0zpBagebyiaN95JhAalPdaRnfHYYBf/+jEmaVjX5t3pU1hhueD2G
R2pfnDsW1SsXFhl2Gk8sldX3U+TL0GYnQORhozcK/+frTopnRar7kze1knw+nVPWLPBiW8zJ0WXP
ihvl2TyPX3fTUErMmT0FENIw8HWy91hXN4Dc6U4AWJZGQKnt72ALogD3aCNt9yF3foSOr4/4PncF
vMYQSziR64Nr9zWwMjL8bjePtfUKqcjYyMvpQzgd2XVuRsY8Icw3N0XVZCPRJZS3slZZwSgtrt1I
oY19nRXCGF9RxubWGR9Bi8ThRboFjOEWCaY5Pa8KlvFLqBzwhx7sFszP3N0fxjbnXeZcaKm5y5WS
JzRd/wOpTWa6eZT63gxjdQgCYLfvA/+15vCi/Np9UnKDT6LOEhkgZGs+muY0DIATUbjxLjpEPb7h
dD406gDLZVMj9I4YiDp/CHWGWo0RpeScAdTRD14p3G1FCnSrHIMFPiOqAhaBZBnUttFQfqD3gaO6
iZ7EcVV9QGN1r8ew/QF2MDG566ztco20JdI2BRZbu8U3KUAKCAZ+s4a4UzEpFG75v3ovRt0yuyMp
+xZdDeLwa/3+iIOgPxrkwLN3g8rA+XZw9KJ8UEDTbiFld3SeKLJhQaxURi66ZY0+ks+kcsSyWIEj
DQ+Zi0PpxBlkGHqaDMdrnn55JdYaDL4SymZuTI1E7ILA+vjpTwA6SbMPpgUn4mp6rqUYtQVIEA6R
/uTZLn8JmXDBsvYck86h2O+oNKSzVAulLM7gpiuytwiMCIW1JwQw0dbKZHY0reEQMgi8Whu4VvvU
aYMjvs7OYR7VezslOCQWMZ1xjgr2mnRDxTwSlJ4pZvZjXHm89g1OgbwzvlTj2pZuXluO7UNmkttl
XGwb/s+y481ihDxQrLmAzP0R0egMDUgiWjh8ZGbROwB6x7690DBN97G68H+/JHSLj4oxLVTNGghs
reGdgjZXolC9vPi8F8Vbc4+TtJPWAwn6nImgB6e6OW/NylYPhTgl7H7hMZHD40uprstbBvksM4JF
45AFFmaF34vKnHq/M0iMO48F+f9BG1Q4zODUKGInesdtrY0hxrHNlroXX7TUtSLrzmpFU/Cm+V8V
+xMXFP31T/5RiCeut0xQyg1nM2VV9pRjqwIVXOWOgfoEgevc6PH9oKUd6UcDKQQMGGpWmWaDdFk5
uzGYCjy5DP110tylhgBntWyCXTVTSiR73ShAJN/rXvwwUT0b7Bxy4Ln5RRnv/Ax+Io/U+hfyXifi
uLiBgUf01k/npJ5l07Agf4ifSRcNnotOq0AoI4xiXJN1sZInwZnCK0NxqjmURnglVFLpOAAJ1Zaz
hsoP1Oh60h846XyP5nQA8lVWu9907ewLy1ODYuVftZL+Sd6XpSAceKHQFI/BoC0wxlR1pAT0PJ4k
GDJtJeRwt7GF2JWy+/IgHcVKqMBxE7AsKJNrT294QNieD4w4jC8Z6Fz6yZehLgmkDQw3kwzgU8Ez
bAQCue/1f/c55LyyjHT/O9gTVc4VEWCq4afUdNii2/OPk4v1bVTTl1q4teSptbRjr/43E7JFT9ff
/ZX0TAEV3elFUa1xcJrmAOqisJVoYPqcc3PbIe3c6BcQwP+N3U/nL6nu0JFBH+D5Dr70gs92pddR
+0iubGy2x4FP9YjAVwfP3UK3T9UGDefyt8R1notzLXk0qUV7/I7R8f4rxV26C1qOT/3zUw7vJ2uM
WNxtC1xI58IZ4OX/VhOifN+35yiPM18Uzr4Mjsrw3tOo6TDpDPPsAuXQBV8Y30qqojIpq9oStjpK
2YS7BychMgxQRfZHcjot2KnTHaksnQ7tezk05RCcrwoz+Vy92o8AOZERH7NjQqabQxo0hAlt/WSy
bryl6vD1q4CGcoWPEvYwgPbjhTeC37gCOf2tknCTlUxhdSeKothcSIi729a6jthiz5i5VNX18Hh2
SRgQjh/RDyf0MtfP3C+M5/kLucyr/d/JT2xGQAcyhDFEcb0+sVff8/jptv8qE6QFMYGK+pklTWBO
g84zOdgG39fHMTHTiKZEHyEJhsB0uA+v6sorR1fCoxM+3H0YeP0dBFZh+UEQvKTp7eBLWFbp6X7i
m7zyEbDbLQ8ivEt5v22P0Ptkda9eXRGd6gnwudnfuYCsp88DpeRUT5/Ff8umlkh8xURLjzU1DRIa
vW/JBh9nCwbydACS/8/NSnNDM+FHEdzr1PvhuYzV7ZLiQdvTRVLI0hYt7+u9ZbhUd+x/tyumK5jt
PAW/LXvSw55dps5Qrl9ubQ9My4IAsk970pJGreWhrYTHvMcAItka2LFDvegwQV/npvE+gQmC7zJc
wGDShk9S28fx7xGm3NpXs3YdL/l6FDr2/0uIdgxgj7Q/a7d2Wx65XUf5gObHqQy2nazEiDYGpgPj
9S3eA2/iEDgTLVtjb3kStBektV0C9j1lD/tyCFYcBb0zyHXWz7TJawRbx3JX20/uVZ8o6SP6zuBX
UouC6L4lQdphQigf30qv43aF5kVSCouG4Q6ksOmViAJUqMsjf0yaMAMfWtcesv5IhejK7xA2F9AU
cXwmTyBes4klu+8nOvdQV46uUifKNXxR3eSUnomyfUg78sgHac0Zn8HiW5cweeweZprKwjRBDvO9
P8wNte0LixCGRuzLUnBEfWvSSNpIUfvtLsRF4I42z8MoxvV0/z7aoF8UU6joUNjZtuSxClmIFzqH
/TFZ+WWiO9HbBxlrPKTctoMoOencXDOgj0sNY2NpBq2tTEmBwxXmy+rf5yet6wMx2CdfheTQueJX
N4VRKeoS5UDTuRlNU/jozdIuYFSN7NQuYkqnI2ugFHAFivLQDNa320isnjyJk8D7PGOQtt/BLIC3
GBhW71VWM4ccgIPIriwTJ4D4/AbFHMPdZ8e8rlRD/NIhKvK80e1Dv62jC4Sjr9QHk1pw0DapqGlP
l0kzAJVnpw1ImF6zKLvfhdbyO1KmkacO6Vx/sTOtYnYZ0lGACQDxDA5YbrznMWm0GD6gquF6y1NP
6UCg9io4joByKctVmgib9otzY0VyWcQsGnl0mXOJDKpD8Qmsh7Oyllr84/Uz/xHcomes20IoVIuz
TDCwrEz/aigveLaaIhHdRE9K3I5WVKK+tLZyFIUmXTTpewr5EjxwhdeJA5GSk87z4uf8qCuliQWP
Hn3zewB19+8E5shXzwlopY1KOY5kcHcilDt7IEUKjULrCSYZBOMfJbbkQX6C0ce5tzB+zV+5zzSc
pkMg0J6mt1aRJ8fErSOBDCpKI45tBwRN1cYZ2KJSzHmSiSARf5VJCGY1SDYIJ9Kru56nDE3ZGhtt
zfkAs5GE8MRDbAXUmW+xqbqVPbSN2Bey6Q2X0Vq4AyBECWglYq+aAWmpPUWErkiP2k1iSN7YPRW+
IH55JgJNm4pJA3kbkxJz87QI/DkvC/N+TRrUCWIWjerCH4VXksj+oEosNTLvmDKo4bWJHGZ85Ump
H5C/oSG/rzLW2Apz9oTzr59SEj2Wj/CO5c9qhDeKQqAKOOqu7Cr9aQmS5TFRMKuLLf/eqP3H5IeW
sJyJebrOlYEZlvimEGFX14JskV2xA+zTJZw9posG6uUc+QncLU6im8sMe3J4DrCId//omDWx0kWE
mwV5hJYSLmTHspYtNmBNwYc0AFHWvX3JpeKVbHKcnUOR2MGICFYSnzwnUFkEiEq5IogLLcFH4FaB
IJbuvRvi8MJznoRNx+DxIPwR+EZ3vXW0csu+C/PToCT0YmIgTUYQcRYdK8GwIqrZwmgKJrjxV4HB
OYPTyndDdbT4LtYN9Ufbu+FjvQsyaT40u9COee6pAn72QepQJbUQSHne4NYuj06YmS5Gltlu4ye8
Fj3qRPiFo+FP6Raz9jL/kVxTaiCNkibMMI/9RZnE260bWVddUstqn1MzRgoH+Qr+NtgGkTVqSzsw
fYzXpl3eVAb4HSUuYOVVwh1uIbbvT7+BbW/6ZLXxad+Lt7t5nlxDRxLt87hjxNm0ymBFhgcfqu0o
Xej8rLzurQ0PZ/hu+W0BfVNPtCG5gVbFOBqSfHTIzMcyBBt0xDYlaThlLoozwqAhVMSwAyIUuzz3
OSwzja3+CsDSVAy5hLjzjT3TUkpoSh8wBpCdqMkBc9y9YbEEQsDJQpPobV+NzCCnXQCqwAJt9p+W
tzyPplVpqplYB9qOTtzDsoS2bbIsoWnsmBtTLeilrOXA6e+rj+SsR/1LJXeY8DydDCh1jslxlh/z
BaY+SRsfZV6TQKyufuX3CL323ZGS+4YAVqAdmsQcUOnE/N5NnDLVk/Wu9aVjnZUhswFENcJklqfH
u/DMBvzdrUeYiHyXqkXhaizCq1YRmazD0zIPhiiuKLscg21SI/YRrfYbx4RVTQg22613uPQLrjkH
eeFvDfaezhf9ruior+Wodz3BPU+cSSie3xAmCKB09upvfJO8dV+vlZgrh4aHSdxB77HIyi3PBVtn
562WID6nsGQhS7F+BH1HK0JUxDlVo/GwFtVlJruXcxvW+Qs7w1zjHXKTzMDoEJMWTWK1hLjnz6Qj
VZUec4oT83vC0IUI4ZISpaBVIWX/yxm8rkF2mvtgvr1zmg9DXLcYLJpAwhL9tBt1W9Xx1lMCvFrK
ZwX5qnBXEnACw3EYIaDuqkIvgGbJmhJFC4UeM1YeJFFQa/XWuKrH/5cIrTiFJc8I9T7s2QZ40wXr
Gho9WFlGzpEuboKhZ4g3HmVjhFrXgEcRNLk6eiZz7oJ9RpPE08kh28kdvAUA66KV68MYEFjAt931
JciR8iEtVg6aeaExJdh63XZB7KdLWNzTfPFiUVDDgl+lMtRTE0bWqySwUrrLV2WlHVyBzvcptBRj
+hgzhpGkGfvIUFcuwVQ9gdU6MZhG7b7m4bPXflnvw4GMMpKuqGnBn7po4dHiFmpyNtzCM91DH3sI
W7NQE5qe1NwohANrpTsNLV9WwdPBbCElZusZusbo4zQRbxeu+7wrL1uj4H0cxzqcL5I5ERlgGZyd
dJlXRQ3Rt5XDtvdM2VZZiw5zBjkGvB5/Mjqm3Bfzqri468PjNpBEHE7BbaDHydmjz8fP7OzPALg6
XlsaSheFfPCUqDvxd3lykfFTb7aqOVVPr2TOmpVIqqeGCG1kR9+drreUnyMfYIvDzE08hYEravrO
9I5/KMs/BhVl6MHEF51fa21ecjEJ8kaX6lePQ6ANCinjmyuJwTUpmIfa28MHWYl+zQLx6eqP/Jr4
sTWEAF3aoJvHpJCnDrjpHShLJAE3XxZsZ1k+I5CMu2SibAouh4nMdoiFsTVYmSkYUkD6k9M4skCK
cVKz5idiPlee4S6san2TARGzUmUXT5syeXKJOlA51NGpED0e9JYMgczDvJiRBOepJES/vUskwaBM
/VVW32bv5+hyU/n5tFQIzBNI/ITn9vcFeO64OstmagZ0h0k1V5kCnlY8KEmjWqOWP9wodTBf12L0
/RQhurXWK98Bn+75SrqtLEfsY1s5VtENQ8O91Rq/XRZRe2ynSa6cJ+mLJAACs/lx4X28VDAv/jvZ
OcLP4kHA7fsZRsn2WJoiEG2Uy+4pTMuarcXRJKceP48CUD9jM+RLMNweyrJD7IV1G6YBBNL9/Bgf
x1KGirE0/TKXRhCY/5uNnfJgBiMo1cSXcuzQdqPmaiPuzCC5BdQK7wrTGosWnBRanVaKt/UPdeQG
eZepe1Q47tVE3abo5i9eNjoZZFRdR4i9/LFGmgdfRJQEIMGjOu/1GZckD2XtEtGoMATgqwNkiOsN
AkyveyJ5XMa3OZPzMzxfQRvXZnKGtHfzBnQZ5nJtKonXxTZlHRPSMck+nysRgi53e+eoFPaTE1TL
BaHw1kjoeNDgonFYEQA/GV60PoaamK2UHi0FWhDo2Fl1zPJdZR9H0uHrQrBfEcjrlyAV8JLxv+RM
65jEb9zTwSrp56gAGKFgSwUA2pbAA/Ovp3oL+5xmlb2nNQ3XafNJkyZkaATW2O3Ppzj0IQ1IP8Oi
e3XDSEvQAYFlcypB3lBVxZtp6LVt3kdClB/oz0/uAzMKehYLSt5qRlNi9t9vtiUUOphy96mvpSMn
GwD8Ao5Or1i9e3c+zoIqCRsTk4AqOStw46aHsFuY+NnmfrQ0Anby/sjABIhH00RXsiRIIU+LuHqT
lHljLA10DLUYAflSgtTqT3Zl5Ifome+w9Nkfz+9bfu3wcDy54hj+X3z+VYHAgixo5I0ePag4seNT
J8X0nXKzcRsHw5v14buBSeWAy4LOZeCHnK8YqnzqpiR0IGjf9o98k1xpJqpoCFCzzmXwlahpDwgy
JntTzPqDx5BzulwqrxzMRInGPoYKjETmbsrRIrH8y5jjpKa8R55u7m3IF7Z95WjgKzoh/Nt7B5V5
w7JLIhDhkjtryZG3Mc4U/F9T8KUFLcAcrTs8M7EdVBID/MljuhenzargnNHWq26vaB5kLjrwNq2k
eTWazQ5TK/iTLuWkOErBFYrRKSmygbsehra+VrNSP0RW0hU1U8m54lt+eeK58lHtAvsP4sw6nj1q
dRTMlMwqfS04e+shFn1ub72UDXf3wGnklyo7A8jGB5tHejh0hPzTyJ1FX3D3gT9Y6BORPD9yL7fF
0TR2JG6fUDGjNto84/cgkmkh+88spGJfcBEcJbikDMmJ/JexwOeuOPSoi4/wIV70tQFlV2Dg0ifb
+6C2hvG4VkBkbR4Tv7SLl/6+/xJML7Pf9JF7E1WiiQ3vPwa5eeXoIVDLw9Pzke+QQLdS13c4eSr+
brogHawl3uux99aHtLbenruGPvQdYhIqNAMzHk/XTSKDvA28kFx61qUH4vtgUV3RHw1goiiOTDFc
l2xyi+x07WNxXULol2JG2v4hoeasEp2+x36ZfPV2rqGvV/4j6rk5sgDvz7FStoTV/r2jWJFFWi5o
ktxmMp5llcH36lAc3Dmuk+d6yyyHVNFqYyUh/YmetlFNgugd2sB0ql5G6hwJeKyoLEhFSCYb/O0I
RoUZUWnEqpvTxiy4LpdZA//Ra+il5d0ZgPNIYdQhZkUtvSH9oVdeUfxKUuLcYZx/ZGDJN+Ve2zpY
8fvotmVCARi8A6XD43iwJYosg+xKtgPKoUhTE9iHQ+ZwCa1koYuPdnn4hA0dudEDqr/2BnNBs9Pw
6TfbMP3re1gM6CYG1YbSl+p+5Y1fj3blOpkyu+u9/CDeT+rz5MUlbc7QSCQn9NTzMro1IJG/4BI1
/DZmCZ89GEDBYiGzb+qfULXyLzOWlc8s/hCCpt4mGUGqqxLOQA2uL4zV3vv69yt26sq8/idobO4U
unLIuDYjrNJXNmfOBcx3/d2JBDZreofCr55FidojNWSShflK7ucX18NRfwS2DXYR0q36kKBbjGsP
I8TX2GeDoIyrz0h/iDe015akbuz8ueXUgLJftrdrFREYVPHRbdb5drNJ+I1nFVx1uweJQo7Mgdkz
ae0ld3eNp189///yeMIsObRFzZ/qgTZZv+sD3uyTiS1/svmQai5WpQmmIzCy/oGFjMKL65k+J1yd
0l8bPKhp+81uOnFhBmTEY4Dn312Vk9ZzEn0p+KClP76ayELTskhAjN3YmXaAwdhkeArA8gDzgx+V
K1VkIzTrX/s0EP0H2IjatDMwOliiLMFKUErrbEX7Ul1qBpz72Z1y8RZUHugO4ZrM4Lr1TvzLGJYN
Ge7pZKACh58IQAqeSgxcJPEBj1ecUBuzeQYqq/3CP7b7/qPtxrWYCt+5+fjjavcaZlU9j6+1WqTk
lwjaPvP/At9B8tv2GQpQSQ17XE7xtqQqsoPUyw49fuTfk7mM7OJ2vaUyRRDMT5/mhYiVL+S008xo
WCGJSbU7YkzBJn0U7t8jpIHX9EBOleu+LA5GoIK2MgY/Qn8Z42GLP0epW7stWXtUBeQ7wuRCXkUR
rA+bWWmNeMq8vLK+b5nAnpBDgmxjFjZHptaD1NvojKryngOZe0vdnA9uX/gTcNVh9h4Y6xwX+UyY
f2a4TCsDL1lgoASojYySKY9Z5ef5jvM4+pNgmNYLoQ1/xbmG66ksk+Z3l+TDK8reEiyuCtJ8z2dk
E08w6dhykL05MYPtecMpTpUMl5dknXIpam/bU85AtMxZSINiZxc2cOCmb6O8f++O4OkfreJuO42C
vEm/FB3sbDHdn9SNV7nxbzZVdM91fhpgpiP95VWBQ9b98U3kCu8u/Z86VPnn57kCpIj/EWDqgrPp
9dvf2xw8sRsbnQS4aXwUYAWW37E7iE/n3oIm2gcXGZS5R/7q2xc/zp4/LSGEmTGLDjzAPacLMLxa
p+of6gmmwNILNR3Q0MWXoJzs8thcPLaTgwup/uoy5gZ+xtLZ5zt0rCGJFRpKlh2kUR5FurLWf7Wf
M0jDHVs4oyDZaMkdRMsckQSVINZYm5HwV43ZObmgUPDDPg+WrulMR5cDGLDxy2YcNq0WzlqVCntE
lq3GXABe+abUqphM8KuMvdrX4wQTJM+skagcgT7jaaYYx9Yjkg796B2DbyBK4wCMZAwWyxj+XrEe
KxhuMpHERxV7DogoVlO6v3Ahgjxtr5/apJ4AJ+uw5OmwtbAIiltP6s3ZekolNThJNNvHe5NJkqpR
kBzIfAOGnC6oNLyBALBjy+GLpamTTitIDcuJ5m9GTJarv5Qcbq55WxgBIf8gIQpZHn2maElLQ9OQ
pKZbjxHZNbi4uZJWA+yipv73rN3SGEueAH4hN3dk4/Qyrj+nqep+/d5jbXw91pB/+ey/ah3nm88u
Mzb2yK+mFkwIaKQistr+Ha0XUZ8+a7YULfeD0UT7qXSvAdI7YgUY2rTROGCUSdDQvmRpP/b6h9pa
imDdldcg8zXofAsxuJmrS7ZEjvpaSmDww7qXpS3D7t8DjEqQ1/hF6GA+CnyRWoz0yURl4e8wubH6
WnVJH609HJfRT4vPwo1dCfKIwt4iRfM3tSqGfa1iKBfKhyKkDBK1WtFcWXQfSfYc9A1X7g6ZNUt8
lv6ZOOWzbMhemNuF3EkwgP4mKMhK6OUJYPeQ0Os/mmTejufitTeGmHh9JfBLiN989T+5Px/JQWys
YUzU6wq/Zz9Ythi7qq5R/voRkQ6nng+1GBMRBM+Zt6XD7MqA5UhzqQpBhNkcYaFBGfl+37z4YqEk
PAsQXIo/sWijuX7l98aVnplqHH5K7rlbdgmhu6LabFUau7btn8NPrMDXzBItIaMBNADkTRK+2PUV
cBrCAQTNXRlUWMvXqVT1UERUa2ZkCQPsPoswEUvZIjyY1uUrOgEWVNnS/d8TaAvMYUOICLCFkMG/
v+tHY/ZtNjDUh4gOHAS+p3JQuma4XMLpZAsQloCoiRGqyEHZlQWAgbiGpzdXmoMOJz7GWWX8HAoY
I8G1xbClwRNznrP9pmFYIeOJB9xjmlv34NFCLc47OnqTD/yTXL+ffSGzeDrYkz0HmqzJufp+nMep
rAFHAg+aAiFCxjBHmYB39X4gcVDn0kpQ3/p+CP7oV9yvMNEIek+TMPw3cd5pBK3bYMomJ0GscktG
3KRyOyJ+p5WICyCBjsvl6+0iQCjfpU/mG1xkev51geYEq9cmy9NTVXY4U/QDtXdaGEjmR5ahKTkO
q2StzWnibsSR09BVCaHhN+SXfnN+5H89TogSn5rqR7a6AmXWcqWV57bnIKXfWExO0ImETCKlDC3l
UNB+Y1l+I6QtoEWKjbCscPxl9npx4Q71oEN92k/KcgVPUbtKpxYZCwMzm6zUkqDJ3sa6ue2+OLGi
NHW1jzCLiDVKCSo//61Ybiq7v9r6SdehE4ClP5MVxludnPXGghaQGneXOqLrxpNF6VZLweIVYLPK
tLxjXTEiXq+O3Rj1WAuvYpNrEidRAJ8Ml8RgzNBO3SRoAwQhO6S5vPYP6f1HYJjCAp9dqEGvMfyb
gI725LogyxlEmcWp0QbYqJGfAZbArCrio94VK7OZZfoNmQCb0fmLTzCLY9eUgn2HKX9qgwuxv6ag
v7SLjoSWfY/bA9aO9NbLk1gI8nh4LC7xkJEi0VKqvUlQ+to+QnHfxpDo+ODIe2jDyecsdq5UtIDI
Vrj7w7BxnFjTniXKjjwfKhtU0TH00b2Vzxt1cYNTsVXHhNgWJhzUYubZUDcL7yD+UDFs11JesoNA
4WXbifi7MlMc/ano6TR+U+Dt1dLhzasoXX9CVomGdDMLpmTF+y2qrn4O87L1DfCerP7rw9jbrKds
ZNSGc60AzXEaPAuBC/Uts6d25uYLBZEKavNjNK2BM2PfxzAYvSfTL/dBOgiqmJTX/Em+HJz6Htfl
QwI3PfVKB6+ruHZD4GRyEsQfrnPt2dZFz+Wey+62F20/qcKrQIO2CH2f3HizGLs1e4CI1vW/IOE6
TPnq85J3rV/8BZnf+J/IAyLAFtnfZDrbShoppuyV3bTzdjOFDY5YSM5seCItpSZzU7Bg+8Q8Q3U2
WJYz/jkwac0438LdKZDY+1ITYOrzo58Zl9q3Iacy8AkzV/Z5IBFGBuZpaWoYGe1dOuzLvyvMUpiI
LYpOTt27H9gCFvEH+o04EJOzdfQTH20GjlfnHFqlw4Mt9RDLxW8hO2olWAHUWPNYUK7HXKKB71Aj
sF2JJ/ZB8QzDjT0Ib8wjQFlj5xbd7p2bE9ulQ/XpOZTPtmnO6A9LsCrfnbB9DIaDpsrO67EkppDZ
cuHKpqrXcOVKVS9A/Fbp2s/qAxtDLODgpMiE3mBvZst+myX/FnboC2zobWdZp89r/TddD1FxNX5D
AlvCklsdx0EqX7uls1tguY1O1wBwrX2wS3kVRBX8M8jeoTJgSj1q9LD8c8uBQAKjtxSbpy+x9h+L
6w/Nv73Vf55cS+SfqECsoB/bvGb7cmFBtf24eBPGupVfWJHWBGlLTK23hI/WklumJuOhWUS8jJgg
p58qb4m8v4eq4yZXVOvSke8HfgUG1uNr/9lv7dPsKfPSzJ7nkA7aBoeFeiDnxjH0arD5huBHyuc6
fQA8rgGAOqiH6bXYwsETuoQ1vCPNMEwIIsrBrMlfXTJvNInlREidpLHv/FleB2jfW28wGEJSBL1y
HPnvjgSx8t6P/3w7BUnajSAPJTJogKLureDSdwiKl0qlb0GdGhe3bU4lPm/cNn9KbchSjZaJ+2Yb
CwMs7WPlvuX8feoz+yxr/15ozfD3MeuTZMRpMd79L8IIm4L6KApjQMTiDUkbCu8cjp6D1xtlO61Z
wR0l4MzZ3jlXZsFr14Uu6HfqyHlc4i0MDagtrmAFGjamgpaVe10gsLFMp5l2TrZZn7aSzqalnPef
CwuIjX5BM7a2L4gWjkJjnk2KI2lMxird2U8TJFsaiY/i8F3wU/lli93hBzW3T31AFDDBF4/DP/8i
rHX5Cdwbq/MZUXEUwTLhyoq86gnEnYfqXn7xFFdbuS1lWMmMand8m+wCd0pBC220GCToKHWQQWMU
8m69pK8vYnmQ1fZSQrCsBQmjAoBMpBEYCfITHm8hX8hLr4Lh1ePV6kh1/DVB96ZfbBNtL9A/NeWM
vSIY2c8OWtfdqvM24a5VdXGdjf+hikx15gZEFWfFEG6pTOv/PWyPwtUmdctZc2BS/Okygxso9GsQ
lBRtc+wrsZrxguS/4Gu3Uk3w7sywa+3wZCPbb/yc5iTJVmvhVSGjieEh+42w3nv/FLoBT66oLuJd
YW8HvH6bGQbRwNSMxrIOCzmiZ4XKEGJAKU8XtQneovB+cf/y4pLwfn/r6HwNZ5EocGdsi3R/KLS7
MY+sOLDyl65jpThXKr8aVevGdGvbpC8pf2a/I6GTN81eG+c8N4gGZEy2K0BlOUbRokynntdtplhK
6zo2F8TkILoqWuR5J0eBkjYagT71DeKiPXB35qaAVpAddehuNr3pcMhbD8SmJzePDZbjskX7gLhg
+0lexPjzXBPDjvyxibsA6B0NTMoamE86F2Pz6bbYwrgR5efbDn+0GPnk7/uBVIt0KbNPFfNMMGcs
VU/Hycs48cNBoAlpcNdBarqGzf3ys7QX8PlextZO7u9pPb8hDtQfY+fRFoJ0PeqC2AWe7p8ukBOW
1ZL3VzNnMzEPD4sa5JFU7RHFz+jvgemM9wUdFu3DXTP5L4eqRtzoTtK0z+NaNeCBwow0Jzb5GfL+
JjbqhsHvg97HM0ktnO5m51UEAMfxLouVoMdwCpcWS5P6r3QX5qJMt6yhfK4dlZ5NaFTyU9NmrAQT
SO4axHKAHgv1DJcEssgUzT5iRbZnEcslsaBuZ9Ln90U3xYkVqEbMFn//OxYvKQpOSzS6vKM0jSyx
XnV0ZAfgPyyZOwGoz3vdIvcM398s7Qaf2l3bn/6vvZ0yR0iK+Bms0yv0G8CZdbJRtd0tIzIsy6FS
kmTWIJJXxkYY5PsDMOf8cY3vVqkC6CPgceiwQ1GtquKR9xDsvn6NA2bS8LJd/y45BdjaI5Xw3E+K
vb05AzWEKovUeBphDxpmYcQHTA6rjuiDdxhbA27zmAD8kEEp3O2NDqTB+5BTnNIfA3atkIyfDuOU
ZvDjcpCnR9bU2UfF+irRO4BX1aLbju+aT88GJAP97LvZHK2hiIakOYK6FNAE8frawREnlZil9tgj
z6kjKSl4dwMiHem9Ox4CmWnV48qb6ORDjaLG9TMQGl7H/7ye4jQJvC72zYi7czC9685l9dC+ph32
wuhXUcvHneA4XnHT29W5C2aJ3JSUM8IS1GAT5Q4sDCIEPW52FLgiKc74KuvW2WD8tRu65aH7Sp+5
H70De0QMynZFNG93urCpSUlqG0H12lj3FRY1VYLuj29KQ6vUljF5zkIjBZ+purasPOFOPVExZIvO
aIsZohbl4YUkcBFOMWZRsily7xRDhbHfCdCTcGkjsAIFE6EFzE5+EayQy33CWfZQD9TptM+kZoca
g/Tiq3UVo966hpYUre6c2NYgveailvHhYSPPzGY/rCQHArOgL4DHA+0pEAxuTvOKLrS82Fa3hPlm
l/WWIJe3XX2GSKWyrkm6mFxSIARlzTOUNnZ86+tX8Q01Yc04G9dv55xizdJMuHa7Sqv7igyNRW8D
Ew6RPY0aLHB4x0cAbGm4t9QZxmVCw1rzSm1ft+8A2cJpMPW3Ns+ybSuQkCq2AUyKN7OifdDUaj70
bNdTRUZ0pBk4pfFJ+IPbLLAHzeMHIsjDHzx53uB0AqAMqvT0JVNTYBhh/6n8Qq0AI6ZsG5qTTwJL
V7AaSZbkwkL0dUE55h8x+55XvENE0rdN4KuptQ6HzzcCMyagHb3PreZZnAjNglupeEFWZdgZ+D1Y
sL/dcp4HfFXJ6pvD0bUS7+HYsAIRYimB1VMpENEv9ZyKAJtkdmaMuNUsTTnHe3tS8aDsT41deKU/
G/aNjxaZg3Q1lT4YiZ6jcAy4TtA4E/N6Kv+khCwvsGfmc9+L4rpUL1ixpjRAysVk0m+Zi5rYIXk8
iQjLTNESEHdiAQIjYC9lrz3gR1iq9ZrY3EXnjCvBTct5nkeuXXRnmbaTScwlSlWgvJvD2zMxtEDI
x7EeWUrE07i+Hu1ywE2agL0cRON/lwzPAVqJeLUZ98DUWlVXEk6TS0GpoMTOkgi4jzZ3QFm+EBIc
40lTMq/OAVjSbLJIUUDeRENU4GmPJ9HC7xCa2WZu2O7SgQWm3mZRjjjTyW3GtrRFBb0dI5SnYFg0
S+2ZWpRt8JSNiwr88zBtWGwph7zcExGMaORtBATZVPbFFZ1k/lBLVvGmulVk3Omlw+dAbrutI43i
z50e0WvocDOIbdwOyAi/AO/dQdXqfCruCexDgtxpCRFLS1mBrfHtCxzhFNBuVV5axM59pg8mj+Kt
ZbPiI0qUIZWkq0IrDlQ+eCAT7QgkaeL4rUerAotAA/YIB4OUagVBGbMbZiZ0B7wyJDY7UC+PmLYP
EEmB5fKefCbtPBPffLaBsbkdI/15Pzh7HsL18DcCvPyfJn4t50UFp5zWnbAseskASp7EE2AKGXMp
B2zL6ZEj2UvYtO+Cw4nO8UOpc8pI+fIzjgFGmbjyN26g/yKLrDNjQcXo5JGyGL/UGXDf7P2em3mc
Z4NLTbSRre2W123N9287KylIKfNUWsgOAcJJqcaiQpDz/0bZKyBDt9N9LqAWG+3d/hV3OOgIN27f
OQDlgpOxPgOE1zY73EG4Xr3NCjheAy6GmI5BPxR9pMKJTP3pXQPRcXW0INOFQ8sNaPBVgT+2DrNF
nPepzoOegj72ROV1L7DGRjVCncYvl3C0JydMD9j/Ut5yupG4h1xjUpvnPtICcgnT3XT94ftpJpQb
R1dywNEb+Y4fnYpcOvtfOM4JVDpBRDUx7LjqbbPUVYmMe7tOlxDFCOibS3m1TPFbyV98K2QISPZI
9Adxr6FwIq7Sot/B+DCFVXAgPsWArfmfp8WiGlBRaZYnnKCDv8sAaGxzya/71+adkdxibg46nev2
y+Y0dA6Z0q3UzHPcdDwhvIcB+gwDDEvGyFGBNFmd4B2YeePatLS3MNl1q+XHlN5s77odxORIJGfL
LXG6eO7IRGPGyfrzuVhFJIe/+o18orjk664CEjzUiG/5LrrdD4IL4FHs/XaTh6y7rvAL0NIYewfA
xGrLAS/r2m0U2WnQEpfkGPHrXI+/+VExyPte5jB98yVrCc+Y+WzL8VyUeY59q3X1HAaT57fm1OfT
7ygfD476ABCktdopDyyF9J66gnMANmMk/FnnrD20OHZ6kJ7upKx67dC0Ov5I95OSFxhgkCrXWyXu
O4CnsfXNy8rO5+7cvbgvVlqMc9bIUCl6hDx1R2/Qp/lljxDQpqo3CWtogWxwSNogAqsleTTYGHaJ
S1dVpxU+XZobOr5p7UNfbRWq5QR67LbckNfpjDxTcEfjEqFkeOnEWpfjQdAgO9lQn26gVjHNOM84
HjYxOGEQNyqlk4DxHgdZ+lTXnW3J5XY36ZYcPb2z2+r6ZimtDs1BUJzUvaVF26gLOHTmoNnTC3dL
uhZWUT0BeX7IDn9wfv1nkINCfKt9SfngUW4vt75spm8j6SV/b9R3Hpo0fKutQlD73S3nCaJY7doH
IQFEFQZDIMfgzQpGmfWhW3vq+JWUSjWCG5W9X5YZZY7H6PJSNT6c4uxlR9DmM2404FqIYFNthCoG
WQ6gJ5t5cqAFM+HMpZN0mlyx86NOf06H5ymsD5sxgjKF2CzSNOxqEVJcRUa3+/kVOR1HF1kcUxJN
9KLOXsOgXk5Oifta9BIXBLmKuYrDoGlyaLm08RSXy1hT4kT47mrcMMJB+oR1jDygmbIkMP2xu0+o
CH/GOc2/C8TIWCCJeN36bZuSr14clkhm9bJBccDh/1vGl0zO/eKZhkERUn572c5IpeQ3D566hMGA
qY22cCnEDIA6SQixxygKPxyeuuIhuwvuizw7bui7GP4H/DJcb693gCw8BRA5hN7/1QnIrUggKCud
/XY5w+QFAJH0FYblO3sSyVrZ/RvLPhphcWHg5VjYWOmeN0ajCOKaVUPmKmyp/LDcXhx1mqIS+Jj0
7JQfZyIOpXmyYCYUqT64wJ/X0CTNBGvKI6ZaD39/C0HqXadcXIliB0uCJkyKwg+PKzrWB9g8HqY9
zoT4q6PUuyiDSTc4GmoTYXLTS1Fqm011gW7HQKakJEZNjfQnEWcaI+R8XSJwmLaXhKaYxRcNEkKQ
GkAcQwK0SN5BymwxewJJzqNYrSwBJSuRCY5lnYc0Lr1JEOpNvYFxrDlXKZjybQDv0B9lrmEOjNUB
hlaJ4WA4YmGr6xgK6YyWoaQui0QH/zpa3//5ji09Trq+J/k/Za0yyRqPN4pAvMWxJa3vuThKYMGX
aj2X20766Obn8wOLTVF7HFSAfZSpf7E/6EndkGKDYk4PXET+6/qbnZofu8ZMpoc/2Mqy9aZkb5Bb
Kp3SPrT9a6LVe8XaMHuxlYlxbuufwYbg79oVXszH1BkTwIIy/PmXEn9dZSpCTBIrNFJ0ilvzAenL
S5O2mm91w6oF2yJcc1EEBxuG30Oz8r2wwySf9p6LGtn8KSyYJcY5nDdfNA7ZzMI9r+UEwdjcC1xI
6OS9oXBSUTzfKLeiEvEaW90EbYaFMc9oSQlBUyaDIoGFi1ef25w7ePbAFIBKnv/mRoRS1mvOAksr
nMTZ4FEmwa4ldC/Acv/OqG1E3OqqhbZ3f0dNKpF0HU8E9Kofv3x3jQBP2+FSNBA1azbcQMz1RBCN
/fS/Q9wY0/FMRMw6hFjRctOLfQVViewlJ2aF6l7kKVKPi7hUKoLs3tQOI9FKkjy6e5zTmSTfqEyj
x1FDBMkrT1Z+JowIn+cfO39EtrOTRiW5NQ87uqELHtbgQTAEzTKd/JuYWywGuvVKgDVWXltmhXkN
l4YmEY01aYO8lwHXAHz8tJxVAqTlEBauAs/UCggiGTGxFhMf4/bYElQaZw7BUvFG/Iwu0hqSuMrw
5FCIR9iSBopxm75vKwKy1knjOfTG6Gl5idldn0/y+pKyvbDZFJ8Yu57NteS6mQCVTfmdV0WVduvL
RXJzBa31yWY8L1W3J9CF4YlO3JKUa9gIYXhDeHG1WrxwNYT2D92KzDwdTdJ1MtLzIevbRAq3dF8c
0hzHZkq4A+ak//OXdIBZNQCnXDw3RElvUxns0WCMI2jnluPOZYWPqjD0qXMcUVHQJzlJYtQGeop9
JUrGCptQoFR9sYUWRvfSx60IklY6hTrTlcWv93jYuNeCuZtzF3Wh7fyOFjvUoER6kPmhnDmyN/4u
9CemJEuk4pofJy8DG+oE7kU0N9Xx3H55hvvEIdh1dCP41fDd57+dEYrSk1wfg7puOtPtMzPeMIx0
4ZSN54fMxzKtoVX/iTu0sq0UyB5NSpmglMlLZKFie/LFyINjglJmJ+MEDgve/Ml/wdnOW4YMYytR
RyZOdRvjIxEgkfFjqfwpUmAWLu4fZLmc+9O9XkPZVcMskvvUun6IA0aE0hYXbcWFrxhUHGbbXsja
8VGwuqCQkuRP7vXCsamw1i4A2mS3fo1zdUhLW/MlISDdnTTSIxgadhsgwpIMsj91eymGYsRDYCnL
UiutqDfp6tBXWvQOgVXIGFT3mHnwLtBUJ7nZiZowGdyZw/IOZNnoW2IutC60Jf/fjPkpFHol312l
OthUQ/PuSEYz6NKNcAOFHH6iFq56XFHed7rdCHITEWTdxHROuhNgbgOUlQyaGQXYxeUjsuES+O+a
0sG4/YX28VwvauhoG0TKvjIsuLOskwj3NCpuTGpvq2EmUhtupnFpyzC4DW2zJzHDba+I5b3+3Aqc
nAG7sKKxoMpIlnNNtOrqExnpGSGLdqKCNPaz/G0aXPLCPHpEjLcQ00BeCz7VINEZrfo/pQR/Lh5/
jTc/1z7OIf5ThyoKXVTP0TtiYSPBtX/J0czcQAiPKdNdDvwyKplUI8IclwU4lJ08/qFBFKqK81hg
6TbrcOsKg+6qyUtlb7n5wikR97Mcjmvghjks7v62sclGQ7RQF6A3wbNNt34G3gegxCYSLxHp9jUb
lb3p9QHcvtBdHi+vh7CxXTjS+CxPvXb8dRuBy8NpsqSQ+aUqNoQDvi8dEF4P3UcHW3Ivnc7UTz91
hG+URkvD38+J4A2goyyUMkflGPaihny18tI9y3WDUeoz40y/338MCZktz3FNEVpqHrzbBb3txTLO
i9WueCT+oBcCwZrxiuFwUz6malcrcwN7DuHsdTS6pIqoMia85j7uE4K4HytnNUB0wemJAMh+sbV1
IjDCLpBt9nY6LHQxTTLUH+4SwlZkBBAUPZdWA8ImQT3KqT+LOE7E8Z6SayRyuH5Qamiio8jvp2dM
aY+8pMzIQntWB2zH14IKjMDgz9tsguJzxJXH5X9CRPzg608R6fR8xNZY0Pi2bTZxDVBioOWSHNHD
dbBMii25m13hPzcXCJtnUJHAEe57g+y92A44QJ5XEhe9TqOlj1mU9vfK0j48w1Y28g90tDX2s6YB
Od39bM8HuLHI7Lr65VhradeBC3IU2HnFkqkzXkQUk+V1pIW4RyskqvHvwx/o6Kg7UPNZs2umZZPv
bgZwmXQytPd5MYTNkBZbuz3zKBdM0R6llYIMmM+GaJ5AOkG61UZZzsjC9oMZ6cQliERnPa4G9tiP
bc97qbQA6gd6MYOFRKyuP1IRuWfcMyLfH0EfRiDo/Xy0C2Q9MBEkj07gPrvpobUy+Ik66gXlpqyo
yJwQzEiimQ7ge2mc4EQ/TYko9Y5dKlLuimg53ZwkW5SFAKF0jYABs4u2CwFqWSJXLi1rBr1IqJR1
fH/jP3X+GoJ++diQWFF/J77o9aZBh9tUf4OoGgvbmTSAqWJmMh42020wXEEmYtjUcs+YeeKY6E3f
CSdb8ttfkgeybqOd8QH1GNsqGk3iL1ptcbSiZTFvXF9l4KI7CcfAxIhpaOD/rSD9fXv6br6+vhz/
WYo9P2ab3MeFDpYvLFP0/5UV//DH+d413WLKGX8hVw9yKpI1N2P2pbPC5Au4rlB4o98bsAU1Wzow
ZZnN1qtNk93JvOkbRx8dmsRkB2vXdPJAgutHM70wym//hXPJ/8TVIdM2RyhmCvTLzbECTuF1e2ol
s4McZOkzMuIAapKRzmtcvhLaLbvlb58uPJSJ8/KgaWLlyL5yeUwx9NwFF1m6/z0AFcguyrWxpRF5
2225jPFK9j6iaP7G6HQkIKvKDy7DpNxNUnZ/JM8Yj+hYGRwu8BQvLRJvHi7ZXH2gHhX61blYZHAF
Dpy+DhpGdTjuXeWpiJctG0LJQUHMb6E0L1EZmS1D88hMIffHv/6EHMHX/aPHvylGdrTll0UHHYnc
2FhKTtx/EIYUjy4sZjBIdzQJ8X+DM2cYCkzDn0LUm7sPhO5QS6OTUYSW0WBNZvIlrF3NCbLO5fFQ
FveroRhtVAogN6I578B0O/N7SlbS4QCsCldAD0Y0vmHx0tejRFWzDcWMlfuTZ6NUELG7PWnSA4zu
OO9ty2n4jbl5a6WKWkBLeacX6nP6AmCgFErYfDzLEtAiCQslNKvVbHv6600zgGvUZHzVCsjZDpNL
BbsbKFYZs4hX7DTLMvoF6/jP+yxSpXgv5s6tmwFYHQo50APvCC4783zVUOIqxB0U06qM0MMGCoPx
1EDwhQ3TFuwCS5HMtP2nxRVCPqW95PsiClr62LJuYt7AYkFhOyT8sRNFEgKBWP9xnXjUOTaVHdlF
U9BqOhSMjFKTEwbXnW1oY6EdsHJmYyY8x6oN8uG2yugayfdATPJ6GiYsRdOts2tvj7A3cCcbdSxc
N9Bh99guzv2a2NE2UQpMAkWR4060lzkjp2wKh9DexVtVUY0H+I2iFiwPBQborAB/nuq780otq0ie
nHhDdZzqizIWGiRBegLK67Mu9kn6JfB0W+0GeyH5cnuXk5moZ/HnWPfrp0e170RsCv6d1HqiVDdJ
fW/6tjl6RFXHwPg8Jn7TZWyMTksVW0ePpDzkyq5YfF2NJ/mFREdSdcp+xu7Q9uH282FOy0QB5hp9
6W1kAGrggyFoLAKWi5uiw39r1JIPILvdxavfHOQY46H+s6V0fXriS6AIWzv7vJJWErRe1iSEodrS
jkkfo0+Ah/GvnyOT9f85HnxDxf6uJq8JclZEr1RK3NhT7Dv3aVqH7ruzhTn6jPPt4qdCLrYpVJbG
CAN/Xo7DFKn0egL7x43LYnJwDK+vssmtGkSmydCVO7OtdD+MRYtrWh59YTC2G130TvF7zkdlyJwa
cAuIi2zHLQIvZfHlUrHAQp9R30dv9sRjgNtwTh1WnNlAhLwo0+/G5QUWxAQGoqEzk8IjQpDPvejm
pmbR9fKaNoxlnEC82RtClBikGyhpZfxOq+VOKyQo4B3v7hH+GB5F7NTXbx3+SLwO4FYDyyV/79cG
u/06ZoPN8CUOmyCOijDwNS/HNYuc19KhjOQgY2KpbycLAvG1Jw61rEAA2/O13VOXH1HtuumXzP6W
KJaikVjs9xtqXrh0GFZyzc+ffG1Bn2R6IKmBbGlAkruFm/m6/uIUF1b0EKSJvoMrPXihWgTmtb/c
HVM29kTBdfOcAXccozuypVwYQ2AF2TgFM3VBIBFoOFNYeWB2eWfIULTC++QHvGZHpeupBlkmZzLX
lh9gVwBGRghX2lP1sxT70oNw3hefYD8/sB5Ubzp6+kur0dA/VpO6cLEShMtM/45jjD8rutdDUu50
vEaw/TDT3jfNEHLTzyHntqkK5XnBlWXXnteqgHBAic9r7qPywI2esEgVCZ7fnICyGf1c1PFQofuw
DgqCYOvHRr2KcoLPEDr4+xwquZq5FtmCpPM1Od+kjlMGbnbCn+NRqhzGcUZBEpJOcQCtJxPFgL6Z
qwF7+KqCyXWTZKZZnYtNtS5LKcAlmt7P2XmEBmsVDtmqF740OazICTWedMxuQL40Zrn8dDWkYLu7
Q7U7Jc5lhLwc0RbjjAPRj80XWPrjp5yQ7RRiM9W3Rd/WJi95gGrAD1OC5ez9JVe95LzLLOjSnYTe
aYCci2SjatRjXwk/SfDotbufPDs8v5K9AXT0rG165GLzrIO8awciJC/+kWV/ZtqSI/DPNbhkXWTx
d5TRwJWBMBQzrbUNaZiWPw7z7pIaYh03Z3Nez04fsLJ4n49IefNATRMl0DxwEPASZyJNTWV7F0yK
xsMYYo7W023Th0f1gjBYYyBHxY3twWFUbrT5JQPdRxDZSuTXrp9wF+SGHGPEpQG94HrUZifPoaSL
CNrWba6sK80NcuH/oJNbVX5PSfBpW1PAmUg7zHp/+hLUAAfczJOSZJvyNgLsWaHsmFz3TKYWdxap
yytNspm/+Ku+iss8V/3I+BKR3k9vcBM5GhQDWg2funKC8rosVTp3dhv9xsyGU6014klasxmo7fyp
cfxbB+/bMxqx75wg2y4221jKuHF6sw+DYk11BOb9auPJ2qpNNDMhXdRU0wt/Idka4WyrK9LUQG+t
GeMAYyI7t83bzlctLrTffQmUS+1AxVAc8yDDomXPiPvXaBzaW/7f2TS05lHbuUOAMbEwZauh+KGY
LozK3zd7lHdeGaLrdkxsHMIg9aPxQ7C4uUCEHPXybwcyzQ7RgvhJVhTKEg46WQlcsJftPu24kK1k
2c9pAdilfRn0d9ibb41pBxZBAKvoBczfx3CoPVlgiluxLjHpk4IOo3Zp98sQBXVJ5u7R4o2/HFH2
au/rV/8jWVZ8Vae0/ynT1Q8mTJt8KaA12mDQClMe4CbY1GKbjp3Ls9OZhjYHpLs6DFhiOkWazKx8
ekxeAEpmRrqb5GP+DZCe7Lb8H+KrwlHnj1gr+xcYPfNS19Js9CoIc6xQ8fEULyzVDPDeIQFtjQTA
Nau5+P0nl8hZN+16WV/tYerBkrc7B0j4kiYfWDKGqJhC/Gv7/36KdFeMOCoX98eHtEHyKJnb9Xph
3pHF1c4kOXXMuDO6Oi1Q8AXUExUq/NBtZ4YmkB9IVxzlrAardg/9baLEjWocKziHxLU5V9m86D1C
mBxSThbR+7E5gOriIaAtOnwGqdHHMsJleIJ2EmN/aEbIada/Y/8CRpHVtfl5Y6jWLbj+N+Nss8Ud
xcChvT7MfnOw6cOpDnrTQVdGSYsUIGKjRc1vrtd23QANieEj+YSE4UtzDLRnd4kiaR1JDrtv4HA7
WdMkVL58D3KVgySSNITW9VrQw9NE8/YcuT9DLr80I62ttEOiBEssKwbJC5/May21vqbBVIbN30ky
cYyd1Qy2YcZ6miwW3zitHLL6KjVyrEtk/FixLvO6h+eDyXpcRv6VtHpjjAmRTGPDIZYo580dk88Z
ISoO+kRS0td/TBO0/fZkIlJcF1HGbocRYuyE6TfvP3+08bJX8ff++d5U6go05awbjVptccuZpyCs
CUwv2APbMGoPj/8+KL/6hVIBWOvqW6dvFKNGDKIzgXekRwz2AmM5AEviz4ZImkmmo084c6q6oysw
hrVBs2SiWeSMVK+f+jnOL2YPa5ENCPAuUOQTIMVFjt3LFemzzNw4cfrz5CRmeFHTYCmAObUHyuSw
dTDt+Rg1jsOxU9VtnpqoaXyIeAfV85oV3xRTOQTfuJjan77GFdCrMNdruLJbuwFhrHMeqOj+kGkM
RD3lNzFklDlijgZXFIhYlXm4AeUDe/9HQwuP+TCHqukAKCz0i/t8SeoReUxHFSPb4C+8UuO6nPhx
tlIWFEDSaUn1k2x1hzPMjcjRJKRt5PoTNkK6mYuc4/2ZMUzFuoZkn4kgvr1SMv3snjZM53EwHImG
kwQFRPPno+tMStu4Zg2DsEORtLeVdmJievJy/6RqmiuMzoXqz2ANEqPZBp/EUf1gFLMWs2X1XzHb
Fmrt82juh8ETIW2Ei6T07jOjPw2Ftkc4zvJ+hQUhJ3j/LCxwp4/gcJmVemnfM4rF1NBSojZ48Kuf
apEdajpjouBTqimL/KD1hiFlPeA5YASjfNp61y+ngOg1L5KVTOuasS5gSBDSs7lYvthNeXpwYw7G
ZTBz/yenlZJqq0P1JukmVN15rk1yJzuYfCID7lyxjIptIXSCN9TckvpP4Eart4UQPcncMDnAezCN
FBF/BNgeoc/PMI9OEFR/9tercOh7YpXQ5zKc6/zFrJo3rad50nLE09h5NOoCeSTbJywVYzBD/YVk
AbyGcl6LmTpdjKknYlSctSdSjUA/fDR+6zJ1Vvcm5V+6CAdtFE8gyOmF0lTf33kEH2fu1jdphQc1
oNavJyBAlr2D7+/97cs3wKpoaFrqhpYM0Ge6Op2Ldn1h/OwJcTCBwdjZ1LJE7SC42eErrdjWof5p
Ht05YmpuojP/3CnTJvzIqd6zFc+HgT53Eux3nAVCmsLsMx8v5OXFXxsjgV3OMibjcoEDLcdkz+HB
I5OiZwz2GCFdqSF/QVvLayAKmeXwGsX4nLFbqDLHL9tte7WUWNNdNGXrMeejc1PvXAuWA/5PlW9R
harCAZQ5FWZvxRSWxJdziOxyUiBaubm+cFydRDZCLQCWH6RuMSTaZr8fiNFnaHWjTk9rgALz97EM
ZfsmH4DQgYI+W8gtd9T03CiBYPWhoVyJXxrMDRUi2Js0AX9voVrEOf1RPBhRobWBNr39o9tNxLq/
6GAJlXw6944R/yJ9D3RxLU4mE8wm5AKFeEH/tVENPq+wclHJcopThJ+rbeAGdI2uSqfFY4atEs34
hKoR3LBlPSBx1e4HZUTvsahCwsNHKYp1Q7/Qwa5qfoJdJDCkL3+Jlfr5rj4BJOsrGhuExjkFQ3c5
tRFFFsYoSDAf27jVhAf5k9hyOuj2eyEyuxxKwNwr0VWkvxc56k02D6kOyqLrXZQ7mBNw9GVYuPo6
YHN2rfllfclpvpASK9UwWGBYcDZTqkae0a11J5EuBLtnObTrJXkzVSsF1c+4ww+izYarK9jypZfC
JvJzxUK56yd+9M/AalmOLjUfep0Zx1fQzzrJ+n8MVo1YZ5+ILpsE/SM06HVKW/T+F0fJgbLLrzBy
R9zpleYPTJ48mAIWDgHTwYN+Z8XgJtu5XOBd8OTfcTZPEOb2hxMwG7aNdO6d6xgXAYHbPs6b40jl
GZvAqJ4haLKv3uhubcWqdz8erENNUKE4waBYv1A1Ae2A2BoL8BuDs6ZgzUf8lvZ3Vc1eC65ef8JP
tPfD9e7Wketp/E9f+iS00awqZNCwPA+03RkL9r5vMNC4jUIQQwPxxhOl+k/92TjoWEGJkLTV2Cqy
D+E+8DetSlf6VN117GHueJq5BmyjEA3qTNBWBj33XuOL1Buu6GC6iuK8ogYTmK10BDb9h5Ky11nk
hG/2HFmDePh6PbnCprz9lqUM5Sqd6l3+pQkH5fXfO57e79R7uf2fucs9NDZREgIlKnoDYTHgfpEX
WBSwUy/RzBWjvX0fWN0WXJ4w1nq886xILEwSD9oILpHnqhIy5oIs/m0OsZQNo3ARxUxegPo6gMcm
DZoczI4IuwM8EDi5SU8226h3C6HZOW0t2Uu9aZeQC7da1MpgZ1xfBs6GdAGSFZVIYakshvKS5XL7
WfFD0IJmtXtGKP6eTKQ2xtFp0Fbcdr8nEGs5YgP1n4iobgCGMZunPDP8SIhFCQXU3W6fE8k1oEu2
0hQrGqkKfJQ6YP7mn6oXRfSUi94MyRRe1XFFwr/+q1apFsEPEQfutAWzHh8o4Sq6TXgJlhRUQimy
fO5wJEfAgcjGZ2foI0jk4FtRd6I4eg11HMeUGANHABIng627oUlUqkC+lQp+alDehOcKxab/JSU2
bm6y6/91xV3Qb5+7FeMfEWMSEoANk2wingPeVQyX7HqHpM1zZTM7eRlued/gh8Y6wG/V3suYWpqx
q7gdwO2s+MwddZPPfd8dhNt+4h8R5/pT1VO+9hWgoX/j+N3QbJZiJ0qA1Sk9fBcn1K29f/98B3lX
1UkSPYgqUEEWvnmulKlkDZ4hDZwiKxG965oxFsbBYSqarP8sQbBmphYe45JnbGfEbcvtENTJMtwj
E9z3ZGAhFYHqPYOR03P7Q/T6mwlVMZYaIWfyY9Ji2DWTJ4ci6n5EVoPJOlBrR19CgaXRADT2zOqi
0SvI4j0TbAPBxhBsJsfl4vEE0mnXgfC2lKFDK87g+hkUMd28ONT3N8/BkVeDgkO8N7w7H9NQc4o/
4x8xTpd2Vyk0mSU+KOaRXAFXdXHhNTuR1irMHkXnNaqaathwCBGW4Kqm0lSofGYRp78Iuweor/Q0
kVFpSVG1pIGPQfOHLkFeagygBAPCTUdYgZGFsRrzqDYxhmeGmxwkLX8/7YzMyIl/p7CwPh/06fRJ
9TkMX0zoma+CrLrCTMkwr4xJAfOIsHHW4ISNE33YVMINUbFwRyr8ElsIiTvDFYLpgDDUYTsOa02P
iobu8yyNavebPPHCN6CtFUDBj9Kc7IIN3Ig4cW+1QXTYIHHs01hNqKrBeuiceUM9p4XNoxGM0Xmo
fMw0tqX7sU5Mz7vF6NEjE1Pf0sq86GpNp8apwJogQvH0YAtgrvgDadS2/ZVVGbIzmrZ4mk0ZmVsJ
soMHyVcGVSVt47q6eLVZYlHx7dc04x97+/51M5a/xKbUbULbJR8Y6LNcs7KABaAj6Zd7eAdfztu1
naEHPBVwbPaT1VNb4fNrDBbCBxk0O7CBszHVjlf5LAzCJJMB2LJHnKf2MbwRye7JdwloiJsI4NTL
LEMZUPQq1FuW5dfkqTeqAn3Hyl/YZ8iQ3GXGq/FCQAJusiDzCEd5vkAlZmXudUhl1FJGIoof6spW
BECXlNu95A/vv29mOo7sWy87RMSMH9zuGAiJcz7b55n2tATj+cIMRDCHeaTkD35dzvftSnzQL1Up
zamjBPrp/Iv1rBFXSHisUcdubXNR0I/aA73Q2ZCfTwd83ptrDDvzEqLZO0BUGU1t8pRBl7Jyceve
W6GG7Y7UFRfKAjZ3IUT7qTISPC77KKRJu9el1sJubtYj5LMtjfIL2YPObYDrTy8Knb+nOZAX4pOq
laJGVgKyHm+UlUzeOyAmmOB8szu3ROJAWQ7nd0XiTmSBwA3PwGfb0Lt+NpPr2R0WO3G9zIqA/60t
2zufFFCqtNi65467YwIgfSXkTDjCot4ycKzTQ3s6T8NjeRZIDZY7jkDbKrU4ixQI2MpMsAWRrnL3
ZJ5S5uoRJfB0NJksQYsRICOkGi3kK4AZfwIOr0U5qCC/CaPsULYEUNFGrqGaLYUMHiPFIsQPQ3AJ
n8GkbgmnPxogoDQoqstEOST+G4xB5BjxkMrIDAREurlJYdohXYo6hOf045grVG2FVGIAwkRwhbnR
sJQ1EQ6GLcrg47IBtzmCQQcryhZLlbcaGqAoZWkZqTB8u6om5QUTqtvhLJZiZw9vxIzF5rNyUrbQ
uijRVvNN4UNouwUyyRBqQ57tzs1O4q1ABZTnymq9WYFSAEWz3YjDDp1esX0qqdO+nVMizZ3IlFMK
MWY+gtouST+SmZzVjBiDSjsC2l3cdoKJx/xQp2wtjod40pvg9wBiLmoBqSr0s+e3tpXQZWtjHHql
/bv9vmVMZb5rmUBOTocRDNQc9vVXRgaWO+pFIQKj+J9WbwEWWje5PD34CyalgsmwWXCGKsEzVrcz
l/WRgKI1dATd/kqnJhF3LzPuBSePnH+Gy0/o19I8Ikn8zPKax83MG5EorJlsaqhN9GxJR8MkDeO6
cSRFB34/DBkH8tdQDARyaff3WtlyNQuVfEZ3TqzIC/XfgDO70iCyoBkFPnRC5l4hAUvySiY4/HP4
AU408ta6G2icoCfRun5IWntiHn2260Xkx2IeIkiizHT2TZZ7XjNo7g52mYSo5MVdH+/R42StofGY
V6Nd1KvIP9dzbuzGp6oVKjCQzYEIZYdbijA2jU/OLaSuzrowAg81J1rMtBNjK/wyZHHDLusZnMF6
pdhH0IfJOiV0G/JEm6NFIAbX4vCKwDyKZyZHc1lc1gmC2vDGaV1rrZgxRoCb0GW6++bNkDJm/fR2
sf+zyvTHBf/whdgPFnWEzwaN/ORCWTPhW16091PjyxPNiIhivyLl4SnlHlehDG0EL+ClgMvuNKk6
4hYdo+DsiCPYeVsfgZi7LTWcALQMNo95p9VaJOZiDG/GkwnkpzP2xYRkHZ8oi+4BqViI+m1ga7iS
BUIP8z+l0qp6JQQPKfJZHB3t9/SXS5XX4nDPOoXf09AKKBuqpuZK+XYIIcb1PB+dE3L44OZ6Cv+j
EztN5Z54mnTNa0TfZoGBuralN3ufgPOpaUgB+JUKoU9PK9JlFmlDoyYxLk3a0wqWBuU6YW8fuL9v
hTQhIQAnQsVukZiqjPaY77rFoHLQdLg5yB2Ct1L8XTBGBMdAaIZXm87HIbH/OVZK6pio/zHKg1LI
CDPzj8g9wG8NknJc2FdqA6NfQgDprfuDSzoyC8L7loKgaZ0ulorAVEhSu2/hm1gXPHekQCiPiFW8
jAhUqej1WbZ9mMcVXPpEH7MX9vTEnzZZZ0Ic8mObnvY2I0Zzlb4C4J5BUSi8rq/iHq5xQpOC9NWu
HADEN9oXL+1shCEUJdQ6CmqAh7HhM0tRJZlV278JUlSmR6/xbbD/kQJI5ESe3Ii4ibtO0jkpvZRz
lIna3NVHPdz/QUbRYnUKv25JKqLPBi+DxV+JlOwFYzNZqJgyjw2Q5/K0vqdDgnqdPpmWLo4MtTpJ
nfIxmV5OBKm145Dnv2JEp6fj4ll4J8uKdBhl+JmOmqQsIvdUy5zsH9MPNX/B8lw6KcCtVd9dvdod
tEYGITDhGSB8WfxYtoyeIxXhEY918gBZVsgN+MDWCDuz7pFOcjEz7fewUuOB8Tn/7qscDQ95FS/a
Drgeg9xVbMXa5/GVHF8++/mPezl9fokkFdtWABK7nloC2LPQI6Y65+4P035BawZvOHsI8KZPsZup
XrKi44YjznQdm8kg/8AeuXq2yANJz7BglYkrAUEGwZoe9MO3KsQ8UbpUQiZUobxP1we+4cDfPB+1
NI9sNM3TdtJRq+8NRA0DsncwmoXu6NzS/XWHVNFXv0Lqd74Do9rWAr0ZTGmGHrvbqLbMMPagrOOT
zrt7E03YgXlDbI/+eW551ZPjZ+/zGQ3gIgENWSiMmtunIgc49ajUlYc0jAnY9PXCcmAkNWfuf3aN
NvHpxeUJSQQSHDWXImUmhM5fOlap76K6Y4KW/tmWTV4D40oL9+nrlZZqfawH6Zj5oZhGSbc0iTjO
I3yRsN5SCoAtoAjiVBgAf23KHtPooxrWpDzZeFIcqIxPKFKASncQIC1kbcXSlABegEGYOBKTppor
JrUJwS6kQGJO8hHvw0p28MJ8ldRxqeAO/IEO96CcylaihgAWtH/Wysc++96muIWzWkLoRt6KuGiW
1dkOoss4xpE6rm8BYGGHE/HD7SXUZUuDTRfnrMMULKLPz+1cD2iECE7aeZ65lGBD2TyPThDJ9dAc
yCxoP5DJmhMHQQSd6QgyoUIZa5o8IdWX/cKNFAQZrAlGgk1yJBTXIFTWeLyA+PcGPdCUEP9H9rD9
YNqDEtGv2XBLjimeCA/I1yI31I8B1K0BOsbPYEAIoltmh0Mm6lmIg9m7tnYncLx0R5+NxS3L25kk
kVBOB8oSpuX0L1eVD2mbIc6C8h+mCPkvF0nInS0Ih2ILEIwgmrVoeWbgMeVt/y8QPYDBYGIxWf7x
vqZYZ88u2YD3kNCFFW1badnLxzQLqlC74Zol2kEbjmuoBYpcFw0wySBPRF/roLc//ct1xLyeHpJR
2r5L8wEASh5cRJ5Iz+2l3yqZ57uqVLgmQWjjFZc861Zy6FjpU+tOWHmkEeE7ACSyah5DWCKIVkm7
82yIKLRQEDMFU5nfjHQ5EvYBmxZn2XVyEw2/qOhSB//kc2M//HN4ZuOv5M+w4YltQXtWQjjfpx3t
M1wcj+2ZTkHUGH19HKlwuD6rKEWkAImEya72auI9QzmFCcmIvK9Y6iEBqyT3HLF05V1ykbM3KE/m
4tG6jcuIQUL3DxSkDCsOI9xK65k9cdhbuOoUJosx1/wjmuOf+21LkfjLLSKwcV+Q4SHsxRNRo4jf
NCshe91jgVTHpOjSPH7aF4szPaxKuigXXd1Y8VBZi8wXX9LJkodwfu56bG7IplC7FDkBxTWwWjcH
RtCBcTTgwqO8y+dgSgElYj7TqiC40mdMv0TXJV5Sd/6tcxkH+dljSv3uvoaPQ7UngzwZvQ9IbaGc
+vGPbTvdEJ6yGgzC9wrKPHC0FSSlJrsp+ZcGZ8v6Ej+xaFWRnHSi0CLHdVaBWu+u7f+q3d0rkW1K
ATslNnTM8hwS3rpw/uzRKX0RyRNlJoo2O9zvKSp4tfmgoDOhZwoYfyLPiVGJrnAd2ojLXv2ZEvi7
EPFcM3KfUnDsxJQNYD73dbM0pbs+RI3XKSSjPBt81HubaVkyP3uJYhwoelRhCF+pJ0SgIVXRQNT+
6sQdjVYWrZdnp/Tg89enKknkFoMfJFaSNhTBDS5enI69SfWjZlG3+vNCKf/UPxBhhCsDFnXl6OZ+
v4Fiai/Aq/m9cvFGLiictSYsZ5XB6unAVaZ38y9lHtlpIEIuHH++QY18wpfC7lJWfgt2LgR//ft8
y64A4YzgJ2X1n+38WMduC7oGrQTncLXKtu98fAV/TxcpcP9Q2G8B8Xnryw3Q/MbJZ3JdDue5FLzo
zGfrxY5HaIgVB9tAtx7Q+MyDGC51FstlfGwb/uTOC1kqCq/fIPnXgXZ5vwEMzbmlp3YH7vBp77kT
HHro9PAsY770gPuVIITqXLeMC0BOy9AaLqMM1hSAMyGJ+yY/fR4b0WuxC+902nYbqohMXV7l3dDP
FcVddf31pWlxB4cwLp0FRrcj4vivtQINo3NUhsPH6YTceUL2Y7AS9pGo+pWV0FI2wiomVYakcVWY
+6tqkJkkcLYJa9q0uxzHCndcSLDuv4OJS0rDUk1DplD9K2GhhY8rWa8C55d5JXJcvLYSQfiKQ31+
Rt8Zk18sMrHOOOsmR+nTxsVLICxTSPDWh4PypEMUXXzh3sMOqGVLZvYGHbBxCeorBvF1HKAW2anF
1yIa7pQ6TB+chXmZaQO5y62m484qU2mrISsrw2xn5ZR1l8cKx2s5okTfo6w0qWVf31Syzy2V+PNv
/SnUgd1HNPCk9A0r/IVIL2rqhsD1l6ddTtnAAIAbtNwFk+4dnWTdz3jctxtHI9z5daqCkt6e79PZ
8ulcbjJ0MFI4xZ31Q9yuNAGY5tPc8f4JrKhzJXvIzLlw3/GowQwJd0xBWvb4LNSqf6MeVQDOu7iu
PE8dlltyeUpaF+ilTENKJweuBNyh2Rt9TbRYC2K9OwRihHwIzeZ+/egC0Q26RA4zL1l2gZrd/Hkw
Ezj4Tah8Wry1jSDafUGEovrlSQXvpPivzXPMM0x4voZNYnYhCAW4qvgqRWcmj3ARmA4uU9HzUKGE
aTEvv7CX8MAdzqrbdG00PBD3Pu85YQzxSFN0hGDGys/HFbhHGEU/HDmWBVFJtljdbHNJ026Epnlc
+xcsKw27T3+kpdfoZ67U7Veh9YL3lxdNGTGI7fW6h6lg3hqbcJevmUsJXdqarVZTLk9CFHIAdHcn
dwYUUFnHRwmbF4vdsOn+CObQGNuKhDf86q9AmwD/bJG0YgWT30mxo6bnzqYdlhwaAejZ001SznAw
pw/T5tUMzSDCJZ+0y72HDiFm1DysI1zsQ+oPwcrLtDuoAMqXEyBtoTa4aGg806d5eWzXV+TMt102
q10dX6gbyTGhrxQxOiLo445Id5LquJyYdH9zodJe9jnCmGhFwwYu4Kl2MKyPT4qgCM0Gjf/28FW7
/9sXPBtNFY2FJWLMQ/OCv19fV3FVNIVRHrajnQFPXB4T3BmKnUP0mSf5U736qkHOuwLJ72iyUfzm
TqsMaCGrMHa7g/rOwZin9LVb113HdpwwhBLQLVEuSIXIEDNyMu/wQ1S4wLzVw9aNM0uZnEGG8jEu
ozf7vzsCxqzPbOKbHQHYrX5I0dVFs8E2ONhfcUY9xElh0vC9aHJVL+Xp5rhTsbIbQ6uveEIviJPq
qMzFxZlUiw08r8X2KYmFhlZqBidh3GCLPxPJvt4eWzZSlA5fE8FXCJn5EIOcZrWqiwTyCGVM6P2U
q6xKFh8omlUCDNaIheN4a0gTkWoEp/cri9UR2GZKtd/Ph0ODSGycF+NsHgeD56cFwEwiU9DKu82H
FoIwblRcz+/uC6/hReZ/7ADJ8cE+rxNA9kVMSrTIavYeSfhenqRyRsuYNCnLErzwxwmLJKYzbrVY
N+SiqqW2Vyn8J4gDbct3aYR3egAySdlS24aU5SAJ9H0w2htdvBgNSxYca9rX6KLAUyxmp/3GnwhF
uPhdqGBj1GfpKn7lQq0Ol+J5KzBLUwl+R/vbDn+2fTA3cF0bM7xN8A9rUW51ZXYY6ZewcnbcxxHh
lTcvZp1WzEvqGO9/6uSCHFkfhc9ZIUUgSstG00B0zUIbFrWRQlvltSrvmC2XEfBD25ypiFytjKK7
N66NmfNMGd9sFhbcsGrnz45xzDSND2GMYJZYSfaG4QQGopAZakBnVsBH16c6BwT4l2McI5lxuegb
Ri0KVFqNF3xY8TWzs2rGhRtXVsQxH9/leLFOOfT81qDGjGDNiyCyb0OCLYFE16xT6KgzqtVXg5/O
iW3Aq2hIbZe/bzbrBNSP5c45xaxZWgH546KontC2KKHS2hY9RXIpiB7ZQ9U5bC4Lr4ux4vXa2goE
OTkApzVa1EhyOenNNRqFPRoAzWf8wk8TP+o/XibAHlt6FXkC+FHWd2Qg3o60t3XSgH2fv3WHLjip
Adh+1Yf43/m75hBKWz4DmlfoWYwDH4Cu5HZCJ2O0kAZ97UDrjnPyfdEQkBCFDaIAgsVHjaqN0b+o
Hg5LXa2ZZZa/AHiEeJ8XZNp8EibRhpFhtIl0SWDNtu3e6Y9fQ8G4ZDtMFVFujNgKd4q17cEiRoSZ
SYOVX+aurIsB+9/3ZI+uc2blDjxJDz5Gxjp8srVNm5QXwti/v4IxcBTeNK2wBFzl1QnrpljzDzIX
PSuwWyCiXFIoQMKZmfQviA4Y6gJYZnUHQd1PXCb6OHBSyq+spD4Jdkoq41z6+ptZLh7JlUUEyuFZ
9ljGd7way3EAQW35qR9xScDlHMUFNxYzDu9zGin0vA4S5GLWT4AoEwICU+lYTu5ApIEEEeSViZYg
7h1h/iNYt9ZvvksrmSMRVHBEOu8ARsmfDqeyiuZa2AgWCPoZ5fk4J5uxbC53yKmNehwupx0U18eb
+D6HM1AopgGEHZKVuVggo123TIYLGtZiClXgelDcI4zEMCotZirO9sjfV6jvi4ahOmbcRhNNfcyt
wD6LRXMkMJqCZxyEj/KvxxmMcSvWtyaqi6rN4WWvQGrkx1iU6SRb97ue/9EZtyKbah/doQLX0Wx5
gEoqEUHAJa29LCjoAcR+5TPYUIDtHFN1yO5JvCXIHNxmnSb9NY8VgdJViJZbsreMXaHLJr3kOvWx
xazlVUHrxfUL2rgI5GxeLV3Bem2y1BLZvSdlCgDBuUnxgYS46IAPDHPfyP6QE3SA3LK53haYSHkM
cZV4ZvSkd4hdVB7GC+8HODb1EzLs330dR6qHBkxwLA/ZM4apuvnDXMWqKSU5kXeeOAfi5J8vW7wY
imkC+dlLqyOCU55xN9p3DYs7cXnYdk8tRtrnbYHYRP9C9OU4q4sy4JiaWHBMloC1nDG34TQ9a2pd
NtNnmItDXn3WvIjwHDNbD9lwzwiMcNp4XtiKfx1hoS3T3oyYW36RziuyM64COyG2X/Jsm9vmm+P9
HDCAwsvqFndP5sYCjDv2jlsjEc6mUEeUyNfZ0ICKumY8M9bpWrj0zRwrpIINL2Rqdu6h9mnIRHjo
WD0DI2kVy0xse0DffHWeLBW/u1oFfajS0mywpnVcr7VYpGeISH01Bm42d8MIN7hA5dxWlpT7P+Dd
JC98k9AYH6J2aYAJ3tt0IBxUaWZuL1dhK6cEOqexLHfOK9inTPlb6wB8723425LZVnHv069tioMu
CfULWHGNLZPdqIHII660VLp3K2/++DQqLAQIw5fbpCVpKRpTTrWtT4ttUwZk/yhJwFmFGquEzUpP
X0Vc34nsRJmJgMf6v9skFisTeblktl3jrbeYVSXJTwiy6FXvAQ22UIB7JFUlB+SVFUzaUf2ssp6b
PlVqUKsJYAf/+A3SJ++cwIxxxPocVwIrxX02rmDPrgOBdxJ7SBqDXBGGtTwwyGyYW3eiutk6GFXT
lVjcfXE5ctLzVhm4j+kYq4QiKiWWLjN2o7bmBg0Y/Syv1INKx+EXTnav9i5BfaQBqJ6HjX8CCudI
eGmDh7rGoFdisNHLi69Yam0rDg0x4ytzxkFoT6Ov+Yo46UB5Y63x7bcmi6lLclACQmnNLg2yfhQu
yDOOkAolRsS8U1j3zs4+0UaNjOl0CkWYvCAf8E1sPoNBTbhyvyfPuTbLStmSbWzc0+4qgpPetXWs
EAjxz2GeuAKLpNU2YygTDMjQt8dychvQD/NY2SHSW3C7/r8rORmJephBvbjiIkMwJk2hRyXDOssI
7NN2ErGj/lL9I58WHOtV4cWDjr6mqF4mj24ylVnJff9gtlUSuE9u30gW0GMmOGtGVoFLk51rxmmp
9bBMU2dHVj6Jymu6a1igm3cjCGGoMRrY+i39RMTOiowH1h5OiEmfBkdKYKScxotI9xKYYJlHWoND
Ojm7rkxOKkgC+vNzcl2k56ibKqfpWFK/a74rIZG5ZRFn7hhq3UB3p/v68Gq83ji4qiEOY6g4M+vu
F+Hc8tm9Ns0p7Dm0vqlHc79kEUeNxUkPGhxz47jhPTsHbJyJcnckac+suwl0F32Ww816YkIfBTOQ
9mkNGTrFXBF6ZZb8AaMBPa9yFPyeqdb/woMWoy7mqGoFuzgxCF05YImR6W94XPg+xR+ZVfZi5TVb
H8kLqUxwW7kwHn0C6RspAIsv4P9umV/iEtYSji0v5qzrrJ7zvtLjlqognIUEkkUXAVIcKlTY0MT7
COqUie9H/4ss4vX85ATgJ7Wg5kMn3V6K79jckquEoVcdcuFDOY4TEXl4awUK65gFnVqAOvergwMi
JFKWMJla9Sgs8qCd17wDSCbQiHEN6frze4ntdvD6SgnezvSX4R4JAVTNKh0s23p8f7XIoSqVgbcf
rXtkfTrqNnvxtTt0YUhI5AiCJfX6JEkA+b5qcgkX//NNWwDX0+mymtHIaOeAJeYze+hZ1m3UqAU/
Z0GPUqMryKaM4BRyWvIAThdtp9GuA6HyxzPwT1vS4hZjKeo+iS1c0eKTk4znuVOsGwlUeET70dpZ
rErxi95nYRJpSCZXL7XvDVVqOI1IQFisOjl21pcLSKf/rhFDdUgZajZWcIlkandTZ9DIshn+upoB
9E3G67KuMVWGvnttvwrHjKj+rL3IcX/nfM6XXVV34Q+SEiBsfXp/H+NPGZIQ2jU9b4aKrMWsVRFb
IbbM63QA5FuppEv5mi1cCxAJcGiwxTH3WXu2rLsPoEpBewGLTp/jJhXwZXsV3r80E1dBcA1GdEe4
SiczVF6UyPDeKxA8fxDDQkZjl9GznE5h2V2pQcUGB1X5/78owoOyUyCPyENjTg+yXegkku3Fo1is
lsC/pQ1atX9+B7urJeAjITI2XiLKEU60zDsEZfUlvQEo3ZRcYOeTwp/KyuslD6Tc5/s2za3tFHK7
7oFTnawW339ZeHXGxpYF5La7sdx4cdgiDEWWNTKsP+I7MhIbw84qv54b/7cVKrC/zhBWvHaDuB81
mt66OYXsCEJgutGDz3HM+4ZatB4hUSgw7H3HYipem04VNZZiH5rqrCgL2AW6crumQeJ5ZvK+VORc
fbWksk+Vv7U8D4ppv/JJO20/ubmkwpQjp7iHLoV3mEWXgCyXY+k1N9lnIgXQHgt9uostrOJ999cF
yrrhKhqUQdFXSqAWrfHKJ/jOPGSq6Gh2i9XyLX/C5qmxBriB9LTgdESPSttSgUqWr0nIOa+eFhOa
Bcq4CYe0jRFduy2OE+5M/w4AM7hhJ45yD7B64gxEdXURWnf/av2wlQtzWTjrFz8piD/yRp6rii/w
kwJPN+FJ7beswk0ZRBvKsl2CLxJwKJtFlZ/XRiuOgCQbWdGA2kZt+cWuiBUqh8mUpz1fA/yZECTK
fbw4Jb57EmzQqrJqpiMolh+c96axQlBYKfbDdOr+VcXvBoclmtF9N1YwNa1lB1ykUAVXRc2z0mVM
r84cbRjgzAku0gR2NEd+cyP4Dl1jrmd2rtlzt7cmJHG1jEpH/DYfMjm6l1MO+0LkfgJYt7nx+66M
dLWut1zDie62/fVa0kpeGSFgSHqUeoYj4V7HO/xSC7gKujKVlJtXgI9ptsq5sHOy9iXXyUnQJDAG
FNlA2pj0q9FMDEEG4b3NlpyRetS0XisyK+busK8CKMVVOFpnNFbqauufuXS/fI33le8QSsQfLCEC
0Yt53rU5ysU866VqMoiWnZmkag1gnq/lJDiVDRYiMykFHPZD1RzwmA2YNQxa4y7GFwcyiZhLdHLo
T07/mqW4WSTJRy0ZlEJlpE/QW43/s3bs/x/3jxC5iz0L/XzJz2QmIsaHF9bl/liySRj/EqFtoOjq
2sAGWGA/o9Gvelnej7kG/e04xQEqaOyw2Emrr9JhckB9HzJ8Nu+K7XHwuv8JlJyxKyPXaa0jP3o4
L/yYDMkE8ptQ2VTGApg/JVfV0HK/XBsqArvMcKNLkiS82UENje09QGoPEKvR++K1u0G5Q/dzQyZw
4VU7c0Zj4boXxlosyxwZytHJ3r1VIRU1ZV2lP5j2otQzeV5LdDGT00BLU98Lr8cRAPXmNarY72g2
HOP5UPK5tC/qqSeIpMPY3wnPfPFgW3fDT5oDN0Bb6YhFtpQikKDbVZxKRZo6ju1XV4EYBSxCYxiR
UhveOJrEB5J62LZVRUJ74QGSgKO81W5oXYhw7BsS5c+12PXfSEmZC1tiAOlF6ttIlZIBm8SIrkTG
hmGozTmxCLWfmemdvdy27Xvsu1RVLeW5d3kNvituQwU40P4ehU3vtMje1kDWpoybTH0gklENjYos
+ki1YF+SnWZ0dZrgspHpl8/KhKoLVGNCm60R27CukdNxQ1+bVCXs/MXrfIXIc1KWDDPsItkjVTII
479LN4OIBWHOIjnfPdTXqKXuWW85Jn04ofksXbFg4/gbxsNAiclImjOSRjQUySflKhDIP9huOkcW
b9iO/PtUEAalYR47er+t34ZC8kEHtfs7C5To9J/oO/+NrOXUxUf4dQHhyCY1aYDWZ4WpdUg/aMKP
YemLLBkonSrM0/dPtbege+g8DkN5ZUCN/SmZKN5vlHgXsPWHqw/DMO6zq5CsLshABRdhZ9YOCeR0
nsWQpLgx/hy8jPku1PWr3y4HMfo6TiUGxShj9oWnXoHUIKi2K/ZCvVqMim6ZRNHuGL/AutoeQiKP
qYkLEGjYULSGf47OvyqEoS+dwcOcsGHrSGmArTRy6zer5zYCaID8OAX7gzI4MEqFf1T88agxFRA/
a8z4fhUxeLb93MJ+/ufdvBx5iQ8V3IgV3AUGV3sWDrmXlrStsE6cibcHRQqfToD1HAOkdcu8G5J4
vPfFP/tsewDbVDZsWWK6M9xW+WNIy/q4YuaEJiV0k83WGxo410fwaKfXhqHk2aWLUidU0KQM/q4b
IMJMHnc+fwRNKXo2psF3aZRhL6dKQ/lAJaD8cBu4nP/4NvoG1KvEihITiSHt0iTKSy2ykhdtX/mQ
es+08LflteW8fYdLeAX76M6HxKrEJPiL2JvmtNIuytTBvZGm3ClpE7+O+BXmOdsjZeGv97sjKY79
Ipgw4mTPTnF4XaLEvyE9MUMuD15PUOZY/r9/XYQNrYWfBE7NOha60w5/JG1J35J/P55ruIpMZMkm
bUpw3H4/ybvztmKetdRZYyn1yc8QBxU4XLf5ZM8gPYlKsC+zSXBu1RjObjIxJlSaITYDSGqc8R7U
EZo39O2LL32TRfTncQ8qpqxF8hZM3a6wzU/aahImIbposBhvN6U/5EGIee/bYFuGTa26t++pg+M9
JqBxwe5wfhalPuu5ejCwqcCj8Obp4+mpkLmVgBswf/dMf3WXw56dyEO0Vv2OQh0XzYuRcqK0yWYN
yeSkEMZdh7eROVL19U9tb0hHsuUv1GaYQljQSUZNXsLdiQhdG+9J4RCiG0fgb9Pijl7DrISjRTM2
jsX71RB6rjbE0LM22zghE12PdNVAlQwIJkSEPRQvNgd/lnOwbWJzdNSZdS6m0wC5ck3D4lTcepj3
vUWnFQYxZE/iqNgygzlPYEwTJASTFdLcKKq6hBKHKP/rAhG3zLtHPfi/tbyP8lAh3UHTU71EDjsz
9mjiOr/NZANNUkwyCpdVY7SdCKOiGsn91/4lGGpaFMEYBbi7CdTA0CFQJVoij3zqwUOH7xrmsyOc
gR2tTHZVpkH9oH6541OFvBIgcZYNWlYPXCn7A9m3VAgILjMUux4r1KvCmFZR1h/C+VknQHxl0r3s
7xdrUILmHo11Ij0Kz1rH0pIMdBfNaxjq1EQ/BDpKQEalYPaK9fafdXR4sDdRvR8nahx8PD268DQH
cYR5hynSpX4Gn+P63iHYdx5jgxfaCRuhWy0fyQGZCEhapi3gZhSgaCUduw8BjUa2UBlCqRDOzTXS
tNWnFWvDmgiV63dYF6aLGuQMU1VZ0zZ3loAX5lS8vrGDpEJlYTLd6clKIwoXF6EVtAYLc7r49Sdg
Y1+DMewsi8xbxTQsTOT+W+0QXytTxZWkxf2hDuUZgvu6CohC73cAj3tzAsv+je9Jnvmwu2K2PGlL
SgLwKxZDMXTWS6xfkU5mw6ix8xZqaoVtEl6iAIh9UDafW3lkBYcAlBMSpi0AIhpz2tJQZT/K9khu
2laQuDzMIr6md2SLeAadwO4681gt37Ax/pVCaQ/nyL6oWapt2o+CSuCEEacA2p8C8KahapsKuwwt
g7P7oQ67FHZ/KyZwRz932rdA4ePMgqgnxQ7xBPvR5hi8D60Geg7B2F2wm2/vPWoact9SVFTFb+Ng
XgP/suKMQlVTDUEAdNOgJP4ZSyvnB1NSelX0wS3oB+47iQlThfRYyvS/ki4OvXNUkmHxuPKPac9K
vwCUAIk4CrdtKJigctTZA0eAacJNixn7vM1C8w315JT5JfST62EM+xpf8mzwXQf98poMLpcgj/db
pnpSpw3H7WRPHWT3gzqcKJNV96AjgN5EASGFn4RxDd09r/ilDsQE3twphUHW3jpK8XJnws3+xbih
lhMfWcFeuFkomWMWxlQbvieQjApMpOuU4X1/xr2SKbikvYs63pcuIjGxyrnPXIOmbKO7kboCIWDR
quYp/kIllul/Z2yMsmIj12mt9S1+sjUq+1MCt1vB70dLBKxOfQvqvRHHcQNO3f1nhD0YXOPPnORm
kPvQhaHg276YNENOcW1g/w7Dzx/nnInlQKxHRemmZXpnwB2ZzLsEcLeOo7OigK1BIgvDFUtABj3I
ByV2svL4L39kZRvcf3tfxSUttQoM6uLk+FVChF4h8uY/8W7w6UfLQ+Rmy2hD8j5vZATu0kby475t
azfgIDZIJtEMXkeceEPPNjAG+iROzhPkvcuVam3yDX7FvyPW6krdx9Wj5gNzGBxkPq77NUEiE4S4
OhXmtVVn+p22+SEdXq/AdRKP2F8xrFGTUkkng7StyIrtEBHnsoDgsY7CQoL0FjlY1c43M4Un3D4i
i73mV4yjoW5wrW8CB8HLrGVHemr7GHas5xMbYAGTposCvEKeuiyH2M+Yoa4yMlSIvYbxKxG6QwlJ
Hf59HscQiOeynKBNxkyt6/sPRivU6G575Vv/7Cu6482EkrvD3TYN+Cb5ooJdh2D5bZs94epd1TTP
IHkT589pcWJKPFai1E3zMeWrJPqEAgcU0hUPpYou9bOgYPoiNUhBWOEWUrLBoTg/kOjV3yYOqqkp
BhCBOR2xVPLH0fYjc35f3TdUJ+cLr5PGQ9i4GlQ7xVd+lghgyiKrom3oDTUSWOE8HrZ1Lq0tfTux
j2ua9cW8RMysQTmZ66JqpB2JLdW6CTSDjkUhgBa/zyETBGhAEt46rgXWRE6BROfhOMRLRmroi2r0
AP2UaAPs7af7Q8Qv94fIvuO7hkLU7xU3qxvxDZA7TCIhD50ctPo1o1fYVTQ5V/oB1EBsY61Bveve
ZKJs47iK5mqe3G/AltDDcQIRmsywj8lKJkTuERbyKxe60VYHKFS0feaZEBFNghWs7hhqpOlfQUCf
QpRvIAPQLSCbT5N6zWCL69fpGj761gOKoWMJ8eFAXUn1yOgfD9O07ZPATsvk6d7i285LN2BUBnqM
zalSj5e+fGC90/hkQknZFSI1qXGbx5zeJFYpXGfpYQiat5H3lHNqEzeL23oeUIljPWQppXe2lOv1
y8hdfjobLjwuSkFBlcb0u4jG8jZfG74FqKCHUkIefRu1t7q865yerODPwNCNOeTRnwk7OSEgXvvO
vDPzleoKDiuYRWLjifBe9e63DFHXGLDE0J0vL3F7o+vFUurfq94QLk+3mihiwzmajjxMaxkt7RDD
ZdzdMS9DJQnLa6NtS7/9uc4AQGyEwm1ohsr/P8yx2XFpf7Pov8ERxvlTWQoo8LWu2Uj7bvOLJLoB
Zlhwx4KplUK/ry6QhzS+jczoe5NHHm6UOgrhLULGq2Le/dUvYmd+JGkxJTcRhPR/eDM2/bpzasc5
y7sVzAzSjx2H5wMZMmui9PsxM5gXtjUXxlFzDjy/MeDnvSq4yL+NyVnDraxuTpSdDXHYOM0vGWZj
LKyi6UIE4kDuw4v2q3LRBO+t/AgxgOF9SolSE/ts2kFbdo9CceQJR0ogMruF7vXKuOjC09Uv0tRn
KoZrkqMRJkzYkG6mEFKNfnENF1R2tiT6j7CKSKUSmlWrioxGYXibIF6MDWOxstOBuxxQiwuxd1sW
SZOPxhggg4LJ1BzPvkl2+9Gek7k/iBYLjGgZa6eCEBm8DPInfMAnl8WtonjNP8GlvJtYBwc6CQtA
MIwOtvTV8wZ4InH8v9dcZSQQYDiD4IjLbf3+oVy1hEKnTRuxJQnA+3dll+gVQTP1c4KHX0L92m7c
/qIB1Y6kqVaD5QBNcO3Odx8UysMm8HSOmMmih53Gymk4AZ9gDxfkxANlOZlZIIiijel5VHl8Svu2
i0mwpzhbVx2UW4Jxer9fx6OWGuZD+K/9LTfUi5wUKpa852lhFyn0X3HS4R0ZxhoI5qpexK96tR7D
pInkdPXQ84Tkz47e5J0FAUbmOoYcQYBVPNDqGLoUu5BqGActrv20yAfCb4gEvcyvMnAgHuj8fDU2
rUK2xAs8eT1pa0BUy4+mrmzKA8MPc20kRQb74c8adZruYgc0QhwLdClbBMow2R4PYgFyQFQL6z0D
OdQAkYJwOAu2Qs30KYGPQdfQiXtwe0RfQTZeVQ2wfaSXpBkswYRLVEw98SxdX6ytvO8qdkB1K2tj
Aw6TwVNRaqetMmlfh+1a3e4qkVruLHB25w++a8KvCrFDyEORy0lTz6mKWq4sNYjkolXLgwK1s6ZH
Hs6NOdA6Y09DCRcN6prkPKLtGIuIvo+Wcaat7kD9KpW/riPfmW6q+QTs+tKXL7wGWqvYrvUfghXA
ycMXtm+afsYkluswMrZTMEt0i6LGo4ZDhJFQL9mP/6edvttafEq/6l5pxg63LvvUefCSlfnq+dal
8JBaWFyDJf6sOsOYD3axuvnWcxbF5TWsQ+BSWDlOaGqZdWGdB3zkDhMfcCgROgpLyR0/VucqRQ8f
Objd60hWBUe3+hebvvHBaTZeH52sE01fLKNMd33lA9N/Nr11fxfPJYAxVaXP/+qDlUAA4YMUVOdz
GFVWmpm1lnEUv3hKchsUXctrdoK2WZCWq58nNE9pNNZJ5fNp27LYdEwe2zvEic3iAnZOchWJaG09
kk8JbDm/gfGNd70p7t3JHqdLpzQkf4ZcmEqrwswal17zGuuoqRIiT7gdckdweSTXA8p69OEZw1uv
hPTlTpea9J7rlAL+LFYmUj8xpvKqQlGTHRQ/+C88Luudt4S18ufabgAS6oGYCPBNhcdeWcszdR5k
3ri7PWDMlY30n+URH5RI0jtY/A9jliSUOrjxzA7pgAGr3CM+sq0JH8DRTDgf+GH5j4TYquqr6EKx
6No0oVSXbfPEfvodfSC1JwTkZZkGfL7ysHiTWgmMxR6C0EgXkBoY+tzYj8KgxBDHt5SD+6GEcAsa
ve+MWbYUEdw4fz8+GrCMInWzqloqYxqwjd94dyMKDe9mOPW9WCeQg3fo5aMkFHexPQkH4KAX9V2S
QtXUsuSUDWeAL9m5TVyRp/PxVensqckK3DGxTvDd3X+ItFxZwAb5quw9cJj0HvKZ8zUpr9Bdw1zt
W81mL9eLgINKjH5BUvZpfuSaH0/RrIaSzYTrPooDrw5VdFbHMEId/DtZfADhCPTKS/ahssNEpo9t
IIk1iZqs5hIQvBc7RwDVMOxt+gYlgG2zsq+RXdp1VHR0eR9T5Bhxr3Yq1HCD6buqOyaA4Z1wCGB2
xspOfMlzjsZ/3BC2/AVF2qb2wqUvUEhGqYv76Rzavzd6jHUHnFQCF868qkcQFvLvI2UDkqEuSzZa
/ifiE1hbxI/GZjVo0qZxRYFBlawq6wuzlTCiiBUKoJ+S9h/LuO7vyk6Ot0KQCMB2vRBHivvrBLKq
jJbqcXdM87izKhrtqOl06P8RGwijltmrXoVjfdJ+3+SXCaLLAVmdE65zop7sn03kxpirGXzr9rRF
IMhwmr0R4RTz5u/uMGAModXfR842N2O6X66FG+ltZToDelF4fhAPwbQy3XXKriSVT/VRJGMnt20h
2ZztXWV2uI6aBI324a4oS/4A+mRj9VhM4K6TcO0Fw5XLOjrdBM3j46v4FeNmevOZdsdK9ufr7L84
y5LHam/r2Z50nbJn/BiManJ6+LNgh6g8at/cF0ZE0Cu+hqook+bgG8ZgyHH98p6PUX1yBAi0aw8O
OIjMfssaXu2i+44qwkU8qeiqEbXW7USuP8juXm5iNnY0/V2DBFjWP2jYQI8N3lV6DZvRInpGDbzh
FV+wF85jGlovAo+PznBYIs3+WYeurNhtnZ0ITRPWT84ugIIBi3EBLiyCD8gMXLK1gteKPLhoxaeR
MWn05WXqQInPuPsJYigxHzsd3QO1WB8yqJ7wf4/w5+RN/ZqGyC2q20yPF9DuRwjhrBbaIEIairx3
yDpqSBdnMiM3PWQzwt5G9C/EA/l4ePJ9xUKaWAhU0BN9xn5IwmzYegjoTOw+twLdbXaG4ZfJdvtr
UxtCZknxOWGXKvZU7T3XyTcduEO/ZZJt1iRo329ctMGo2YGRCPiP9mmXg27ItRoPrSudmCVXUEab
aCrSxB0pEpd91SVXqUdpzdVDYVRUV2TxdlLvp/ZLEoaKRUWCe5jIRrjR7ja5M8AkPrI6cmUucAuO
rWDZHQaY7o2M9itFAnjCbI7zlJCxPwonOmkKhMYitalit+4Bg9WZDoVHtpPuvPAWpwJipD/xBLA8
IMJ2NBQNVeYHbiPGvw6D5+jTM6GxEAha3PVhnZ+LQj2LE53c8SEmMTeIrOWTC+3mzOL57lM15bIt
A/6Uh21LlspIvoQ7ve/TSE3sBDOcqV/ma/MQ6McnbH8AlX7HRtKDU7jL25QIDmG9aK0kh8Ee3N4A
rH6MOtWN5lpNoPhNgt4uykywO9DpM3Y3RLJOT6Du0R38CEQz91mxbyGJ0a3Iux4aPH0ziOt5FNrC
EJdyuIVHmvwIvSoxcJHS0+KO5JpZ/aQRX4rOnpWPMZq3UU7irIpFm+byJLTt68uj9hHLJ9oQwMcq
t6NcF6LYa9h7WcYKFpPHWBrwy8kwa6O9RWTmacFLSMkmgtQZpfoNGzoxO77tVZ1xBxzDXpVRkrrL
IDBWEQwBPLjTvsGbsyjmSlge2nqNIkOKiol7PyoJMk5NGP1RrLf9zvm2Y/K7/dFs6SdnywsobhhJ
R5e2XVEpDy3UANeRc5n7qa/XvMUxkQXY6cuNd3FAth6k50+v7YV2oZli23Sd70vAwW5tnQ/HrD5h
WZkBCLARfG3JgqTKP/+RMtLYJ2j/rUHRwe7+il8osDnE1MIpg5iHYwstOcgN4myUgYivGS8QOU2B
XitUAC2AY1fb0w6w1MCzdcFDzsnBflRESu8lViSHa5Th7hA8vfIl/ib6q9CEjq0SlZUbd85DwrZV
queTu6LoFNAuiF+rEq0CY55fwkw984Ku5oclD43QsWiyvFjz7sAWhCBx5QYy3mKpQK3sy7Smling
TVGZIYb+P5swE33Q17OYYImPW1gkOS0ovhs2dAKhM0TDR+TzQlKAb5mMuLDNMawNlmiKENpdg56L
0btKJG5V2TIbAri0xg0Fbg2ZZ8UDwJ+P3KB6GknlSJk1Ozs8HCYtXC6jiH6FHV20ba38KZKdkHUs
ulC1QnR7Yu7lgiPps1Zzeb9p54NgfFpFxF+L2hXRHhhhtiLsY6BGU4OOfQNYYTeLNX44sejTPuXq
43xJi7o3+FDo5h088wJ+5jyFwLbtvmJdPQm+RvXKC/7zdWPBRH4MjDrhZbR2vCU80IntefEWMVaT
s9/+V4wqzJ/xWdVJncfMVyRs22IV8aQQ+3P3HiFymxW+tmwRZALqbA8TKmnYRioTrt4xCianbY5q
xRXIFLVMSvM1/YYdgZFSQu+kGpOuRJjkfJq9vtTQfNt6JsnaXT1ji+SXjIch68VquTTbokszg4JA
VACB347QbC3qFawOFCxLtuNG9ojUey0zupD97dH6xT7kfuafvc8V8Palf5BrdhawqrLnJ6UJKK9i
Vw+PUYWvcGsFhWy1f2ylHRxrm1KeUubHAz74F5QG2E8EgXyTs5RH3BV72dNqj2zh80BfSFMpLdnw
3nbQDRZp333m7a0FOwm0DimbOUxFTnu+y3mukUGrXyIdfTb08bMI5+KqKN4qfSmDEc4ZMdbP3AGV
EEzKRIhLM0sT+h03381ZeoF5wSnB5QfO1CSusZpEXJICaJ5eykSQIJjq5/79dctv4d7oFonm8m0S
Eo3yaNzYRQeKNJKlyHRqQVWEX94ZQQ1tZomt9DMaUcBFx4MIz9q6KMrFK0ZCpHPT8LkWLzpSuFNv
RAAzWozop7ME6TMpoou3vYPboaC+TCkWSP6fwpxxXswLouERgl4iJJP3rRjLW+mRuB85ZadnyINE
gvfSk9Sg81jtFagEg0LtQD488uDc/kBDtnMeD8A7xS3FhC3GSy8gR0N7nxGiKQCZUInYIabfVgIx
IMTmvMD4PHZSjh711HOjJbqtuALeWzOEkgpdrOx39FswBfCDPWVO9v34R/wSz3QuVtOJkGpCfFOH
aZFRoWA7SyjTYV7RzbrdMU4OWB96xmbRLpVZMyK7KTqVFpzhlABjn+M+5AsfZvC+08NQ7YPgV+ST
5qpH4MCIjneMQMTD0qsvuH0EpYpqConRFH1+dJXSnfVumjd7cu76xZysDLUShNxEJEyExlIQUEDh
HifBuAy0LdzbdGUugSs5K5AAmnR6pvo4taJh/1PZfw6yoNhbZ6dCpk423Q+eFpoIktge4I7QijDV
vd5SgbhONhgoFfUGCm6OJ4y4e96jSx1Gw7JodiI4cSQ9orgwZFyFbgTJOJMjgQuX3RtyhGTPh3+z
FxMb89eYijCBWhP3eNErzdwy21/pVwhOiYncBQ+X7PXeKClnDzVwaM2JaJvMgwQFlAjA+LYaoArU
PqeNwVnfd5I7pA4G5gfsU53hqlK1wFg80a9hpHNHe5tEdwjSOU1Qt28MyU5vQFH+1q0OQCakr+uV
WLb7XTwUamNLgE66a8TdikfTFd3SunqBMwX6Sv0SZdpyOoLRZbL+CHr4tqMbUXY/cfIq+4BiSshd
Ef/Af3mUmrYsvLirLLkG/9OpqnqtNN/yBH0YahvUvW7zp1TLCNB9mKTLKx5r6o2EySpDwYdKQsOG
cp51Dhi2L2h3cAFBPrSZ8JOS2ZM8N+q/EzQd5aLU685tmHkTaWIQz16ZmQluMIsmSsigMexSTLxG
O/rRQCyQ0/HVtTzsmZ5zWw1kGj8t5rmChq8uoRWLMJfptkUOFAJTqemaVRS06OsHmKuXWLy6bbmN
xSJTYn9LGuOILQPh2rUP5CF/97J/nnHIAe+MhRKkVYE2y6XJ3kniB1tunaKvjPLzxbRyyfdBjixj
mXi8DxBMd3FacTS6Wz9WpjTjeTb59ff8K7narIq3vCtn2henvWDpQv3Lxi1MTWl4Bn8g5E7fv9x7
wJY4tSP0C+VnB9mmFcrwYV04ABrUBFNnlIMcyJk/KPW4+cIE6MkvIHPnjUJcCKeVk6KQiMy44/vM
aTPGkDxtWpb9MMKxzv5gTV08SqRmTsf7z7YvYc+OyvbQEDfBEhohOdOXDrTD0PFR89zRyrjlTAbx
upCZe2LCUsxsgOdMpegXTEHhmXCgNU9TcAsg4UkX6yB+qMfmMYvD6uXRrgW1oKKuPK/Y/KOCmx/b
D4PS1WVX/PQBgcqPj+Y17Sq9lZgcu0mbft/qDOLTf4AFEp26IYDH0bSgGC/7IzDfhC7XMQ2ajVao
TnbihdxHdrse9ytM19HocF2KHonbG+Cjo1xOIvtA9hm9Seagxvbjh0Z91dQd8qKRVRDCVKKoZyT1
cti3G6VJ1tR+mh//jlQCSXZWQolZRQFAsM7lp/vDrK+gpze/HOm/ZrlGgX8ZKpeypkSIeiMSMWh9
I254Z/xKH6iVlTYmYr2bFFDwiXZi3VVsZFqoFH+JY9TvyVYMHb2DgXE5ZwkliWVk1vLT2mwr5wLi
gXSNjdHPG24cjnovlfcxt3nk7yG5dv7rG2vcSqI/rpKaNpKQMczLJG2V92QFcqV6zdmBPusBmDEo
9UoEuT+wqXet6W8XpJmGewMyacMRSoepSmDvldWoeTqe1O3xw2scwtAPNJz0ZIgJ7q+2SLjcCgKH
x90TEfWR0GWqz0Bv28K1cC8VdUKcRWO3XNbh21+rfjfYLsxcS1/LD1MNeHvxPt8ZlWUbauTych1R
YMhejP+fEurhVRdYsTX7b9sK4+eWwNLViCrfWu1jExTwICWDtNkPWIBAxgbBGDoVQwRCR2x8/Iho
JKtVf9t65cM9tdtSzuYqxYvbo+XF8nfBtvP6kaiOo3FPMfTiwZuRwhZYEjsP7iOR6SDDkbdV6X/U
zpUQgLgDvuyYYVwI3P2AfSV/M/TJyb0sxmpfIuq8HgC8NWElNW2KtpRokbbnS4hSuh40vQy+MjNE
r7sYu94xfbvYuOEQhWH/Hucx+ej0pzsbSj1KPG8pOU++3rrRTgAx/N4CbVpbDN7axEpGyF2ajUCT
+Axt/cndnAnd60rdXLfJhNz/KU711rgz1Eh2ips7XHxsFBHJxZP1ubu7pvub/ba1lpvh5NDL4cbz
LOlES2L3oZsEarNsedYGQoQvoeoYrmdoTKg3WTqxhwK8lclTvVLsxByfi0weQ7S1bOqCtx7rwLAh
zRq1kU/gXQzHPzc5xjM1Y1TNGP5wfH462iQNWqzKdpqF3zSfJw3nFNTh5HLvq1lU19hYJLDCwcwc
OxPD4kdv7o3FUMes3DEuU2f2gq5C9ar3Y5SyrY8G33UFAyXsCCbnpfe893xCGOjmkPyfP+LJg1uk
losigHdf/GHgE+Se1jJjP36a+Up12G39JLBW1JYsajy/QChQgi+BgSGp7Mo3JQNoB0ut5Id/DSZT
/62iIB13rfMrBDcojo+lgdqiIokeP+vdPx15pyq40Aan4g3ULtqAKhmZ4N1zY8eHxJ3m7MUvC2vW
/M+CH7pqSYwqAMy8Jb9f6KVG+mAIKdCrvIvMHbpgmjGsF7y4SSP1DuBYmGXbdQbqWTX7GswiIvuA
L+8yXI6ali1P6VPJV6o+4Yb4MBTvGmFOeoAarAsyHLZ7onXSNG7DRXTfHcf82CmIZgKF4LItiAso
vPycGruh0l2iCBUZ35HlvTMucYK1SXzkV8FW0YxgZa0FsO+SlEezkBX7qKqGi6LQH4IHP5aL4WV1
QeeKLsnO6BWtKQrngO+aqUbGbvkThOz4FHUtHsGyPaHqFne2vPX7Lhp4hipPiafwRFzDBbEYU4uH
uPSs3lFrwM5/WKaIzVKjwWBUcaoCk2iJegOMFhrDb3AnpYSsz+Ijd8UM7XxhEg0qoJlE43ITe8lO
QPxuHUF5vIoyBUB0iQBAivt6OUPWiLw98UHeH7dnDHAhI4BMJHJ0XYm2f1SIAIJoW5p10D9RcWzw
pmbaqizdI4meY40vlyo/Oc9PAlwQ4YqueX40CzHbZ7e9BhQhYmUcCkvWVI4V/2NXKBHFRkITRS7J
ONkQZKIDsNnO/TYqkT/12IlK3TSsS01xODC07v2/bFtiSiC+Gxy1A1gWx7DLnPTFl3xkznFNt48n
1Yed77HtoC2VUbgljjkmNVaoyqMNhT4755XozcvHqQKb7aYpivbqKQzYd9xRz3E1pzVB8W0jCwJg
azwqV9sXhT2k9aQjeCU5nnLMM6YieI1+cAFXxys+U5oWUb2MYhdN64J0PHXrhU7w3K+fD1G+4nJX
pWc9Ay8u+yiY7OXOjs4Kb3H9lh9TEkNS8hMgEswQMjDeOyPE7E14qWyjbUwNboJ+AeDyRG4rKaEO
C0zFoEoMYmJK3IL8mC79NLo6I7xSbeXbOZLdYPBIeKt29NOqa6CqhHMSzSDHTFoTl4LPKJpB4YMM
0eDBIu+hHYvFMnwTPsOsdEiIkHR8VgZAfXajbedFX+t0ALI1JrAvsLRWz1Fy5eaStk4bPKCzxFB5
oHTH+isT9Qms9cBLjXd92QUL4oy8ygTGuTP/RjFop4S59nfEXHI1xyTutG4qz0dtKxCIZMMbNGZ9
22IFINdpazYT1rFdiwd6aSdjAkGvmYOY2EoZjKZWi1jJLay4FvG1mNaUBON7kYjqVSFFXRlMXiyO
dQTNxQVZmCSF8XCeJdnwZQiDyzEd7dkqxMONyUnkOhzf6aSb/dYfFHOR6NctXEgkb1GSwmHMdTR1
MSauSy4K/F1461FriMjLLYr0HjxVsGTBlqBZgRTmi9HZA6p4Jeq3rtYAQ33pyzm1MIV/91VS/eD8
CPuA26kmv/vtBtd/5rfaj57qGdCsK2Pt9vhJh+H84O8Ca3Cm9IIvehdCs7gIPqvWCxh0luqZmWN1
3b6We9gmtskM6vh/lc6gGJ8sLN1S/VLzD4a+yVeWfW/kn6BG6XYQvrWREUTg3SuX0Av9bEJAUULw
NOfrF/sHZU+iI0vWj6iIeyFMayv52TD1vD9hQF2iu04WZQ2GCGXlsjJFTRhK1Dt++Qe7PnIFXO2B
bBjtoi65vfPbqI1fqjQH/nUx0WvDFNF6TC7uI3qrGf0sSK2xUHvQ241vYwPkOVeO9b4piToc+y2P
+1Op3XmmkwklIlqXdm4XHSjulfmJspgXDNzmhnoCnrOMkjCDZyRRjZPrEyj+9i5+t9VgIxX0zoH6
r1l8hSjV4y2SRy4ATAEbQjBQ2HCJ8SEnnytUnKhwXQ2WThEAeRXGryRf5MBkrAOnj8c3YIT2+kuD
vFaI7d51wPWt2E+qBq2QU7HE/B+YMTU4FNysJcWKrWXjgH60IxSXMJTEHmBDrhbp9I6cVu0Q6ruz
f2FQGb7a4Z0xMpJnan8bHJMVU272M41r4K33IiC4FiLse+1d7LB7cjgmyc8ttIMdJstIknCUMxCX
hQ8taSKq4UzTijwCGsQXSCGMYIJwhOCyHA8qpdDvZCctJyQYBWk3jaCuie+8iqgenasQBFl71dWE
yiqpCBuP1y/nm+gVJ2Sc1HNEbrIHG6fYxdeFWMBDblbyO2/KNgwC6eQKrIZdv3DO5nOqFbnevKkQ
YNdsIftTjB/vAM69QK589KZXKg9QiKAtUqeWZMw7Bbbf6qUufmdm3FHN528Q0tOuCSK7xWCMdkLD
s57vLM5+4RhpICzZ/5OlUKPoKdYefP+kKpkgIu1tpdUKCy0xN7zQv4ipjYDkhCWryMkCyR2EfkMN
w5QeK3CxXprPNJrVYJoNnnS+knSbih8RmT0c3oGyhW53bjqAXD73L18KuJLI3ZyniazToSzXhAoy
y5CNsaV3CtDFSiRCxOnHFJKgLeIyK7sKXGmQXoUxZ7meIYxdzQQK6qgf4o01lQb4ITXtkaJthYwe
AZywDCT+OUMpIFvEHjEtm0eU88g8naN8pIPaTSEABv8i76uuq7bF1n5b0AJAC2y9R6QFR9878Ou4
+F93oi2YPJAY9Gr3XMD2OZWH+JHFXMmD85ht40aAgQ/kmNks5xGfRzbEy8X/MyMO5Q3iJIXZmw3G
uZKWPfyFWFemVJLPtmfUm+yOpqBu+cOgwLVmruiCvXpZP9728XxG1IEsX99Op/qcCKfHyUc91a0g
jEGQPAA83yFMyvTWJ4EUXSVPdo/7LddC0doj7yXGlbONx38a+iM8XaJmuB1EiPJuruA1JDf3NqaM
5xv4Qu7HczZ/oOpHHo2B/KGWKR7bF+lHvFXvCGuaURL0EVDu+nEpe8jUomOCvUlwqiBWk+ZS12lM
HM4YMbYevCPxReSvPa5FxkfY/49uhDf1XM6iBFAkB9XFJza1RxunusB4oU47BRuKEVFR5LInB6t1
rPEvpqQB32/kWEtgca2DO9zWfbE/WHp9qZqO9O525IgZ8XWnvdM7cR0IALM1SIcOAgRq+uy6NO4X
mI5vyrgJafrVeVNsSJVV7FeDEuHfEUtdpr6IrgIGgGHdAeK7c8/jSudPtgGoOFPTYiIfBR2sLbup
z0I+2y01cRatyLTVScAdtojoppMJ4nRElsap6F3wgloF41L61OEzgFZ9qSPCb0nfKJoM5sn5eOVZ
vUdkIeCUPKUcTF0a70gMTWYD2GU6Q/4o/en+l5aILhBw3bh4bUA604SvZLWYzVsRq4ZmI4jz06p/
JDEjJC5HQVPfA6EpWNZ4t1HrXtFpKxBdUAqCSZf6qCppp0xihvFjvnoVkp4stQyDinrseyjK1hqC
R8VY/fq4Ny3yRM01rJggXH0HCf+iKKsKsOXOnJoQZfQKOuB9qv0q3DRwaguCALgEIf3z2NorDfIB
gafoDoOQ9PX1fRzqzayX9d0fymiWrPWHnC3Gj7PTQcfzJPbucO5kJR2vQyohsfNoeMZWXL8Xak8K
8Dbr40jLfJ58SDaTX6YrBUKn+6QebxAQAd/5XgTpHvnQI5F1Lt/cH69znRwFnEwrm3JNIr8nA4Na
44JbiXJc8g3h7EyIWrYdrl3j5es5X+4h2ijJJU2QL2vK1+fE6Fk79w8ECqMbOG5pbh1JZ4JNSYLo
2GGfHYAlNrrAFqTCBi4NlYWhy7sYhorx6I9OgHKoVIWuX11gUzI62NwqGdvIqluazhmtou/R2/Nw
7htHIdSqFmfpOgp9MUqt+LqFwb9bUWxbIPttWGbaYjej7sJhhoh410ijFmErPJOrOv+HHCVh3eIY
VS9W5JF90YFMEfSxSlatw+ME4ZqoIEvcGGkoY4OSH1yX6HPV2cu5y4mBj8JS38S9vo9YMxfRvgqS
9cj8Jx5ZicgtZtWGwMRRMtuSOsyTqhStkabhIlwS8tf1t+MReyZ7xaxy4fhlDQLEiDIpDuy13SuO
xNyKPuao6Xc1C7mNhgZzLylT35XoMUxP6Bz80CPKVKjL2jtTnZY8i9GB7OO9vPR8EcKHi/v5xtH4
oqWpIG9Omtncqfdx/esYLitBjBe+FbhG73Ec+0aXthNK1Nm2N/4xesJPGhhcdrK3/gkl8G4MhHnr
dyCnRiAzEffd6SrKYKiepfAsJPV6bCbW+qibxl7BHPY/Mb3awQvCRrWmiBgWQE9bg7Zoz5N0dejc
8kIK46j9hmjGHLYItAXRmxxlcKKlGaYwAwRBNJik3e+op68aaVH3ZrxjGcm3HA6XBlNNS6EuCrwb
6dLuhcKkndI8E9SdFvERzTp/gBucEPPYme3U5EywyUx30vyFxGTKvEz4/QG8hu9VXwwNV3dJOgCX
KsrBmFTHqIIMONAR4jA1sDKArmfD3FWahCcOdY/+Khm8RoDoP18nmOTHZWiThCHGsnYzMSUEhpEV
fVyZlIWqJE5eDk26vUG/kII30Txp8kfUqnFAqjhoGN5i0a/qID4RT9eSFF5SUZCvT/D4upCcG7vz
xKXGelZ1AqeLn01yJN9PXaW7cQwn8kK0cFeazb6s/3LybH6WQdcQa8yfySpIN4XGwF/2nqXdgrla
HwsxGo0jHPd+cLtAixIMLBjGm8Vgm2v/mzhwHO0sn3uvOqQvrBzguHiB0rwGXAE6XMqloJs8x3VC
XhmqNE6yqleNutESroY4r6X+S+6FTB7qcnrNWmj6BvsynCTITMi/wjBd0ZNPRCSqYhjgY3op+jCX
ocukSklp8XRzZ6M07dbPxjeAPXu4LvqyfKp3wNcOuH1FO3s/DeGoknhKx+y4SFISsPgN/ZNRCR8E
S4N54k1the9hPCRkEY1v/fb6R/8G7G/jwmy4Lz5VgHSWY9FlBqiWuCdEiD7cZzzSp54F3iWEjQBB
AJR47uOr/VqezOIeWQadRm3Na02hkzTIUaGssDtlfnlvNHr7bg9gCUUpWw/S+vHFfkaYXV291hEK
udqHaMSTIbl4JTuKoMQaN02YffIW06rYv7qudMDRkpEXWSCtYruL0sI2LLMjZ5c+I3z9ifjmGohs
kGWYNulz0Rs/+vKpC++MHNN88SGbOyhuBF/Vl9hTR648TAUwCIrLSKKTysy8EeisN2bGSfmJd7EG
qglQSE/qgO+0IpF4OG4MZQVgDdMn+/9dL/DBjb7pgB2k4S1om1XwzvpnkRnY44GcYNqMUUn2GzZC
62/dFrzwef5LP+Mnooe+jEnNKdy+YtGXe+tBvZOcaPK2NwtBJSwN3ANkEIv1PnlSP7ZwpHU3aU0r
ZqMRSVA92nsXw/8P1BHvAp5srWozCaS3Uwapo/1ireKV+UQ1Zb4xXjA4uyBaQsyVpGqYEkY29A6k
uvoC8F9a/Gm4lwpzOBsKyFQBcCCZJa7SLpXKDD6nqqZbtlPIU6ybRudnByX76beCkQOJMPJ0QOXX
HIdgjPcx2caxnJBK2UZ1oUFYosXjoTkTq86yocYJiBmvkbOqP8b10PldTI++wWrFL44/A8TaCr4n
q3y5hqx9J9DnG+PkeJ9aL1FosckwHhYTVwKANVu3vPavcBmqaBjCthx+idWKgfZIpUynC0rDCV8g
VMSNR+5mvRYbXTpG5tob7Vqg0x2KW3hLl1vmQEKgl4jZPh9PkE8tV3N1+7YnEDOqPtufdO2ZKRfZ
Wb/HE0KykkTMD3VKT6xf6njrYARJoaoVeAfSHtuf+Tx/an4QWDxQwqCWAACzrAB49MxaBVEhIj3R
X1MT1e6vFneH0v+9tGOygBabVN30XRIhCDZRp22p3SU5R5IdzWs3h5JIhRBua3YU81Khwi46Sauy
5T+hcTFGEJEf22s16RtONds2DdXWjHeHRezL4AIGe9Js4Q+jxUpT1LtowhUD81D7JbwfOMkSl3/M
jOBoRCGl4NKWBfK96kDxjxmFW3HY5HprDdp5ezVj94en3+mdDRiaszK+ZZYHhx9kt7zQXnPMzXOZ
lZlSZ5DgLG6He6zSKheE/22fcx0KdLgtn3UjHR0ITPMuWJvBxLU4H9Dwv/OXpzF7ZkaqaufF7g5y
cxqLFozPMMQqadvx/oTtJpvMtp5WJONEWrWUf8nAeIExyeF/vhB6jWzMdCVuT5GgiTLoCyWncwy+
oUqH5YhTO/5gSkqUd4Qd+d431ibwhcZ+ooEH8biTgB932um2GWS7E8XpvrU9rk2fmjYBlxWgz+dT
Q5yFSpd74opx4Vmr/NrxqX0LKoJVySEayAOFFnja9HwweL/Rl5RqSCru8Vwdok3cQEhMP/2QLzou
17y9ftoqs24fAAX3akkMPQWVjEeVbda5AD2z9/wZ0OdjEc62AGRHd1l9Y1KhEvL3dU5UD3h4tl/h
O1N+XpkJUXdDUJ3JiFBKsFEltdn7Z59r0x9gu9LdNy4tSoFnMwc6cPuxXsvaph7HTnPMkX7EhYGy
fvfd3dcQc59RbvxBxXTZ/0LjlZIXeD6TbNohggE+XczNsfJu+rvnLLx/WFnFoq4nGsiUMvAMJTtn
BG8U6ED/DoepVuHln4A3uWpaEHw/CJW8aAACTwqTW1VCsLcuibTc5OwFdauxDWJy8coApj1IEzcl
A8jbwCgAKdWj6wUK9vYjCNIWgNbFIx8stETz1QOiRZ+brCQAX6U7B/58g/Zq3qCt37en0fZKvbCG
HOYL1M4w2qc02cVqev056cVO6B98rpXuxDXPWVSOGhqOsk013rNQexbAIOD8RmkPxGICU7z6oxNk
NR2xQmhJuvx0pthioVMuQnpeeiSvZ7smjvDg+BuUlo2V+Kb3Ogu8FD+JGkUtVQV+1BiYCJsSmrkN
jMP3lQ+TeEroos52XZmyPP4D94QjCo8v8Xlxpef8A/GDJdwtq2lx7xSKOs2aCfEVAiEo4y1UN4h9
F+ytDq6tgqabNwIYG2sHqJAZ3C7eFHqAhzwSlk1EAX0FTXfeuM7VZ7SjabvfKVh+HGyEu03bGGmY
YgOqrz0wqXV1K5TbeuudxLUEixFgf2b1Iq1y83T/WnNLDbwQI++X1ezoMXYSSasA/o7MhLZMMSMj
mDfyDI9si1kKTz6yItsoxW58eRHp/1JWHQHCBNu1ZQAk7JD4THtP8v+Smef899COeiwcomyXGerA
1Q8/tLmROfS320/CO+Y1nQF9LtWRXdYC8jCqqVEmOPxBL09Ag0s58UYb4EHczg+imQmYa7ZKiXhU
srHeg35LpyGbQ1qNVCE3c7B5e/SQuObs1mNx8qttmfAv01cfeQXKCMn9FPdczEzDCoAXDsAUbM+0
V4PISNzZpdbSc713xDximd6Zxdm4cGu9z1dOvtMBxLx6CZI9JxOVbPuuKclOYUZj00UozSEUHYxA
PEu0EAOjUWQ2KlpQ5ZFvlm2Ue+CTHcnCkXRvKOOPAaVObtMj+kGAUkGZ4HlQ/zsQI//RqFD+6r/0
gyho+0BoZaWLP7Wm4sYeRXUQIpWnVQsn24E53a4/HBOnoy7yszpHbH4hgjNnh2ncqcU0Kbd41FLU
swsaCd6awCmowfe9fLnuX6yCMxtwggv1qUbzNlUpgooUnr7X2Mgx+W+CHV+5fIhpUspzhRZ38mDD
UwtX4EIf36kpQ29iw8ScveJCCFwoSv/tm1HNN79AyNFSUk8iKoKDYgDdrO3bMHytEHnZXfMHffVg
7CxOFBmYebSnSRxoFIgrxZbJwO6NwKQw/KPqJWrl5r6l4OOJNDB26aVUQfhcrJrANgq+NGFPQKm8
xNiVcMa9Ys8Vnekn13svI9vBiaz8Fq49+SgAVpvmDMsuozgIX9oDRSyFwreXbGeMI/ncTRsuNEE0
v7Ip8MsGb5TU7wBsNDlx2sGGxlR5oQVFLrsKjsTcN8zBiwikfa07hymtlt5sLee1wPT/CuySvkbo
IIqfiez5nZU35jhhL757a+RPn+2wvn69h0Rz7n99dvDeLTReEbyQ0UbVQM2v+S9M//zT3go7pm9r
DeoCRJFw9HQ/4jjkGxt+TF1HkoNKaWfWtlSlcJi4nvMkSywOytryLjqSK1zMuTY7BEye7SsdEp+w
RR8Cqku/SMNqwiiExPHhB7HPm2KCUUt+WY9kwIHwGxsETrgzF2F+v1v0IbnbDMj+cSS7eoVWefi5
Ww1veWm4QELRNM5UoSxCbJyJljI46quQfPONNV6uUTyryz3+Ugmx2x/lTmoLpF0hCfW8PW0aKY7J
4tT6pXLjTTt8VsBrWdkFqj+d6aUE9rlcbtjoCayDhTok79D1NMFMrdkE2aVA2ao057yiGUYDKsXW
HlDWOdYgxeljlmvgRnQMhyAX+sX9R7e34JJKwfHEIoXpDY70f6IpXym/LOB2pyvW9Do7kwP3R4pm
xxQg30mibJnOaV0PjxbauKO0PCCuYHec7WP/ehQCau/UjNcgCRa3TLsFqgnlNdRVcM/+citut5cL
lfd3C2qJZ3pTCEi8rrNaFnp1gz+JsoAR9cCtauHEFYEEjGVDN5DkNVrz0XXGy+WYFRFp7Qd6nrae
ZCoT4uMPlYvUICDrrxJ/SsDB3WYm0Q8aUr4i98/v+PNeRNzth7nomQ9ZGNnrkGE5Vx8QjZ4hdqRM
jFl0aWmZO4/wtc5URa9ZqdNyHOfjJOlgPvoMbloaZ27M3TOKw7b5Z/cc5yoLElAA+etPPoHILxqV
Vl05/rgX17RozZe3AvVY7losdN11TcLzbbW2IdEjMNeB+1htmgFUH/jnuq/kZ7KO4LZIgra9nKBb
R1QZLTglgfLxaQm20EHRldWoGdcbSSuAPaUnZcmlC8rjPSVXA32s7FliQrUcbo/8DMTWL7dY289d
c3XnoNGgq7OjeASGj3zdbXsdVXCceMJipajbz7VzNm6yBk5RZUnxbMXutfJuL8mscvMHu1b1LgFk
npRCMd4YYgpBd1kXRtKr8zltoybwJokWEZUnDopUZAfw7Lc4es5dnXt671UFBlhtbog/YBMZahys
fMvqcDuL+J1mAMkT9e62AGBQYDFQ/Je/DmhxNGfskij2sjiftabC6qGTQKMUC66TE/rC+b6UfSWm
1kpdkgyGo84/ypiajCcvxJvcFvST4fGZR1ZU0NswJ/4508aV3wYFGcNTjyzIuC7EB76MGSduYcoS
slrfCyJVocXrDSp9HOGOerb55cuN6DQiTtUihslFRMj5896mxHWh2rrgnJkVnSNrvb7fOT2qmZE+
OWGX2YA0P65zRwEer9lzQYKkjDMO1F4BlRfSprqeYYWJEFYGBiu0jw2tL/S9aLOIs8xUJqfBV6E6
lJpBudFFpY+41MdR65u1F81+pi4bGdLMHD7JdpxHLiZyT2HWczyXOtF6cdt4Bu2RZyzFF4sU2Rc/
T4RLtxTE0YYLMXyY28syXtCs1RBgi5BTYEQ56+cKFkefNiYL9J1787J4MnOuYTn4Kjik86eAkT4X
BGNVBQamt2uC/BzZfUdZG0olTrEaJ0zAp+NpJJ8i0+QZRQZjWVmNho5CIgDHBnt9SQBVItndLuIh
MrkcQPRuWeZatOZ0YdIgzQlrb9vGY7kvVDdsWCFmA+WrbuvsxSP3aGyIOCGQy9Buug+Sa9MqIfBp
AJNnurimxJVwbIurl0BHoZ57+3bLYwBLdiMZ1eSaEaauaNhc9gDZFjK5zN+dxCfabq5usD9CmDD6
PTNnihIpl1tmZccJ1pFijzOsv2D/lUz6dgW3GMAHtk9CB+1BF/O1rLQgHFLlZ3A8cfcZvxFsjnKE
qNKSYp5HNfwDXFA5EDyiEQlhu/vIcozomLgFORaUmGILasq+8L/QG13Ezd1B9Iui5EaYcgpgEZLh
AeyoWYa+H1ACMam6oSHSEblPRWVSDw0gkt7OVZmolmnXk9Ue6YqOxvX3eQWl+wZP9f/FYhozWHMk
QJRxrtxviHWbXFUOoYxxrNPCXgWNt/tm9mI4+VjJ7o5cj6EssOooYEnvX5WAt0d6cem2K9KGtj6u
t/UApFt7+V3/aRyEjQtf0e+8ErXFMBT5snJ1DYWlyhSn+zXNpXjVBzUVKSiwxhQ+eRg+UnefYbvK
NBJVGg+v2ySSY5WP6hnL8qfd3Tkp11OD8UNRG2V9gPTYJZdDzn03YN5liNWvNbJvI6ZfgrfjCL58
fgeRTyfvRIyR/A5wWBinUxbQLWhRzU/hr05WeKrPgj7pkDR8oMlA7Fb34B37CeWLY+Z/Yz+qBT59
HomN4IIeUO5Xd+COmlVE1FRn1dFEhfGA2G+jwFfgmW1OI0ilBkZnQTdAdvqpyVL+R+O1u8Ty+lJV
n5nfnuDVCb7maDhyR9oTxB8511e6LlGOYGQ+fYoK8R2C1FAHJcRgNt+pRlHIhEo5e2nLIsslF/cJ
16JLzdYC9CcF1HV7bmGKYO0lWyX6BHKs8stmsjibq1sXWvovVmz17uxilZC1aBsIGRrXRzPibstX
94FmzbzfiBMYvsv97LakvwvSu5jw9JFW1MP/8/jr9PnuvCubhswf4uPKLlBgLrlOavA/NpQOtVHE
ZnyCF66yZxS9PnJbt7nUXGNWSi8BTJZ9X/ftb35qS2lVvoqwQAB4dwLDUhKBPX8q5LMaKNRwLP4+
y6JvJzo/M8QGCUwUn7hvBW0b0Q1CGa+08oKAujlwVGMHaYesf15coq4+1iz948TnPjRKt39Ar5iG
hUoIssOVcTjT114aQ/DZjBFplCp5pLPa/nbts2pnvtjLwahkfFKCxdT53iWjh/kAjjCtKw8J84bx
KvRnWDKGD9yI2WumZyc0MjBQpE0o6H0OBPJCupgiY+rXKhuzrzc8j4LL1voAqrvbWYg62ZVPHklP
GPUUuUcjxdse66GzFTlZwny+8MfpADDy5qpssKpnbkVlyRz5loFSrf6GcReCNgHgILwrGCn1/tCF
4WydITs1iX91m4573i3HT/vGzoMQs2Cp2R130ZoluDH33ZemfSSHjkk2avEDp5WBHh4zbMVT/FGq
Q5MIR8WcPPEu73KdR5QxnGmdE4+3oXfZzo0KyLfgvmLluRJjyre7WfylC65qbd3xUcRq1MPiOYH2
8PIftspmJuPuJw4nUJRb7/mDR/eWq3he1fIQZ1xFrkVkVxfdh3agIiyGJ49PC1m9DbgeL+c8lOLk
QcUsWKKzWWnbEKhQIPR48bv2kY/hQk4XYmjG01H73+sqUXEARGfIKxjterq0mkARbkel2qihK074
453GuES8PZ7N2VvIBcNQmC28j9DuaGn/dVnQReiv12C5Hrhukr306TyorVIaYiiy7UqK5q6eEROe
p8e8TeDvkiE/hVMwdatB6cYogwbbr1w21PjR0WZlYq4C1695SYorBcOeb1x+P27OhqTQXFxr/xwB
tM6Db0XXF/+lhYxx8dXxVZumjFQQBoctRyQRsmUY3hP10W5CknQ5qtM3jTl3c4u58XUhNOs+gnHM
sJgQ+foZR+bPh39aVGbCsJ0cxfqkO9b5RL4wDAM7btBjXtmMF+P1YcJipqJ46xPGBWesBaOAHCX+
XRsxHRhwyKVD+BZeDI+7TX9KiRp2LU+cza4a1ArmrcYiKP60yq0fq7bnXadqVb7DrUkX5YrTz43E
1cZW3lmf6sT0/yTmrCacW/U+VLlj8IBzcvZVf7q9Wff8jzFo0IFnsnJC2kXo4g1hVMfvH4i9fWoM
lTBX4lLqRTBVpI/nco1PN18Nrkv3y3LAxliQhKAHtohZPYULStb+T7MuqoLQZzJe14yfkveMUQfb
be98S0k18yTiszIYN/YBAQRQ+64PYr3ngErlfbUfgV+jdBgfIW6Uws509Ha/iJ2FXQQXwjCm0IgV
s1Uwpe1EkYBCjSSd23YqVeXMTL5lUKDSy0CoMTJBJvUqEYcBSaq2vmJB94M1280R5NaMvgTYIKF2
JkT98TYUvi4WM+nPN/rAZ3fWdjU7k4oeNoSXXaoxVngwRw/f5oYn7X8O0miZbcl3d++Ik8g42SPJ
wo02gp3gqK6nv420IJ9QhbBNF6PAmebR9+k2e5dxpmcuNAAE5el7uk/3/mVRsGsJRU24m7B3RWHd
lkI8AuHfJRF1LtITQ4BVDMlddmlFLgC1PhWF+pwzs1xwnDiUuQ6x7i7VdVsDc3RSkwfLZdvJFBRp
vwgLwjAZ1tfUVHf63vjVg7MljY6KjETwRNcCBrJjvPAepmEVzTO7sOjjgYwp6uUuVSH0MpmrcujA
taWMP7FOhqquYTjHr+pe/t4D05TbZ6+9/qSgbZ71YYrxQD49KKJ6i46re0nsaI4aKHyzKcaSCySz
HIXLSnjqoJLIIxp0CyfeCz0Al4ZQff1OTeklSFSJeF4+dngCIrdb0ZND487InQ6S8bdjrWFEeTBM
1CwHOV56EwwcvHaRlk4qj55OO640oLBDFfmXzYK0AWSlUFwPlgGPuI6QLzW3ktNmmStoAaTGqfcO
5q20wdewQxiO4unbgqll7MO3lUaEl3qsJlCdJLLmCrmh3/n8VVMFcoY84byWa8Gz60XxSqZa6k3r
ATuGRgZxBpVTKeL06Tu1lGXFaVGZJA2e8hjW+bLZ/04teP/YniJ49dJdanHs+h5Rj3Xtr74cwR0W
c/STEtu8KVWkl/LQtLRfCEdfYDBMudoUsWGmGPEO/y0Sk78F359+y1c5uMrtpC52uQaaNfD7M7sL
Wsg1JDaPwMI4X2LhwJvVaev7QGA6muhWR50us4Hq31J4tO8jrbrFjkxFkGPsolX6r98s60fHPJEO
fJ55tPkQ4dlGi1Td5UiqB/LAHV+s7+8xOc4S102HC+s+wOYR/BjuRn8rAULb9jcaWktSq90NmiU1
ppU/UZ/o3/FNUikgTaX5kRkEwuw0WAai546PPSQDPQJLwoYFwmbtYwOjH8bYL9JMeWjyGNZ40m0+
P5UJ5WXEqL4kWKKClicVXDnmYEofFRpto0kneW+vOTTSNmYNxTk+Zw/09w1SFpcTGeGemliCeqrY
XZm0tZg1B0c3BUeUDj7GFl/9liNy319UnoavWwooyOqJHaRGAK71PqYrQQH7xTbekDsfRJr1sd3e
thecBu6LoOBZoc8cW7Lr+r+ivbol/6NWWMmnWskJHsKmGeNIGHuSXpZuNWITT3va2v1q/qszUMFv
oHytLTxslF7sCtWGVa3P5LDQlJUCodKP+irfLW99dsX5iVTop+Nxf4YOp8FEQzjTjXe2mRwzbirN
Mje0Anm+J0OQuwyFmD+pIGYvoFApAbGsd0Ofx8/KK8bKseq1RJ6mIrizHMw9KgXk7TLgyaWdbrnv
PwvjxcHH1gwqvCGGqlLmWfeeGRADv3QOy737YdhlphkDBAT46Xg1kMzH6aKJuI8OuEy52R796saI
1idEiiex+jaxPun8sCZ9jAdRbyst8s+TVCIRxh+hqhR9yBI6XIFtaCYGQL0tkKDoq89RPJHruJIa
RV/obzXEgSO8oRwCVS5befv7ygHq4Pv+KuZ1mtqG5F4cxy3cjA4Qb2LQgAHKx07E0oNmnUTa5rhZ
bHo7C8FkqrcycmhLpUA9hZRhjBhGpEkz6jiNQVEOVA1nmTD5bVVEmmz7kH0zXPbN0lsqEQPvfjqx
YgjV04WOMZsOxjFU97Ncd+zOuAKAGRR/U/ZAuk2PzwJWSZIqJFwDe2YJXNHfZPU6b22Q1mZ+tWoG
1u2VSkezZzagNGOV1L+VXl8v0Y0kag+DUS2etybjsnkr9invvrUmCcuAUBFDeQT32KHcaVj3RJgV
hRxWTg33Q9m8bHpjgiZ1THfrNdD3LVDhXkMrK/M8KYTJWryCCeFLWQq4TuCHbgzHb2h4q/XhdjSF
2JwxTSQs9DoS9LxIKR5cFJoVUmVUqnT28aBVFLjOGAI1LYXKz9kFTkhW9Otbu8M3zsWjz3WO5YEs
ohI0BRSd2jpHGMfGYs+QxlIcV46m1sVaJOtYmbtKAJ09ekNLOPTKOEppJBRGeLf9oMtjzGgKk+9o
OBwupXCqI3mDPMAfXiMuB84OVEMEkryjk2o6LhPkW9fd8ytLa4pTQl9AM4nHSi/nT/A/5IEDzvbu
/LCohhKFUVgM7G9oGSw9ejFZHSTw4+ytwAM70oInNSlFzKOxrTbcQsfqOJWehtFYqPITari+kZVP
goSYxA69q1pvGINo43IKZ0BR3YT04mtw69vw3X0gn3PLdqsRv7LQ+iM7l1zqtgzXhlfnt4liMpyG
4xf/ee8i40GgyIbjeaHGZpuOg+ky4P03TQt+oLyNZMxBfTcQ/gJbRMRF+d7xM+meGtoPVrVCjmRt
E05+MNVIoYNBjbYRxnBIFd6C27t2VbAwFt+0LF+9v7YTVQ9VSRgnxXLaO6F2hLQ9MsVDsc/7qIOl
xL7dSqIA03mIAaA/mMlMVCABjC0627ZzS6ecAYO4n2lzDHw1TibzpxqVSb/EDDkHChEleFJsItav
NzP2LG4kmIl8Cehy9fbNTCtXz+pjoSFUeqkbNA+LfBgtltrdy8r7jm+U7P5HLff5e5hbzEuqvK30
p0GtUVZaATSrgPDGEj64fLvFJ/2oja/Y2of4PNFDwIxVdsi+0J/+V8jPEeKBU+4pVdwCFtocxXdK
NCVXBuVqzNogshWHzqHaxtwClMSKooMaNp5k0aRWZpxNX4UNL/k+ckruSiIwBIDe3h9m43nzhf6S
Y738mWy3SyB7UK24DSR0l8EN4w7SIU5DBunTPOkVhT8xPqaTaHTrmzvRkdYalp2sFVxd4i7fKaAG
SPoUIAz72w8K0mjZ5mNWzOTwLLZo6b9a1kvSMA2pUkOD4bsQHUA/mNcF+iySEzo6uurjjeyQsYGE
//9qqHteeVYnll5KZMkS5jq9r8OdDLoe4i4LAmx+Ai7kAPGc4H+hlKhrOHXkDcUkDBN7uXrTlavp
LAZFnF/wBB4mm9vMObVLvyg4Bs6+deKWBe+4Ud+NyosxO9sA7FeS06zBVHd3YGjC58kJJTXbcAWV
Bojm/yTJLUI++ndCu9riL8tI9RC59rJhO14wgKbPXb0iQEVy3zVarSnlj/Ev7xd9IKjZZGSV5PcB
UVzlhWw61r/3sjpBftCbJg3Joj9EBIxWqBhEHWIRMrCIGzXh7wFSxp2jSirNgMIwHyOZG6fHDNWK
DS6llPTLkFLyYx4u/tlB7i7954/DqQ6Qjt0W6QshGBihoYY1lWXkQ8vj7dGa3qAuWp6xTcTootcn
TFbYSI7wsZqJN8D+C7v1bQELfM5Ct2tNPSclPZlh3Q8eVI07U+cilCZ5iUxa/TJLsGOYQEoeYY9G
MqNSPYS9ObtpsEK8jw2gQ9z8sZRUQf+ThMCoBpmFw0Y2Ac8wpt/lLk4NDIeONzgOApGDhq5B+Efz
M9GyxlujXVKCb9XUnsaAYkNDDUHQFbaXs5tb9z2ENFEiecJGOSwjWSNi/4oTgoe024EFNKsAfooV
oZnXXobtY68GV15NFnXTGoJUxxlU3ARvPZ+Nbv223ZQvetXD5US6Ej46D6VN3wru445q/W8mR63a
ve7yxK2xkrI4QFwX/BFo8qIHCAjyeQrBX+jUMnaJFS95BN4hixj7ZO4ilF9+nBmS8fZHPnQtFNtV
IP/QFiqYmf+dchl48qZ6FIbplPTCdsZkefYK5PofmZ77pUqbMIgxHahywC7W57kZf06p+6C9AVm5
C8JAuW1+c1VBIKEFLZDNXDExjdqHoh+pJr+j3nPSernprCEKl0PTgizEeRnJoWVeXl7JXTZk+zU5
0nKk9djlSCQ/l5M7dgflGybXJMiK1OLk+YKdt8eEVaV3UuDFgg3i3OEIv7OJCddo+wBxbKhkhD4G
BK3SWlme1b6emz8w4o0B4E+hbZaGAuw1ebi7g9H+lFhZNINRs8+0cqRknCNL7R21NObOy9u1Xku8
cx9OTDC5yygrQ9Cmwujzlkq739ro6PmjWlV2uNAyqUMHV93wm2+Uqsg6+LYhT+bL4S3jDsfqsJwJ
syLYPGVGQZiu8cMxSiCNE4k2zCrTZlAKUcVqh+UQTYTxOc+vZ6HrRKNWb/cEtdStEZ0gZ8w3Gthg
krIpa1szIYV871RFM01N5Sri3lI/d7w3icKzjoTXcNzZNa8JDUNqoyNjtTFTii0yYbPOJ6dZpehD
5ZpmHufrVJkGyZ5udv2y8/TAF/u+UTtTZZnAwD+mNlHR9SL9JOgf0h7VYIsNdLBW4MQvTugbIWOf
4BrppLW4K5A9TAVB1W06Q5igVV0TV1eLgSifGU2YTREmjaZUPAGyOALdJd0Rp5NPhPQns6d764fT
09TqwgnVnbsaAAitWVP4Hqsm3QreCE2sT0yz++5Ertvuqpz4oEPEOJLvKzTzjT5j5Df59RHlZasv
7QcwrnElLtT/tMl5qAt6nVs2Ilztoebxw0eLVlDK+NKaj83gBzDoCZ6nfQO17TNPg4pLNR1By3EI
sKvAA+X7cEy1vcGwpKOW+27q/4Q+ZF0bTJHerX6DeKixvz+emvw/+ed+0Rm8yMyKI5WiFoTsE8G6
tTEzdL324ioe1PsYMYF5v7SfD8JRUUtuGpIh7r+BUwq27Cv8Oqj8uVIMba93iVhR6E07nHuuSBDf
sTBiBViuh1gvQL3kOoKPApwFsrKoSn7IzvOlKmPdVTVifqmbBtPjUgxDimASPpuL3Fl5ZwwwiLnA
Vd9aMp0WE3un+c7uXzOr7mwLL9Wv5BOcgQfhbk0N/jO4I45T0At+BsHyzpOxoVIZ5jmWIBTkZnIW
HeFcUpMnrFNXQuenTenJUNDd/zDLWFdmTKMLk34AHDiYLth59X+hyoZ4Ykocyb/488guEsop6ecJ
NIK9DcIrpKkWO+T4E28MXmWdQt23FLbDCc/FPb8zTVU+HTiwgqO3ovZiGDjj2S0lcUIpSnrgaLJA
8l/qc/VwHUd0i7FMf1Owyv7WFGUhgVD+JDZm1d9+poSlkjPLIJ9bH6SLJLJO0HCRvdgf3bMh5Xw/
5hKkQTsUFrG9RsVTH3d6qG04BDtCSaJtZxxqnGHEIkNo/pQONt/yGSunuYrs5Sj2/8hvL7SPRhLT
pomUJ/wVf0rfhU9TTHy6/BO+L6vTPl6rvLv/20LQrhh7l7bwvY/VMCt7cQB0LgAbtDnQCbsz+fEg
hjxQp5eeAszCW1RBcsnejgcB9ou+f5a3k+diysiHEzgc1lxwLM3beUJhV4AATVIlzi6kMHTIIuAn
gx42TxrahAuu/N9tsPFOTXHvT7rG3boy8zbMR1BbqiT5ppWNXzDpe4ch2HmYQF0r+ayRVQvFWXLh
hbDt3kIcAm588HKQxhlm6NCsAi+4m/IE8BZsRRqlAjn9pa9mo9v+nMaB73nmNxhEbruTdT0Ojxh7
fC3gYnqRlsitO5S81g8D4fBH2u3HN2dxUHwfo586GriAiQx5hTyfdyuxqbAfjp8cy5H7OMHOJqeD
zyn6s6B5Q+yq6AULeILlZWpb7H+qY6adfRdWzC4Jto1CUVOO4uR9QgRKNTbiCBHtrBt0kZ8fvO1n
K+lzlbyLuvh/pw0/xbr+HLeu8UBKHDbAW58D2Nw0uaw1ZCZ5O4CBw4TmqRGFXUgxvIEEnp2ZZDqA
DqScqTRb/tvSp0XbXVt7CIc1rC3kTWRo1Uvp3XTAgY/l6l0u/O6U8ueqQQD1Jalw5ca3eQfR8VjN
wTzSTSuuSTiWhrdAkqLTiVbXne/Gko0q6MPgiMG4FE3wtTLe69B+no3h7Z3uTWAEC+M9FW5DQDf7
fclx9oYtR6WRxC2S1fT1LVSLWx1Q75xaAGFWuoQ+lbgaMfcPA1/8H3TMIZlPU/VBKqqFNFa3Fu9V
fGWrcdmFoDgTnQL0BNtclZrbhFgmZhsyBLQvN7/G/MpoA0v1BqfnZrCcqa5CBZpz845mX1zjO0c4
z8IJvxpSLaTPAV92vRAZVEg+cnJAxkrIKwwaGFYS0QTf80grgobSe0mKiu95p9qAyHmM+eaohy92
sKs49OaQHtIGKDBX3AxKh/dG7CqecK9e1fSF5wuHrhJh0Hno3cEqAZ6tLG0ZC/2C2pHeDpjwqNm1
NJW94DRbMaIbn/cAmB5LLBUjoeQTq4g37sdF+PZXYzYt8dLICpN9ghp8WGSF6yn8WGvtPCvZyfbP
iOlNmM/S4Q8TmQc7YlafyR+GnHjSSBULmsn6FaOa4xyE1mja+v/fBSPwb93Y0H/+Oxbvrhgofuxg
gGhIIFIeNtTo80btF3u7lPIRfExym162zBEYXqTlGPMZIqfAwIEprXxW3El9DL3JLlgGX2xEUJAy
86n4efUYe3sHoUcV3LrMV3HXQqASs7bD682BLJd7BNZDAORV1VaQhQj8zNwsF0anyHkQicZHrDVH
ablGAC5IiH8KQEMHj4EvhAZJuAKOUvdMKI/6Pd3+KgmslIvLhLgBkVm5pXoQKpHQIliUYhHcmQ/P
U1vN9SyuBaO1eJJQ3xjv1IMhJ3Xp7cU9gf6PmjXtpvCKT/2/mWsUigZbiC6f4f7KOMLTvDaUM1Ps
g56jHOTP9d47FlBkWXHpyPGobtMQ+ie3VNoSpXkJxvMW+7VoVXi2JFzPOaHqOljnPh/cJJZ0m8QC
bTYJx2wpCnxsiWSf7vfhWsVOIPIbP6qefjebnaJITAZT1hetZqZBkjg+84zg6Pwqa7ddf4VD5wbO
5WLlthJLqHp5R5lOAdtSH1Qwb1sjGiMZPDsBo/hByfcm3LkPwPToZj9/PHGyTUQzeEEOzMnq6uvq
tNYCmdzqEWvxcBo6dZ7qUEU34pY+3grEMVSLMHSOj1NelP+wB7Vuy2QbtbQ6ZJbzT5Wmdw5XBzkk
TOxSVLLPfH9VkwUZJx733fnhWZbq0vXOcY8u7rbTShoBt7m8+zZtrbEomWyL0ig+E6ZwZDCJdwW6
A07jbysdD0eO3Iwhq6Rq8Ouxt18rWmac+XN0SGVj5H6Pea1CWVKVyuFxObGrOo+mIHRwwVKiC0LD
PumBqHtGmOlUbH0saZOwqDojMjfaIkugmbmxeVL0B8aCweiEQwCYTsz2+M0O8wilBkgViQunhwgz
EQMpbCg++lDTjdPQJDGACYUG8jGoEyZwVX6tOmLo8dnU7LHZ7Y74TZjnhooiHC4sFqp2sW+vTTg1
OMGtIqAD63dDR0uYZBI+Ouzhn48FFdH4miDZvCczsAY1SXuynfBRmMAkaUFko5a4Wl7Pf7+C98VJ
dMm4eMVgJeZXoNH1hQbOE84KK7S9Jbb7v8z2ZegwibWAlbcMh2zTA2R2ZjI7D+h2vcw8YJeg9cqm
qbahFl1mgy5b74esddEsMTmlxPJi66tcBOOmLNy4YGldp1v7AkpZuobT8bQPGvwLD/PEeDWgoz7o
9+bzUGnC+lXSNrZHhVMiEEoDUkCVqSEa69rlSdlP4Zks29C4VKj+luQSbXoXGKAkcWZfDtJY6eK7
HYqczmgQP+deT/a9wiY8pMgohOfnBN0B6SLjldJ4CYG7dRvfqnUe2Ck0wX45pIp4kpq4XH9TLW/4
s8SsmnDe1UoARjaBeC6TEsadWTfQT/H9LKQSsHxbpQvydUhKm00HR+wP1TLzJOLl9gMTLRH3RHd2
3QaBNr4dcpCBSFwHckwYDyDdT88aQ64k+2hSvyhgN17xfOIv1WcpiivMKAaY5mk2VoKL1w4gASlW
Rw71zvykm906RQ+bF+yMCJWFfeVv19HkI73MPpIZ9HFny9ZLtPUNBizsTq3jK4ImNIK2ozLVqNFq
RpVzfV7Qw7loZn4C408JJ7fveWQav4+z2wKPBNY1NTlWUZyPpj42br8/mP47IYlliToqBa6AXUC9
Gzwn3F2zf6tdeM/c9beUMkfZGBTQVztVvNe4Jj0A+3kZnl2eVPy4gzK9wvDFLsch02sq+FVob50A
MmSKbuopyN6CeBuUsTxcGEfKnZa5bOgm9C5SecHyUVlhKWxCzYB7aiQLBrfcV687nZt3sSh8aJob
B/ShAon4I+AoWGPjkIBOs4KVFoK2Yjs+i3UVkDl66EZ7filJ3JnQqEjWLd8LN3RplSL9s73KmQpA
C/I0uMomnGFbtetnPCs7pBM79f0sJQKUb7Z70ZiOl7BpliLcoX4WRbmAOr0ANosNCyFUdkJc01Sc
Tgpy+Qlnrra2+y9SlwF6m6nbGV/pj32pQRFJiZvjiZ+l3ojPmtVMJTSdcypdZ2o6CX/se6ARE74Z
xxqIyzIB8Smpoa37zjEj9dRvKoPVdeRp+jsX7Nb4hM5MevVaaX/icK7ew9WTQcH8b5dQI4XFvQ05
TksF8NLPdjHFJUGuVvRhBkuTk/8ENf4rULxyZQiyOoS5oksvxu76z4RS4YNQy35xXzis32G+HbqF
UuCsMiUCdSgS79NpofPwqQldq5zE1AWWPaIT5X1q0q2Minga8qbLBHaxea+rRj++PnNvlv7rT22v
Xa+fw9b68G5bt+JuziWquusbE0k5OlZiF7N0QBCp/7VK8X9xEqhe7gAZnU8qU4ADA1F7xrMSOLFX
AgKr3UtRq6898pWg88GObWtkV0Vd+ByNrW1lL/5t9bJCaLPNEgb91+5SKbYwP+ot5LlZkzV7ZDRQ
+vapSV6oq6BsTjC9ZE4QRb78gFV+fGqgdCAh3tFgoVrRXihbFRPTsg/f0KHquU9W85LyfpgdSKf5
hkp/TaECcb+yISuvJpJlabhbbOcQLQ39OCm/kR5zkDmfSwFLRrofVOWQ4SpL/IHcbmBUVNOOohFw
hsfGDr7SEeNyr4ksKAXQ0JbuiJPrbJH2CrehP2db6sev/mM5TFjER2UvXozAu8tmKL6EetHltN2b
X/r+C0kCsIzmAJ6MKrup8pC/kQO+cZAnVzFAz81gNMIxi0ve+X/AwS/52KqUkJ9c5npr5lbKshz4
wdYLTGsEr4XfXMIZtnaVlxN/Mw0BI3643sWhxQo/ZoMWdcEysdUSKK7F+Znm7voQxIC+vcl1vc1V
w4MZMpmDQBMDuo6FSPJxeoLjgviTGbO2DDizJcDgs1vY6JUX4kGqXAgKLvBSUs6aXZcZ+pt57WvY
smirMECbwsJ7ubvZUI8bZFPhM7xj1trGaPQ07aEeTdJEe+ysxrKGdrqg1XojnkAOuc9vI0Mbi4GV
qg0q/CanDbJU9mMw0RbI4WdSlKIGI6evr4bUa1Lv4DoUp3qyQn/GHD4TTaKd7d7Uiyy8ZigsdMyO
GpoZpxpG9RHUlGlDMlQkUaBhC/L6L7DPH9vSwAZK+etPSUEkS2IyB8gIz/VSvWXFnb5JZOuXUuHb
0lyqvIdS0f1q9kt12mYHxQ387k3Db0X4BIUoThw2ATluS+7JTrjeYkeFO8lH4+jM8IvE462dQwDo
z+B6Y6psCRoFj5M1CskLqf5/fYrMiY7+snsGJ5l73pkUl0bgomwj4kV2Aq1R0IfemHQksdL4jz9I
/Mm1lgrIryuSC2hVim1JlF4u+JHLblR5+PU11Loqt/MJcyKxlVYspkVKkcw1ExPIjRZnwPegN4KM
w2NsRMYuvERRS64ziuJ7g6vzkiKXLOMT1dPYA1weSrj4QszzUyTBX8BhN11RFpfHbMyz1JPFjBzj
mKnbQUT610jg8QguRsniY7QNG/X5SbKLS9T2+LcV+LRlQDrDAlR/+mxQaNCnTOpXjNccfvSRX7n8
VKEH8OmLLj62VM/KuNJq2Pg2+5ZpYtiSFYTat4zAi+JXfHHVxYfJvAxSr4OcrK9dmrOBIWg2pYXB
M4HeWm3nBx9ztcDIm9Be7ps137eYjtICHn571rlb0eolQ5H7X2ex3XL1lgaGDD8rzp/q9eh4Afak
q57R5wBxmGuOB8EOdlOmg4O00CFFQas3Ggd2xcS3TzPpA5WT2EzT+PJbHudznggN9xa9Laahk2b4
/Ch8dwexHagN8jIKCf2T79AHTBY82FHpxEeTS4ht0i8WDgyKpNdkFStEAUXNGJDg/HTfUzBj58x6
lDF803dQtTZZxBRY3AChvCvZGBrmf6jmy4nr9Cl2qK/+amqyKrHBd/4f8C5jc51LvlfdPS2T/IE6
R+UDEp9VgPVNo+rM9y7eKJdZJqekp7Hifn5fPweW62CHAbwmml7n0Vys4zbzZytz2fF3Jh3nYBLt
zMmzDZlzl+6R9MHsqUXaa5wkrBlxDCqLqEJ0m1e1wU7uiBP1+uJYJvQEcFmmu247xP7PVqYrTmX+
GCTa+5RP/J0+JjsY+GTmrbS6S2r6rR+DL8ljSVt8OKz9TW57feiRg0Bi9l6QpiEhmHTZPhZTE4tW
3nrebhQkr/QK8b2x8iOB/1R4NMb9O7+tUtzrfy6qOiLmf4bSi/62WTmaf+xbOnfIqbd1XkBXARnb
YE2BXaRN4j74+WzKTmnNqyZTYZS/Mpilgyv5F+C5V5OzdO8E8zXy4T5O20tTJcObslioqiJdolYi
MobcuHOqEfEvbP7AcybxPWGCydhC0syhgDiEXtjNDkOzJddVpfpysMukXRgz1WbekRInMNFu6GIQ
mEnHGdMlzHO4aNN8Vuz3eEa0JegDI7u+stiF0T1LNPIDZSSnXPK/aelcepdMRYfFMm1dcuWMTp5h
tLHglQ+PdQtr1uFQygHKNBhwbOMlLwT8y9CqoNN8D0oenqXnm3D0DkQ69FcYU5mtpPLPAMqijrMi
2RQC5iRSAScjph3GXKkpMUPne6O9m22c1M4YNxIB4wu6NEXCR96FTmjcb6SLzOq1lGOIk3Q6aiR4
BIjqtiHwocrAZX15dMO1TdlJKEoDwS/Yr0el/W/DZ8jOH3BhcO9kQ+rNZXSdfrmqT5ctvaHuVARd
i4hCPNcMzKaVIR1bZ7jZgBrqxE8AwTLxDNoVQ6GC9G0mHZW0iq843FS8M3YpTn0/vRFgKrKjr/L8
C3ktfIrQdCdK8Gd8ayYrceocl4mKk/0mreHd8zehuwWXpe+kTcFswSbCe1I3WzRfjarv8QYA4q0l
fmVRdYYZ+Tvq1dc3e3Vw2LlOJz1JEyVqIiQiBfdLyugG6DlJa5NKe2ilHInhWFy/q4NmPuTwU0aI
rbtYxL/15CFT25Hu0M4Y4ebqD8AQhtraqXvbUThWoQyQRnbCIoQ9m3RtYWqmTH1+RYSh1cb1pv8n
oJjUJ7inuMw95S/YZBvfw3wydnasIGijBWXzSoNzRtJbDolXJcP3krMu4yj9EzRepF6WDAB57kZa
zlr3jLypWScVxGrOuUBkzoKS6NEuxx3xIXY/WhVmPm2rFBFpunKO68Op09DgIHT2D905dK9prW7m
2ByURE+ZF/mq+6qyJVruWENBWCOuLpXP8Q5LjJVDdqTizdYEZwU/vMtym+kO8697LLOEv3udaeNe
M3f0htx66C7mymAfZOJyVgXlBJdegHT6uM54tVF7aJ1Wvm8YSUu3bUINQkRogm1w7DutxlfOOKfa
ZfVToUXJH99zu1JWSfjw1+tNiVoaXcSyxIvXztoM72e6dc4KfSZLBxD4wDArjCuBDzQZpq06OtE5
RwuuIinD6LKNk67LYbUj5JfF/WfMleWoD2sxusxx5qA+/2bQv6I0EDn3Fd7O1LSE5+tAawcxtlKi
FsOcIApO8jMsobQHv5B2gSH7nwM3RpW7P19F25McKGLakU07h99wvxavNgHa1rJGEGWqV5zUtFDx
SrJCqeJ8+aU7C01wrqOcmH92C+s3+XnEEOwY2FkjbOBUIit2HLP0Bf0xUAL3UupSE9zGRV3mCSLw
/UskHiOfSqPrY0Aq6LU0rYtUza4IY8QOrEyui6vo7nh+rpw7cuPhy9ccSAYsGOHQK9sg8oCm1XWq
VIX7Y0jvRHNqsACZ5a1I7kIAgrh3lTU5XzyxMX7Sze3+NZJnp0036GS/71XcE8wyCOdlYWXl0jsx
VCgYLKV2hFqQabZTrYOBSAv5FdM3hCdV+YFgPrrYMLFmTEMmMNReLenuE4F57DsfBaMsd6yUCSn6
3qK8rO3VM6XxpXqirtDwRWH8hzKnWrlU2/UkCUUiBUH5bSoCEL4y8CxW7UYjOQWCWuwDSg/VQwFu
IEsLr1/bPV05Vxws/ONHy0cjffsuQxvlH9bv3o4B/ooDXgWiYQ5icz5FE8oaMkhlt91vpQth3bRW
fimQaoYSyfP6/GXDul6eIuDENqwzY6arTRAm+AiCzs3bRKQEcZ3WmjIsYSScm7a+e7XQi4nVRI2y
+8PT/DF006VD/LsGekRNHcFKKlCjCYABidiYXt87/bctjRfn1qAwgsYRpNOKp6y+fKztKHl/i2fH
5NhZ+HQXr26mYTnyqKvczxe7NxRRL5tQdSiiByrP+23zZfoEjGBfJG5KnO7UpBS6FivtsfgU8omG
Q3Zw7Xtc6zQJohAUUZkArXuiKAkg2pTk8HW8MUDzIDiZeUUsBeRwfTRXpEJj+hgnItu8ryGQ8wm1
kBFr9T7HIxNSWLKCxwYDmTJpX0IPgaNdjvAbyuuVPRDoQPDknNCHsBE2gpi+tM0T7AIlYoZMyOpR
cF7nlvgqANDtZJkVkS6GY+BTu65xaWgB+Gr1s/Exfg9Om2WLKE/lIlEbq/rpHG1xqhgpU2N7co9y
/QeRbKyn5NfXDepWgRkZyyfF1KRhwnQWlx9Vtdxwzr6P+FwNOLCawIkCzPDbme7XN5QD0dF9S4PJ
fA6+3z2rua0sEXNNiPdfEO5SExFckUVlvsjF84IgZLRpMi2GFJU9AIMka90F586qg8UQuM7RHzh7
7ahocxBD4MiOm3+XoBrZnRKOX7oShP+NQl0H+BftT3Aia86ckcAYPIBX8b02sb+8pMV/2P6A6Rjt
qSLNHy6qVXkpiz6WwZPJjJG+Tu2SoIBqeYZTIkH9kV6LzdBTpO2XQxdzOp/mYwrqsEx2oFwIBWy7
iW7xjU8WyDHON94Y2tS4C4yaDms4fCQA8KOOby9x8ZgfjIPAOPCrJp0YwVhYBHG1Ai/03Xi/rcdD
KMeWJuXoWkICKYPo8Ia8nLrBzn/O+bngNBnUx7y77bFjsG/WdZpJALHljpM+KvsndGf8jj90m4/7
cVIPt49iQh63Vmum9KSZC/az7clqgHzVwE1dWrnXUlq+ppCaPI1qzy5Jvlh78YkD+hQ29Wk+fCCt
5DQcuW5UPYQfP545kk/fEq4hjRw2B9jZ4hnQFZTzkdpVWAMqEeWQbtUR8RykB9fupkEBIV/tHmtG
SXYoO0zvpKc0059R44FNTEcLSSpVSrN5e0loOYVZ0wAWkscbaOhc9fCfVrIqsdLFm7X9sGNmYwmJ
MWt1Re+qVQz/nPPMfCAB9ssBCnVSb3V8VEhG/nHysTmPY3wx8mSpIMQCszoUnOs9BrZiOmEajHcr
Qi2OR8P2y7xzENvrdOpVVTSGWSHppC2d+gHvupohHNEWfCO6ALf1oMr9beaYBnRkUVkSVZOBZCxx
j9ZbK0MaF+YoSF9FpRxOBUel8uzqoUlAAiMUoY4ye3fZrDxDZV8Uq8UbHiyc97G4dHtI9njTlqCS
S85lYGGx4YyzNei/s+7VEdA92y/LijXWLNV1iH7IzJitxDxsXEddp18i6tHzffFVXGnLcwK/xtfc
wkf1hXwG8bQ7NovlMehVsnfaDtionb30vu4ivvVO4QeBH8jhM3tJyGh3/g3LnASrX5w2svwLfll6
80iCyLiz2ODURd01HDdPbxoKp7yV+jpaPOnhhjfiRYBl7ebIVuFyimolp1VoEh6VfaqXCvDUD2Rt
FNcGm+wPlMxVwzanhgeH5IrH+EGFnjULjAZHxLDhRhV9P05lRYsuML9JCoPy/Uw+TED/gy2yp0TS
XMSY3Y3DHdEO2efablCgwbY5LopPtAq4U9mDi0USyEK06NBcii71Ies1t3ob1GFzagQe8QJpBAgF
0ONIpP9Zz/y6v4mZlp/ZgSxbl3+xjyqeth3NpmWEcQsir3j98uP1lOB8AbINtjitPZ2BGmK0bvHK
hgtnzkS2duz+vBF99zcNMGQPLnaf1kwxleWVJ9q3xuCaLVeWelV8Oq5opLnigbG8eYpbv7wSKcE+
VtzPHPYrbMUJRkIceq8taIGxsE31OG/7+CW6w1Hk6YJfEZrPHYD9INehAAIreA2pJXwIqJtoGb2m
IqgMeLrqAZJ5YjOx66EDoHGAS+29CbrCJaf8nrS43V/Utm1v8uA8jN2Z7VmabG7OfxppwibX4vjY
7b85jTWQE+v8nS87QhugQMIEylnlo2eM0Pq+hm/dSXf0QCECZtLth3hygjpsrB3RNTU3Hz+Oc9Cl
zbvN4iQkbKryAeczc1P11NG/ehNrEduotpoBiSh8VTnJgqi1BXTX1aqk42GDAwQ2M+2hkZ2Ljk/P
Q0lvfp1oTyhF9if9avY+xmuXCOfGvKT08TNZ36l7QktHMxuB+fcSVSgPmOL+aUEn8RNJzipzwCaT
j4gJnahA3XS6MihRHMg0jp8X04ReECmGPn9Ko+tlSHUzLVUReQspgQXW9JgbTR9McWzxff1YY/aV
5sZJ/pvK+QRTzx0LKtwQyHIcIGEv+yOB2N1uDMgwRnvSBxGwWrHIXM2KSTd6wTl71zTwtSHLYM2Q
KEqg456wSmKAun2Hex21uptHHWP0L5RL7bgkFq8dt73KLyv/q+rDNxfUDa5fbQsvGBuSLgQeT4iB
KjgExmlMxkrJJZdGn0Rr+OtAr2yT3eGyYv+PS9qGRC0nAqNoN5Qm0AfjLUxaRTt2cG0YcR2xC6SA
FVH/l3561edX2D6767ZDfwmDQ49odYp5Q0nvgMUgswlbL/CjP6518vg8HTxsCWFeGlwtosz5foxi
Fc+tgcVu9eW1X4erDO5aiRNiau8JexHa4mgisUh91n8thxyFxXMm2rbNrGts6915bykY8RcljS1R
w9kC3YGkqhGtYsVK+dx6Zq27g17fhh93031JhjKYDRyDToj00iSIEqOXsgqMU/Z78CWFb8wkdvm/
3ixZzlqOVl44n9EbhewdXYG0FO6tK8Ng7NrICZjeOThb+lkCJMHtHWfkvFn5h8GF/qlzlDIwmhFd
KXER0TuFwa7Ps+Iq2B0vDwZDugyzbjwac5FWFwI52uRGtClkx+Gd21QS3Oyjv9uOk5cYrF4ij7f8
I+M+bgKigpELwzCwvTkvyKxTEzySEac0gFwU72BjsMrcawYlQMMCAPlHRlWwS9Ba/R73UYBISV0N
Y/eIioQGqwmRb5aBrFqsv7romYdz4lQavjxhFR6ApjXDQ2lexc9m+RKMFRJYu0hZxmqu69gG9/PN
QYuqKh9ANp1LnddnXTmCG1qHuwlz/WEHpt2asZ4LB3OvrW2vXfTUdnBONUzVxXaysRqmVHj3t2lk
p5bdjV0OPyyEe516grV2aP/f5C/afzCEh7KywbZpbAclpDJooD9PgqePD+GhBteAnDzts8/Lo2U/
qBF3WAvWHXPQTX1DlH4d2L3K+jTqoH78ymdg0oinI7rQ7VpybN/fAJqSeCpx+CGNuCzuAX0Pu3Ik
xCovfeKbjVfzFWGPiNGiAq1SsTN7iQXnnn7pbZWd+MGHIJi8mDVBuiP5GiTHbYDLkig7EpBB5dh4
1R3h5Nq9NmRNZQRd+VNwzAqqoCYBXxs6NI4lJKpqnMZvcGdWNLY068z7WlviZ+llnQDjiccCBs3N
rq3wl1l/pAIax3DYvMbq6x8uf7BZrxgIbsv0QJRdnznDm8X8XAUBTJI2gS7bOSKa1pYm8CMyj51A
n4M3raavG/H5DK+RYzn5B6NQEHSYc4nCihOYlaLLUrABUJ7/D50MOywYE09FVqK6bT7kWooYiyKX
Tb0fi5xFhi6BB7lncBAUFTdM5Mu5Msi17dvv4lMKYJPWPqDvc1zE5Qk3lpWWmkqYR+k4o8ZbUDdx
g7+uGtGJQCc1Fuaa5h8lhw2Vlzt9NSLU166xvwUGYZ2kPZkAN/Tgnk8sJdcpKiV33XSNMn0jTM1M
nzUQPzRH5wIU97v1SAaaaYFf4ODpARkqiD8XBxfxERrYNpFi9oympYkGwWKKlRj9DVLSBTYK+PV9
LyLurM7M2yID4pkyumSg2XFREbrwEp+vPTt2NIIxG73k0Ye4zeq+khxG75obIo/QempbnJNy5hYb
F3UmH795AC1gZIWHGXdH8lowCLWJp+NLgJOrPU+7LTD1vG0OvC3rut/K2LBN0RUVUF27Cjzz7xqy
1ktAitQ4vcdxB0Hg+DpcZeRGXLGjWANE1U8L3e0ldZTkWyo6U2jOkbPxjz1xxst8l58QQJsrSggV
HRe9yYMH7cR1fdPM5MO3CimoB0iDbqLg+a3/Ab2nizlILLk4EQ19RMuXqCTj2eZVVZOmbtxgkfM9
ER8RNYNnsm0yA0kqI0iYgaFpSh5z/f9S1puiJOrHXYgT2qfFolWhiXQWuc1q4ahzywjyrCIbmp/m
XjyeD+dPv8WtdAhR2FFM1F/zrS4fUgt66tllAkESWJ1ftFVRUXtR/Pwt5EiX4P4+zOoFFtUM39gx
EPoI+4hzyOf5AdZkRlvW5q1d4KrMIlnzH+HKIwEP6cLXyt0wK1K4OaZZNeUcUROXcwMycC3XbL1r
QHyGlBP1WIdtnYsMLV//oHErvQzSaQbKIFPtSUiThW4th4uh3jqLA0G2nnemrVDE0dJ1YyiInBCr
X8rrwGyiDzvBq9AiR10ib1RfzxTOE7MO81d2WPozkwDpnO0FPKZ654dlU7L5P9Y6Z2D0GCm1hFbZ
FXalaLp/oTg6IPnH9A35zhmctdCaKv5eFaTzwdk8v0buV1+IgyH2EnCzrkK/mg5mjNgB2R+5h8cM
cmAovrCH5aNluL0nWS0lPMZLz8CYmKtQ9H5VBnp2KkDXzuGyIh0lg0LpAKhUk/awdBeUaF0W/H3Y
8JXUsT2PGkjGI3pBK8Z9EaQ/5ZSjLUWjuXhecTlkaBli2mQZFN8lG7jHZuR6eHnNbMX2RMt6Hljx
rFJj84ewIGEv1guUhpnKWK5hJry5rGE/jALQXFFZCMcTkoHVVBhFmMbxq47X6JdjVgEoqt3iNYnt
dWjCWgsebIcelUY/vmHMUQIjJ9msnhr5Cgw1jzaWDRc8A/Mypai5twLrzDdR8kOBB/jX97wulJT2
iWm7z+pmAEhBM2DBg6/Y9JuEmX7Wfe8CxczpYCPZ00cZQijmBE4yEXpV6YmDXuAJV269JSWkM2/y
NA6LWBd6Ycqr1SXDO2nRaqtX2DEizQYhe9uzXUlNx8bhhJ7aE64hFQ334GSXcaV+Hb+Tl/wv7iS9
vpH49AAQUPk782PAovaVsRUoq4qOeqL9UP/H9c1dG0sLC0KfrwPwc1BoOCPr8O4pLRIj2lP/L8eG
uus2WPHxA5XuLPwImpcDJ5X6/Ruzsso5wB1ePrlitjB5E9JjqKnJbse7M+aobUFmzwEa5/x81uLJ
mp/RRwtaVks1L3Gs3Pe9AapS6LJZUqJS7k0Xowf4N++bFDHeQkWyqcyvG7+OuWFzyVqui+JysQtU
ypHejzDyADTiUlhDlRQ0tUhIq+fqGViNBuVs7obj4T/+b3kWzBhdVEI7wTzIpDZcAupH/AyQ3jk2
bG5DsliFxVSl2v2og7l6r9QrCZx6nefqTZOcwIdEbCsCkFMTmyopsiZlE02DL3x0bGF0DuCoO8jY
TQBicIrtRnkX8Ap1HINKxF9EPe1qBw4eZWMLybGtcYuqsN5J/9op4DHLogBww+6pjvx7TBBKKt2G
FCpYugC9V6+eBpiVZ/UwyBBKaFox6AOnqfoAgUFXyIGfM9J/oadZlDLVlBBNN72nqnPMU8zqBH4v
0ugpK/EZPg2sgfwstf3VhTUNYNaR0YDriIUS6qzlX1tt81dejOBYxC4GeqCEs20F45AR5USD2wOn
RMA35cbgWc9HEf/0QdKHzm2L69dsIhTZ/RpYJgEVPHtBoJzlsD7RbAdtpnyQ91GiNr/erYMhvuLr
KYR5xiSpPylMHaJtZgpcP6p1kPpaS5Nl6bLJnvNtlza/02IaxEKKn2r5aqZPJTObS79W+F+Ljit7
iS1ZXo0otNEE4lijbIVFnxteBeKcfFu8FiMB/WNez0RQ7NRHXyzxEZ3ECCTpl4dcrqhet+BUnueG
cUBPe6TCeVaNTm8lE+QoL0JKmlVQanUgDu18PjMQDBpYi99T3NwaRMTKJkhZqs5EW63FxROWoeZ5
yq7Yh583OlbHOsVq6ZPqXHZb/POz4ky7jo94gIIPO18flxpq0fSn7/qQQNfkdfPw4eRrXxiLJpmn
DCTalgqzQ/JAU9MOEJKqjlA3SEuVadTz7MTTneYSPGqGmABoUwa4mjO3x9aRvO9APgoJmDwzjI7m
KwgfHLl8x2mdYcQ0RC3mbgqKZSh58n3i0LwT147QSULYpUrX+ZqOGclq7lpGomd/0T/fZbcGbv0T
rDZbaWKF+UXI1yhHnjroCEu0fcQs4X0a8yewfCnAoVvg0L0Vb5iUSspl3cK/qO1PPgjvozQtnI7l
i4ZkOuRKanBVdtPELlruBpAO6Wtng1FbhR6/aaBGV60zD8Lh2NLK1VfrYfsLw+k6dgQjktJCTHjG
ru79WVvnvZ17zNMjQjuFbS0Vh7s/Q7UR6bUlKhza1JSBufmkgEsBQpnPMxBrmcHvyu7l5P636PGo
Ykaa3hcsUPTXJE5bOm004lT8yjVN9XAqfnF9O6W68O6Pu/Tf7kAZDnA8Z+kgQ47sKxqZf83+m3JX
0YvpkZa0rQj28dLAc4LARXW1/BFKASak26mY1NppwXQd0jRn5ptfz8F2ga+vKn6KeJDay8dRBkXf
lkqjzptn80mH+aHoBjl2cXi5krWMVEiEPQI4XoYivEcC6YHGHkMrQ0UqSwv0oDRG4L45qWhLf060
I9TRS1rBYKSg6yhzXEr4ofljpjgvLl9vc2dkbE6Ok6apyfZApBMMyDI3HIb2TW9u3pbWNOQy55rq
BYCRf4Xz0mqcdFkDoDKenF5NRfGuWqkrtzFL9SbF8C9QMKaqbPBsxBDhaIjzkebAne1JUE+oQAVi
3yXww2K89h0cE+tc/j41VmQYRZYhgNbOn97EWjZ3E6kh0fyQXDH/6JzgA052G1W9Fyj9sP5/rYAd
fnrXGOSLORbp59SZVSGg/VzDtHh2aVKoQBglyAwmvr29Y0bAp5M7xVO+efHC3JPTY9ThbS5NC6Sc
sbcAEgj+AIy0XZzF+S14LxH4iLeFmpHVe4w1FhqhzPgOqmYdCwgKA2gQe2du5w1zM9UfgtbbSgw4
5g9Ap64VnfZBsUH4Zvgdu2/1dx0R5PMlObgLxDASFg7I9Y6kRJYSO/74pvbOMfoL9u3dI+Hc7QSH
E7kez0DjfuGkoI9/c33pWE2rFinBpTDQgTgVyUpW611X9Q/Ad8YpDJk2y0BACwEtQPfGaDi6/PdM
oZXXug9OWidEEhKKco8tDAmHdrYaZfRlYHxiVbHcz4hKZOae9XmaMXjz8dU0hWDUvoiPsyxuLCxb
h/PFfcy2MtGGYgyddwSKgMGX9AsSP13QDUslZVHEqE60kb9MoBSniNKtrKYHp35PTYu817m+doRo
90fyhvU/Ee4KnrpTHqDmP9OR7oJjppIMOwsmQNNXZcZCY4XH8Nn/0kVTRAgB9J3jAM2Wp7Y6tL7G
3wRFKraALmkWYVg+XhjowRO/X2D6UhEIymrZxsbK/uGUt28w29HxAmF/DpT1Q6tM+nMIzbY2Khkh
p+gmscxs7FE/m5zqhrEu3gK7FEPhPr+3EuIJpk4L930w5unmOMJiN/yd6+La31bQD1g2/7GbppFW
Sglznz4rEBud8LKOZzb0Mvn/E5nN9hYqMGu3qD+BP79m4IXjDhJE2hRRsUiC1QFWiuxBiacWFUCX
YiTaTgnm2sGts8WfCCoSpbKGGSjxRY7fLBPQXmLssqQm6DyLZwRUu+ShZqozgCAcZZBefwNwFSSm
QvkxTS5KXki5UcEm/WELyqFM6CD+WIQPVyoNl0+N8Nc+2ig081XOWsHTU16yocnR01UuqOe/MMb/
PMwJw46laIsQvfRt1Y14Dc3borf0stPx4ZRZ3GeYAxaHR/qoJ+Tkf41ROwpSRQw27fFNK4e3K1ZC
OO7+XkzmfHjY5mIr1BhcWL4SN5qPFGmsv4jeQ+Q/XwY/qkjceor/Y1TEM+nZtSEfkSj8JiuL3pYe
x4m9ZSbUSEiBvmtlO085UnFiAwGVKlIk3TfcEvK3zqqWLPAePAArM5TRUuQUQnp1PbRYAQsqqvDC
saXMhlVfp6VTwqMR7DkLRB193ffLC7u9B8+Jqp21DK8dKeN0TRoG62bFkHNMTq8dqUx/QCtlMP/S
0ShMsn3qdfXHglY3nXYUFiLCNpk6HziLpHjeiVmClaqvZzN9Oh/Ik1Mvbp5CQi6AjSNNwZFkxZNF
LQbMj0IqsZn87PEXj+5LkyKVerb7Er2En8JJ/0hleB/oJRhxOPxBjoK1wWLkjDQKUlpslJINDjrH
fbMO1RWdjLoXUcmSjFTd0hrsIbO2VF/jO4EgpLhkLQm1vwFb4KOWSxY4aC0E38rzZIduW6xGB7Kv
5eGv+zl0lNprDUbIOkLuiN0pMGx1RH5L5vvBrfo5pA1OOHa3FooKqa28qLdlwl039+tDhfwA6EtG
ozlSyxinyoWuyjt5ldk2Agok8j6zZoxyv/N+3LbPAfqRKd1Cg0fZygc1646WTUVK14L0zSpzi3km
ZMrLw3jtA6hOH/ezlTEaod3Qt/X1fa1Rz5Us4Z1KF8uOuraVbi8BxBXqBzmIjk7KjYcH1/r64QLD
+qCxSChp+mPBthasFkaBtYizKpUqbpGASq7LJ4kgWGTGgg1WKRvUMIYk7flN1x/Ye22yg58Nqg3X
QBYAsCcBJCjCOeM5VJWSlzzdB7pZ60JfxH4IszEgape+WbX/IrnsxcVVyGu8GpYwccVNKXRV6ybC
RISJhoebI2UH85raJxycOPUOgbDHHc7R0Li10pEVbOvI7IOnsh5pHVnQkA6EnpCZZB1dtSdbFFFE
QEkT6Hcfk1sxFDomicjPMnebyWwOpplcROx8xxaJd4Ziq//l8Y2OF27BpcYVTeHqpF5KVCaszMir
5f5S3jNMJH1ayDLA92PQtRXvGq5MhK0x9yi9hLhZEKy2jTS0NB1QcLe3fVIiWs1Cdsdh8CrKEDES
80OZq/2Pook8mX4qoj1S6LoezphNb46oDQtNj43d1sUCwkPj6CNa/RhWiVIYaaS+mt1OXFJDTKRF
iuoYDbpltLXEG3N3qE26UqkJwmzy1xFuOkhJGQThfY7krdJhFK1rNKLzVp//Pb1wDWfyxT2gr1vm
svKn/4YV1/7fQQSPAy3JTBi0xSx9DdmBZWcG9t+jjKEAPzbQTh2lBlMwn/Ya4QsKQ0eecX4mPg+h
CKzg7ZMHsg8W9S1frVsABLgGgDPVHF6TwPgv1CQvcqw9bzKvEgvO3Wl1klOxhs9G4mOoDFrxlN4U
b7xotmmeHL/+bMEuWRKSQ81h7qJO/sL0v95V4SDSezMvwxh7j98J6R36figtSvwSWandVTdUU7ZV
x5wMG1y24fjZdhKjj0l8HNQFoRz+BtAWsKdNad/Bv5U1Dc/lD7se7h+noc/Vj1RsTDiILyI/rCMG
BjgUj4DzoW5iKNCcqkK1FoCsMr0wLQTPdnuDdr6hlmQ4sZE+/lORx5fQQro60bjydgw/s+bPJ5MT
AfKRIFaKtWDWrXD9YIDKXUWnlppCStRk4ae464p8TI8qLftgfXGrry9jE53Lku4Wxc5QEgw36kD3
t9joTvFU5B/NE1bBL44q+3oIHwS/umlM2z8OrC8HwP+RyAKlRJ1DOXh5Ha7JnbzxzR1y8yGXyqzu
5HEdgtcxvew3H8B4sGkacaWpSX8PItrCefGPv4HNmUtO467yA8oeMqJzc/74VB+zlR/zdGeLHPve
AQGSlMpDUnU8CrwZB5Jo1Vp1XJwcjSexc9Xu2uQ9DL/xgIF7+ANeaZNIJQNEIf0n748TZikpP+Tz
pU7f+grNTydT42LJlxmxnJVFUYKIYL3uw61ABwSqHe9/Rv3LGeD+MOqg6gGtNPx8i69VaWkMKRFr
WGkHvChP97sM3vwGlEk0/ZKqSD3fZw5PMDyf3eZ6dSDUblPaGcKeRnZyYeLxmGT/TufzSOw2Rw1A
jk8+KA+50J/nEzh/IfFtrkHXqS/HA5iTPLuHaCTLf4ZnYBjGMkp7TRtGf4fp+9r0cXC+OECDlReB
JLXvdMVU8yGR8QrDU2qReswuAnFRoAYXy/LqioziE29p+5eBoSo788ksCqOdTxU7+EdejxI0yx5q
Y0Pd798NtZDRbWzTyPirdY/DXDs/WDX/r971mgSHkwqu7zLHXJ+tygH5jP51PCd6/pwkIngLDINS
6nFZxj30KplADWgO4HMUgz32tILXBxAWVnuH18TGu3thQ3A7/qWKI5EpztDmW5AFk3rbpSDT6wVC
lPyIygEl85eeyVGJsEs1i8QX2agxF7FfWTM8/BGP4irbPOMo7IOKc8EV8ZZoZnbNvzWzsQOQpKjD
SSwFc+sBUIDf9VKFJOniYjCldqLdDUQdslPhN6Gz84+5r6gDBUMVfi6erXpOaiyCLb+EtnsS3DZP
xNcx6f0cp6WFl3yodO92KeN91giY4XDSxuOuff8Z/raGCsd2gs0AE2NrhyIIP4TB58G6Sp1k27BY
+X5py5V/aJUq3CJJAX6gUIcnJT0ticTfVKzWsXUCsL/QsoapWCMcO2zAgnD0GRqHjYtcYRLXtMrv
cW84TFjblafQMFPUCLlKVbamWNWAwA9CvyxcRSBnBnaFfPNdUafyIlrHnfWStDw+wKtjBtFuvfzg
e0+f8R2XJipVDbgCASUHcz0zyUH+Lq1p+ZYg+E+rNj3RPDISHy6sWFx/cB1KafrWm79YtWjmguAk
/8sc31SGvslv9KTA4MfeJu8ESX7LZ7qxD81qAbeodh8MBmvegwmLzVcBYjvjJySzR2E+RZZnZ/YS
FWntO1thVWMLV41AoquMQUTlKbwyVvNForc047SBglvQR8LeDxH+mj7i3HxvQSK9QoUFxbYUmPMW
WgR/2EaR8ag28oAYrUDQ2obqLQAe0YskZh9yoP5bSXOOexT4VOjdMVXjmI6ZFlpUhUT5e+9dlU5B
FEvWMooHp6GNycgRbc7OXuzhiFfuLiAOIdA63kw7k/HwCeyZdQ6sLPqsFS3dbEZVsQWpnDbNAXcL
J1WB6bt0DiLWzPYBDUStM6X6StqFBTOq3tYuw9fPFr9OM2U7K2HkaSYlJz71XjU2hO9M6iC3u3LS
Hxx+NVeurkaHJv+77AoNgAuRpB9igTpdVw/Hy83aM31+CudC0hzPWIXR7KTWn8jC8dpCr9+3YAn1
NYZ7xQ0N7sRgtrUXVoCXh0ZztRhTIdEqX9tkEnO4wf64wXGqfJMIoWaEKoBgFoiyPpXNB4ncUiMG
/C3TTbY2vHwNVD4tG95pV+3VlawAYk0anPWwvNL2XzoTCXZ+YNcaP2LtJzr1ej0Lq43CxeizVquy
oAci5ykMTzIJhCLM7A0svPrH9sTpA9CX99IKJIZ0yAA2wKerqz6ai/Zj+qBJW8SJSe/DSqOU5fZj
cAvfIYasWQSNebF6wfmT1W161Z/jyVtDMFNu33XCAorVhAmDPEcAOhYR0weIw0Iry/TolgIlAt5/
X8pdTMxiKXg4yNQrrShmT+V+gWCuBdVCuKicWNHCe9uy0GRWFzz7pj1QbWnpyF5FvZ1QD8BF8KaN
lRTGcYriZ1lIsUqzIzRamKxRN79jheqE1z0LBZTywVi2+T/5xX3xMBpA8vnBpywWPyN1647CKzPb
WTPLz2mPBJi0BVdG8Q3ZvOxN2NE3IyZGq1lsvZt9kC1uP/p36PhjxcSugFA0XjeiaroNDPaIVb4S
0inVoS3DIUuYx4aeNUDd0o0pWfrfXnA/jVFpBunOD0BavNBuvM5Dcoo4qUonLgPBhlk8SP9TFHqK
SyN7HlqLGPBSnj0Q6QVGkUy+WSMSndU5mV3myl5rAp9MskzjypWMox5XcqEGAwLDWPIuMOWb5FHI
17c2SxkTKBjIKGWMErFLS2oxEQQGezvTe7VkhL+eJokhaoSiGwL5do80ZBqRxsaQUhYzDx50AfyB
gtroXHJ9tTlTQkaxGSkUWnVt4i2s9hagS2XXYP5wDVYPxxzv5pVosKRn1pb5/neh+YBM4HbyXmba
7tqAPhQ6mwMpdk7evAFCn0decIsSKk61Hes4VBLAjh9FgKv9TV2dFK/diXM5d3phYd0rMnM/8VkA
1OkC1BmLRgxdCKiKYpB5rJxQBRm3qUefknCu2htibkXP4Q2ixJC08GpbU5BO1GbizT+MekAiQ1Rs
KMeDeZMb3QlrMd7rqXlChW4fE76DVY90wZ/9i66Thw9E1MdkvjX+NZkmZzY3hf5m0TEFYtNdLUG+
3wpFlz6WY2vr+Y3kNuz6gaZ5kxlrXtWPfVw+qmYpk7L30MhWG1B+aQDh+9fl27rk0WCYmrvhpJKs
AJuZRYkittZZoGMLHrALOwrAIiKvDcH3x6jtVnEmpjoCfomAmcjDJdRFmhaBekW70h9qJbfNaetC
ZpvvluH3Fi2h7FWDGdtWPW9Iphq2/y2WIkRBCylq6pY1QqvbDfOhOdD/E269GMDFVS5ETSV/Zfc3
vdY2eIcHukOcQ/BKZ2qkpTxZDSHO6RZ9fmQxi/qT593AQ9jOjnXMysqBm9NPRieOqvbXo0jIpdTg
/ymv4PoBLVAosdTqMZ9fQtOotgRBgj/IPlXwK29Z1u97oTz0ohHBpwOAHx28bAxj82ip1w9IlE6q
pzMD8VDVgXjMQHmUIbvvYPy2I+lGGUQtQ71I8EufQG8MIb5kk8dUa1UAsdzI5MisoFyTn4VrrC60
h+YVL+RH34s4glPVdUjwKrnt/4izzJp5zYCyKfCi+TyYuitknBRwREpTHiNQ1ZqROooN4swwhXwi
FqIEy7qpHsO59lWhfQLmce8rsVQ+cQVpAT4tmQuzz4RWYvPbmLLVqrgZkZwP8lr3xB51mkczI0RE
p8ApFIPJEyFr8hd9T+PFMFODc2XY14dj/qOqMJzfAZdj02Zn0j5rOJf8ZXoj8q+EQentLiddrWWq
FN8coPIZGjX4ojMcI1Ks3fLH/seLZFI6iSRwkIxE+quTA0N5DmBMwMHsxTM5OPvpAzICUQ16MmFm
vlwVsInwKVhcZJBSie8i85UtaHX1ESppAhy1BbkF4xxUn59fhiXaqHoirV8HUK5usTptsRA/XTZN
VeapWFYGVrXmDpSEduMEb06QiNF6bXsPw+MHyla2+NJtOkf4IawWGlZcEMBzj9KuVFk/ZY8lhnvj
rF9+TKOAE2CP+UtbrhKFyWkHmrE9M6NRX/HES9PS46mxq4GEIJTzNNNXiJcFLyDHbhHU2jQKqv9U
MHoSWP2uPkTGukWGWwT9gOenxQZoyr4ry8XO7ZgvF2mF6PKmYmFwdOscYqTR3+8ZIpk/GUybRJTJ
Ba+1tY5d6trAInawCkwhx7ewwy07akPJgqpXSR5OqP+0yWlAoyWorfAfvFZPo6xWvIL3O240jyBt
AWz44Qha2rrFZGRk11mDvxpsbtfe5CDhRCqUU5lKFyPwAeNMEitghVo6Nm/+9PUQX2Ecz64DG3cY
gvJbZmbilPDQs1rmU6ishEvxh8QOuIsfWw0HjRxRr7gdJBYNkMurVxIFBCuxZ9cQlVAniUQGmx9F
7FLAWCnJNrSC9F6yhriE2QEeRHMl3a6kNm2m/h6HJw7NxM4zgPZqvLpsZc5D0YqgwoRXQ1gfq1QC
TiUiJE+kKLvzLa/h+sXd9BAEVVGLiRZsxG8T0+PChnayK0kdSuiwemrnGrnYZVhfRQo7hkNkMIbt
EUnssuJMJYrogKZwf19tXBNGzqqaIfSKCgEz0+pJRnoro+2DHia+LoZbn+cvSHK9VPEDJXGuOoxa
YynBU+tzTPUDpdbsP1ztNwVVjOHrr25rfRFQX3SP3niq8K0vDr1xPV8TSV8+x1QAuCTlZUM0EDKu
5OPSriBzyc8AQWRFfsMj050Za1JLnAse8BqdXk0YTMdbE/ftvf0ojy6IIAn2FfmpTyuGzTnn8hnI
O18I/pUfqYUcJYrfmntie84IgPSC+zUjAq0CYeV2R9tMO61CqBpITN7yAwQgHTIOB1Zi35iCc7EB
s2kUyeLV/SwzHbSapO2bkScvJoI2eFwrECQsg4fhA3gqbFb0asoXj+3zXFpQAuU4+GSc8EDxeZIi
nAHYk6CSDiAjnAEtOnoTz4bXU+kbf6xr0BArMtK+EnWc5MvpqpuVKo4RZqG8/Hc32xAhsdVRF+gz
5n8RybaDJ9jImJs/CvwtiaiMZZt8ASno4XPCOAG7wj/krORL8bCxjSd23+JPi2SiICfkosHfFfZk
/qF50lAprZfSIspsVH5AkkEkoQFVKxOoMpHZ7uQvp4M+8XS5TTgKI6DktD9nnEN94hm18DveOP29
o/+pUgB9sLrL2xlEssbiHR9Yjthl6t2AHP3N7zZtF8o/MCuJtNc6zmCHOzVLCB9QKxrqYt/LkXrm
+s9+1qDI8WaqfGIBLd82aeug32p5pLd7tdVBwBkgRNipVUVJo2pW7TNBhcLnpWbu27xgCc0jMeM3
izSxbrD4V2YPDMTJVH1OZJgDdqedm6eSPL8INIngmaC0h33GC9PFwwIN2W4smV+sRBFOCcpn0WIC
ialvrExExcXpn9q6Og0+Xnzy8+fhlBIk3CPpjV0xOpd4an4bZYVAtmSm+wD5bPBruzmAG1jT2V/n
SiJ53COFRG/UVl4nJNILhZurDR6toR/Jz+HGirqH8LOvG+Gs2UrAN43loZfbd7yMkatmVUyZXNtX
LZp16rgO1VAc6v3z1qWNf9mQIE9GpOw/9ZFDblnfcVRpBnV1UbmYVJjY8tVEeAdGP0ibY0qA/7A0
K2fdWpWsR0MCkous1qy0iU1rNlc/QhjAhfXVdCwODRxBtv+O6w+WG/3LtysD4EM2WXMX7uIMggrK
HFNygO8p5wl1GY5dhb6J6XkpXOgqzOH4e83kAqOb2jSMDY3YMx0ZT02ak5d7usE59HyDg4jNfWe1
fmJJdNHVWIdeD/Bb5H0F2/pRekQmxA6zaIo0xTkybr6fiXTyGWLDqQUpcfVJF2zgIHJmWpoi/Bn5
93p7ruLYUjvcKkyPmA/qWGvjjXDYi1rWnrUDDZ8ftGUUni2/MsueNpcdKeSyma6IhIWJzeVodM95
wYQXfaZDjRgjp1qoHDYwkIICJkiB9lPnxfLFT/hYI+2gicw9Y0Kl+7vgq4OvEPACj+wf01aES3P7
iISsHS/GhbwDfo5qVugG3MiQKnKl2xEjN/afT45bO9cy9Ba7IWhVE0ky3gdpfbxVvx+cMsEuWHv6
7pjpN2YpWd90W1N2DXVThAm5CjZVsrmFjSKv2PN9PsMiWHXRpBiollBEPITGZrsCF7dCdYosLSMH
5yxanUNTf8RtATZJVxS+R0ckSzBZDvVlwjG6RRgTbF/cfzHMOb9PAqhalKZtJfYemwPXPpGUFzgT
ypvDw2K0RbFaVZHRmqaqs3wHJtrYsSXnSw0HCu/uBFzwgZoomJZ3qYkY1vCCulIpgRZXx1nDAkz9
bncEFk2m/D87SzG0YDNq2G8j3RKaRB3bw6M2fTG2DEDH1EMLDqUXFl+8Sl0P4s5CTH3M/Rvcwobc
EEgrtgJxLo8AmMo1b0hDbM9n3oUMwZdw7PCybPLbwzw4HOrLjsWz+H4OycGQU2EUuH78OSEQHtlL
5koUfHQ8ya0LKh7TtKS1keIVFvGTfQfGib0TouPaH5Rj0s/4EbXMlOYvowfx2dxl5Z75FpdeLQQH
9JAExP5EeJz2fKxdoIYyH1kKOzcmVWZdt4/ESSejhe7MkSI9xed3Z59dgwFB4k9Z9nJqEQKxaX4i
ChgUjb4EXi9lxl+gQhQhxvdNPjj6G6YgE2jHEWTVAHKs3/WMSkvPiO8ru+G+hmWJEGjwd1Mk05bx
7LehPeZLDBaDWEyX24JJytkijFh2SNLjAgZTHtnVDbWy2FMQ36zITpzJUou/eDbkIBnZqjRPt4YJ
mrKgLbMuuIWMuWsF8xY1mCUCWZCfhnx0B3TZ/gkfTF4SY635kg85F5UeMviNAdbqiD/UKdXSoDOE
B3vJsVx9Lw60W1PbKbaopqHjkrscPoOp8yagX+GwL44GdbeSgXyXYYnydGobxnPAxSxGolJ9/gbg
z9DVJE4qK92nX7kCxnVbeZjiDxIaOdW7FyfZ/tQbrG6xca0xgDxF0yBFeatZekw1Mlg/VPjzSIVh
pG3rR9YxAxT5gTcjEqg0DTiwB8ypz8D/YSjXH/YFcPD6JzwRkkCiQjCe1WpcQV30DS9vWSJezpIt
TELoctfuSusmF+whMJPH9S8Xj3KoutXhemNBcTOhztFoFR/2M4ocJ/5U6TB7yRjdJekQfqCbB06s
D4jxXHAWH5Q757EQrVXKtP/RrQ4ctaJvdIVxm0n2iHmgVTnPsGFRRuT+Cxk7utTYibk/sySvfdhH
5r6ruFhKwUAFn5nehgeSMNdQ86n7v1/oJ4LYWZG6rG52Bl4n3M5luH0e6cuboe+7LwyvrrVwGgec
vjO3FxGqTSpu1TJ/p7QK2ovh93wYHdquRB0rb2zA5mKc7oQq6uscewA1JUVyNu0s7PhyvC50NdpB
X9WpkauVLGND70m48z+EhvJYChUGDVfEy3sN5wQ3U9c4xdZi129QTH41fFyNZ/UJ/DiMWz/jF7s7
Q+yJUUSB0KQWZmT8JHXDuNyycQKtr/rwgzSsKxBwtx7kRaLWXf3jeXUEs28mGkTNeT07QRn2INcp
LD49OrZ7uuHd9544ffXsB19sEqHqUyvTEwWkJi2XOwjOQ3R+KxLHaB2cfFnT0M+GmhpRRPsIX7d9
gMFFUDDwAEfZl9aQtg4NyTWdgneQ4LOVW6Do12CdemAUNJyI14fJPG/ko8kK4sTATIB7jbw5B1ue
FFKOKjJwSClNX5mLsD/iIqzEJezWvmtN1F5arGr2FhEvQuO2Bm39ro7g/p+ypYW6oshcLQEEKSQd
TFoNZh3jCnpyzVq2Gkfqo/QAbzhToXvfdSZ7h3SfgTaTe3rVopvOg+tptjvNXBVBNdESyieLGsGX
3gfbLqRAS09nFchA0tM7lksBEz9gggpXncmTO9O9CCwsXzRCbVbkIwU5ga9MAfzg7Bfn2kUABS4O
1h9xRCmQ8aGsMw+UMKT9LoyQlDDMLWNMhi1e9Ato+668shR6pA0BFcruzzuDwYIHEM+oq+E82ftg
kSaicJ1w/oYtf+o4E2T5EUhwVqDduzMcy4S84X1DWHkHlBSybYuM6ZXCMwVeR+Dj3IXWmCKPlpQd
kxcOunX64STAEak7CXz3n/nYAke+9XqL36245Ebnzi7IR7yycrhpYhGESxabpN8B8yRvow1rgVGJ
3Josp1RP8nPIseUIWZChv0Em1/x8/MEGL1BVt1lmBB3JP81y3P+bff8N0mAxsU410NIj3TVxNiaF
1vTl4mL/G0jco9ebBlgtvf0wSQ3HsPxMDy75U8KX79WfD8TUKHvhgBwgwdcM4k4xLRz0laAqE/Hn
p3Lek5k5fLmKQsr9PTtaN2bOPljdD8R624ryhcrPJqAHBv3YuJDRt4gzRjr7Ex+pAjadEbjuGQ3J
gUBqePDB8Ep8Fzrf6j3pr9MNZ9ui7Yst5Pmv46JGkc7OgQzuT1zGAO3yjWdAz1TzBxQNtHYAvGTw
xtpu9V8i9QNy+C3FHHMnXfOnQsD5kGI9Zoeohja5+eAc/WIyqGepWxTkABxBld0kCHvoJDqf7Jy3
ZP3IOD6K7kaa754chsCFwFiy0yw5ZiCmbUkIslpAgghFtOzjri/E1YxqVDqqMCS2jL9svYjeEAqk
2lIGn5oKQ6FcCWapKxnuPckWJ2QSaIYoAeyMMIkYh6x8sT4vGKp89VdgE3Gs79q1GEbmUCzopZWM
myAwlG6aWmvURxmbQp+3d1JwjcYUg3pIUPpmgrMOV42vTL4ujfcLh11ez18odCBs4M4HeyfgqZNL
D9WVzVW/uUybn3cgqz9qNHzW94U51BFwgaizAhapHYf6CJiLJIrnHSJgVGYtabdYci5kwt8WlN7P
6sD/ur0x2psUeICpJBNMQPq6yfFb9JTsCBmAlueokPhBboKIqym6t5oYsdrcES9dGTsD3cW3MOFk
Jy4nwjpYHz2vrMjleb8NPCLdZWwDir6R4mD2UVHQHVyssdTYmek6IC0L369ZX4XNVY+CIjMstHR8
ToQHnHsqrnzsWRT1BOtjDtm1pFTrLldXwRMAdQq2v5UWn8jMiNjpyFvH3GWLLADZImEQfHUCSjia
Shjdx4r5/XZsfbJVQbYSzF9bHOSMwUmJXkWo1XkshZMZEtjGXOaY29X4sYaHH5Fj36rlpWQt3k72
q5Qh24zbHYj+t2L4ku1V1tX6EXcg08nQHTmD63WdNmHsfNyHORFAIKoqCppVndI9WNj6sjYpUnlh
MbgyBEBZdUGltsSqhmhat7PrWRr++WlXfZv0F2TV5n2DXTpcFkHYrmB4SOLqNXZit/XM/hVM55Mc
FEqyMN8o9vZUQTyAobsD1vmwbpnN7htyyHgm/EgrSkBRKUZOKmu7kXzgDVRDxWpbJ/eJ0tODQXcJ
6sbMZQMuxPX9Tg86ilL1/krz8QCpcn+D6cqU5YpWAyzjRybgNkge1srVHFOsaLz7f002FdYXo0lJ
pz2RO0eukkfEIC4gT4kPpjwbsal49Udr5JnwMG8grIUWcZMAPCks/3axjfWcO157MVuD+CDlTb9L
Zm4MJVpozUsJh/qUleJaFw2wQGd7eb8T8PLhV36uQ1h1pmNJtUbvz78710MIIRPv13Z5hRMNUMel
LGwIrcyhehLwLalSrnv6nHEgsYX+eVcrOqms4G8fYulxiOkY0+g8oOEb4TgxuejZA098hFCjAM29
hUBVByS2vS2z3h77gnGjAVx8kyzPkOltuv5s83TlhTzSYjCV/OZxURJCQPbX+r4yWMIpKU2KwjE8
zHrdADB1Cfm1eFrUssgN5yPnjHbLE4aqLpK3WNupBs6dXa9zeywFlimk8ZWbe+i2CF3hMGn1Dz4X
wAJ7XC5N/luBDsPsWH+KiqZbftZR/YKOOtKEI4XAm0qG02nmrb1egE55+WHbhey7TAKJ07SrPRxs
9zwUUovA7GGAslEkKiMfWoy1v+d8q3+KdxY9Mkq4r/gIth16hQNQ+6izNFeBIC8QlqiZMuLEXuwS
T3Lq73wFpgLGwFhc1gr+N3IWdRF2GnXuRKyksH2DWA2zzaJcT85FGyVE7hcSl4qNYqZdmin/JEzk
ZimsmKIlPyJDwgyG7s3wFdDuYzYqV7030KVIzwHvvOTO7HoIDQIyiRWMPAiB2eNCgpun3XcGqgKI
UoWHZRaxf3lfd5G0TXLan9QnRfYMGikSzB8z41G1OyicvVDsJve/lX2cx79uFTpnd72eT+lJ3Boz
qgbQ6Ld2JGG5DY4mW3QgfrEM7je4qzroI6EAHnptFTq+hMTsMV9oYtSeVEMvYehxUJB3vVYljpZB
HPwhkTP50S8m2Y8KfP4wKDgXgN/3pb1jtmVN2iDoqXXJyMyMy/9yWU6dfKIM7FB+vfbApU1AFZ2w
5M7bhH1shauPkmjBLMsMx1wGQ4hRuKwfwTKv0dvpVPJui5L1xBn6lp4wkX9QzFGSlln8JilBHfGc
URvRfy+HmP9BYhsCb6psCSqQVKLP0mp5plPjJ2LXQIzDGoMy9RnDQWljuQB87FTs0X4J8N4keIwa
4m6HqTtxLS2Ox6zsgaQAZ3Swfb1+smCNLQM3OYYE9xqvmtDVARlcSYqyeEeISZ46L2oNYj2Y5oq5
cR4WMBvS3fXULCY6FJ9LxUIyX2DFaF+GYN+R5VtcsHhbLZPx2VGp0SzXsje/NH3pf6Tf1QS57pq4
Sx1IGqugk4ke2RPV9YqCZYC8iS3VohPTSqZDVlIBSdIanxpYCfsjVxn6GAmdBw9W8Wkt5AguCefH
Elg5A/rhOMmdNEq9/zybATQeE1K8uGocfRtFNB1289pjIcjdWZmWcCWxcTmwh1TcLa4v+QF3RZVT
FuZeqzORnAjLY1CY+oOGXeAHXug0E/LAW9JRcZEN9qPuCKWi1M9UG533xFnhGmCZcVt05mJePBey
w6K40yhTCHKf8+wMjDVCZqRI2VLoc/OQ5DzNk6nV4vDoU9Jr4Enb3YBtYBxc4qWGKUlT13MLdYAs
hUqjSoU9ErScjvNRyl2Pfp/3MRFr6GVmmYZYDUgX3wQxBMsmx/3ctGlHU4flFGBUb5+ggIIvrlWl
y49V1hePt1E/jFs8zaPMtkicdqfoajrAZ8SNIwItT7AcshoUHRRoqCqQqFxscl6voswYzGRXG2Wr
cH+flBp8nsrFGCT5mkX4E5CY+fz7Fniq1tCAmMnZdwha5Hqrh6Y4oCBzL882qKCcgzrKO9jTG2AO
LUHNbIh19betVowGWdYxNHbac7Agn184neUi64MR8C4kbTZ0Y4UTbyDQoEBE8A/SXD7CBG1fwaGz
qjaD1nLH4EVsKaKRUJLj5xTEI3C38ADcQoYZAP2comaX19Mcl5EdT69uVl7CMh28iNxQkQa3UAfl
uH1r4/CgDGsOJqRETfgOAGowgltwKcC3efQsKNcErYFYfj9TaZvzsecXa+SS45VoZ/Axsh89Vtgu
EhJFStjl7Q9Hi22BM4M+GK/DkHWZLIZoyqR19GOr6+yfmkKuhRLjZfr4VJjUF5KcfQYJggl/+VwL
OUyCpCptDTtIzqmz0ObuDk43/ddLJatLomaqkQLFPE1RYRKf2ZzRruxLhRzXh4LQpjKiAB5aNvgx
v43jI9JShhRNUstVLud8yN4iwORcIu2KEbDtdyH53/wupoGgOVN0Euq88sszMh/MjEVRFdr4p9oF
spEajCKPmbxNEzIqGqevibv5i0Ps0uOjfMRdki4IXtagq7/NIMDpYtDrBry5VqM26vK3NHqPspCY
2ukWaIG1aUV0maOYaOSddc7It/FUfqVvr4kuCuUJ+ieyw2djFcHsRu4H3eX6aeRiou+MWXOemgKH
39fX6seMZBldI0+SXk8ilOUxw+HbuJ9A+tpPJTouEm8hBdumYeU5M/Ze6Mr0Rg8dHTvw41DXKlS4
MJUfIQCLXhtRPugQAuA1aeo+r+0r79M1VJIHslQnFF8DQ79ZALMo/m+XaRwrt3qWA0HGtDxOzitj
4C1Y0VXUQKR7+WikscOqNvvYzoX2YCfE6/PvBbqhP5podwLrRa5EwS4LsML4h3xd8SHEaT7K1cm1
5Snuja1QaIiRgiOizPtqzlx3BwZWTYV5NX3s6KE8dVcTwB87xmTmVb7Sd//2bQMHeUMbKaY3cd23
nwkQcNg6NVE/xUgdylgYKy5pebyFDCfpVtrRAsYFkXlSrugFirdrK32eAX+ydUvI/wn+c5i1xXGb
GrmeXTb//rYtpdgQapvwcMYP3KWaEmaHMxdwFXIBi+5IT0UBoa5MN4x8a/S1XuhGkSOLHQHZo+0F
UTC4Wh1ROCCEz1h0TNXaMSqQSe58cW1/roi4RbRZl0z1NAKV4289XbyV6Pg0584qZ127B5qxPXZM
2ZC1vf5r1Ebc1Ylu/f0Jg8QSQS19WiEMsu+AYv/9oRAE567mhcA8i/ZOtw/EOmoyJMkPtfstXwqW
iQ9w6b0QA0j61/fuGL+D5GCXWT8IAn5IG3G3bAn+URiFhKsooQU2ES0+dYP1i85nj4qnErFcE3O+
9wB9p0rJR0cCiXLeoNqgudtixWujGrVTBhbkqJNLCMjhSIE3q82bKz+4pbgCC4ViepIDNOgAPtA0
D9QqLQVqB/5y4ds2QBkqJLB61aayVToq8rZEo1pkw9V/htAWpJk7rYS5mhwJxn8abxOYt49AJiBe
LpEsU9AphcBskApkC7s/Iwc0ogvy+X8oZPmSqZdK2gTdCG3fZl+TR3R0kKRUnZWI3jzHVY9W0X3w
/W3St4/rbeFdZ/h1sAfcmbLpF6s8hJ9P/ltN5/Ut0Tgzo5FvtxSlTF2ny+2iD8+QIkIqpqUuheyp
p2LPddK3ITo4LyfLck2TmkhbLhMy6tJVL4AuddlUTAYWR0gEY2JGMYLF16OjQrfAXepIgS1twCkk
fA5g2ib2x+Wyg9jQ21V/xSEFnJmPk3FaL7M2jyYyO7T9JCbQUziBpe0jYOi6bKAJkkfO/xz15Jfz
c7YE9A43RkPaCjXnF7XS9hZwqsM3f7pGD5ZARFfuGQqN9GnIoumvytF4CL7M57DEFchgl9LG0DdC
JQ8sjAgMtmwfeTaOL4CmBhxQ8d5f8ITPAoFKQFJJsODB38s497kxIXemWmwWBDlL/TVPePUU1bfa
RqbaDZ0BoV73SF+GkkkOqslpRAo1HoSN74+1SVnLQMhfUrPKnVa5jcO3x9GhjxD6s0fnPCsFBoh0
GtTA5pMf91vUuP9k9LUcF4vtSOdNN6yTdh8yjbwmL8GL33kEjG5R7D3Nnicb/KTIBK/Q5qRFut97
Qrx8PuRek9zTthZXm7Ey3Wy8/+RJ0Aj/X3IxC33gIRW0YtQE1im/syl2IWytWlDYKHOxoOIZBWMP
fwYN0iXK2b9Qg2UsOI1x7tqYy0M/XnGOemznYRLy1CKHcRuDW8XlJ5gN7GjD+sPF6bFcr1R/BA1r
CkCNKmP9ZOkLU249thTmz3Z20cl4S4R5/aC9QP2m6e7FiZ39HfNjBs2jD5DLrnJN2V/gvlcoETLB
ePL9+/aCrkFun2L2xXwIf2fQWAqDqG2wuPCa6W8zK37XW4ReWMJqJ0gqBmYesjPC0h9uoRCG80MI
5s1hxGQXKHX3AIxEVdIplhWhytneFDg1cHl5OWYjIX+mAuvvRgrDej+KrKEPC3kK/yeFb7ekaO3E
K7a0v00wlBdE7i29Gmr2DPicvuejeduMWtBA5iGpzAsfpP5QRNZVrGXJEOjp71vzB60awC8datdl
+CkKki9JQCjfUjZ1E57BzF7bGP+Hs16wr/8rJ09Wn6xrBHSdx+habsHLi6EUDXpWVXi6HTObgCSF
Lv0xjJj5ICCuA7S9vZpyRl3cxEcmHLeb0Q3z0xZyCH+fGwSx4F9A/OiCxENE5htSJno3/XWU/TBc
jdp9dNHVcBUJ4P+FECOK+yH5P+aFVRgFMhUk7vF0eAekhLB5f4nn7ugkMtbt85chrTXzHoHQqhVd
e5FoJq4k6hFtVEfZtJhs7PBsYCSbqooH1nBOF+8cg2XbnGOwtQwocW3TDKvuRaJTt3ebvKQBhbYo
Z/loSJPc6QpUnuRw3DVts82aS1m+++bd+K7X7B3HHo+QQnqAGnabM50eAfmzyg5T7D0Iqjs4utap
zFPzIPw9iNeDU5UA9ldxbt4vOcsaUGzjGAQBvrpmv61ELGOixBkKE67FOZNzyW2Wu+B3l52sFVxE
HHua3mqpho1e0hV27Ln9dggue771u1GBcwNX5f62iaqqllXPe1wwTWRKIL6ZKLRrJbb0HJfwnTMp
5+/TsGvDjb5XUNB1e9rvKu+imS70FF+iQnOZZVdiSIghwOrppm4TxVyCmMM5tO9XNDyG4ddFHNBt
dRxiVmIv5yhU4Phjzchv+vAZQ5sMzcRcEZxlcMr6AGfHp07m3NtlO7xnKgLy1MY/QP7q2Pkw7EAO
sBjlpkPqvEDVffpcgPUY1mRkqU2ykJ0ri8pcOhq2oQVb5xv9O4PQ2YYSDRBi0Dp2xZifpH4BcjZv
1Osk5sApm/ypuXsEhcEc7cmOV12fzeYQ/Y+cSzIGWqleL0PDYCFO2GhYBEdZaeL6+ecKmRpD9SYa
ooCQoPuZ2gteVsYMofsWhWafSWR+ORATjSX9iTFiXy37ibKRAZPT2eDrlUNadSpidkZBFHbzd1Wr
Bbd0oMaX29CI1/Wv/wDIBT9z0MjIMdABXqekAtvLaBi3jToDo7c/xZDPTdBrOIK4dr8/kOsUI9gc
FMd0tyUAbFdbMPSMfxEp9nXUqVhkUaqs4uwlJPF3nsKnx2Oin+5N6ysvaI5GnzFJ+ugyntxUqGzw
r8370Jn6WmMY8A96l+P0/L8bCcgLC5F5Qk5ikSl6LymglR6Aa8ivlziFQN2ciJH7Bq8bsT04dO7o
joIToiw5zZ4TNeB3q0UkjzRUlKSqPORQ7syL2185xD6fA3/KN/xGqEb5BwDALQ1jobSj/sXyBHFR
erJVX47bPEs4uOwFZOdUq98TyJr20ErnI+YgrQSKot4APoXSodU3g5HZnVD0XPdVQROCBLPvNRtM
9mHqc6S0B/zdQJ4VcRd+FGULDHGM7fSQXTLjk2I2P0aRzZK60DSnyN/+PBz4/UGF9GRUQmKByqQV
bKuo6gDXaqWPpk/swLSfIt+QzOwFuwPQqqwgemL/PmT3Gow1iFmxdADT65yHrpkk6wUA3531Wjbs
7NXYYHLd8Efu2vrECANYPXyQT4WP1Mhm20CQ81aO3KMA+XAqLH4hIvSoqCUCvFwNvfRWw/guQLLg
+gs0RLZuLGFsmHNzq+9E7Q5WQUoGtO4G+m+K+3PuNq6+J5DiQ9mtmDBpJTK3/isSCj1AWsNdyt+S
muD4FaCOrH0xNC4cLsC1GEmP4o9GeivpLGZr6APTsnWBNAYm5p6u4yZsK86sEcIvtzmJhT7P6BAl
dCewo8cB/yHmK/YVWheCWCsBkZxJ9oeSTHHvytzEHDzijqJD8+FgdxOrguNXrw69LdHTZRbN0SQ6
vmombepxE+Bn47WD6Cbr5NYpXIWzj7n0/86mt4PvKdlPBJYm2/3hja+EItf6bgjH3gPZKPo6jzVC
8HAr4h9xNBb4Kx7BZ5Y5fM1uBj+PZ3FP2OXsyjbMCNIdFp0bFV5iEggwCs/gMNs9UEMYcc4qZTar
dtNtAWlHJHjIpkOt3XAdvP/uRpLhZERPe5Z1SW8aWNSzh/hvTkpD1WIlf0dTdHYegSFnknl05j52
RjQ2H6ETR3k9UidKB0l7GcD5eBPiOskMNAPW6rIooa2ymc9IjfGFpaD2Uf5fXLekS0itPqzumAjf
l90lzmydXlCEMLpjZfaSCPegRcyuVt6sz1JKoZUBumEgir/UhkTHQA2qpbM93t+1WWe+aXDgAoCa
3/vfeZuplDdaqnVL3JiviHUtjIX+SH7dDFoHlZAdKGuIfonNkiADf4YkJbSHpMJiR/IUvxChid/0
QYJevINE5Kjsv0HaWXKXEEh1fDlE4I2o8a0YjbhHH+ybLiRjJ5iCCzuBCoV7ALi6VgMEpOt4GlEY
MdEHCWR+poYeZsii2T+sAyEGxq2Ab0i6YX9K6FS3s/wFbt6yifoyHuubzSLpvPHDKyHtrFh5HmEw
i7zJ9R6PgVO26Vix5RCDMtHfzPoPSo4hXtjhuzFLxyTrTf0f9XUOXI0Mql4qFmeyBu8J+nymVnbv
OBE9dz4jGD2/Y7fw0m6gqQE1Ru39m6VB1crETHOTbNQ7XmE2KKnH1jJO9pjwf0QP4M/KhnEBTNM/
FsdE9PXnDnJYt4ERFJPqgzufYPCcynWUyr3sLWrXxvj6FQVmshnOgXbgQs3dH4VASAdGQJvzBO2M
T+K0u/erlBAJGjAYgKD1ZP7ueRj9HM2Q/q1OM8KOycNDqMTBUr6tGY8BTwo0qRbP9lnWyF6AVfVD
/G3bwdxROMXyAP+N1vF0JpLcby9u2dvH3SlgOcmGAZzcNWYNmtR67iVfl614/rKVJsFKacZbNxzz
gtQ5n4a4vdB1R84ss1AT3O82S9b2ukR1LRHsCse7BEZYr9rNXKkJPeCkugpUVqo7iE/lzRFU+iNT
HFzpTacCDd6G6o1JhAkIvXoLKrHrq0616ypcrsn3CW8aYTHi9cKSdkEGTATpWvvSHftJ8qHi3dh6
L3MEuZULwv+FfLDqWf83nEPEqdac+QcJGJeqX8IZGZCbP7siASfATZ8jSSuZB1Krt9Sv2IvZvdf7
KWDKV9obxXSrUppTn7EA3HEKU0vnsDKQQcT8Kak1nPk+e96nFVWRoozMgp07lUM+pdKt/e67Ulpf
j2L/UIlBSNrQjOOUbCEmg2aOERmsjdtHX2bA/3icAqsUDE8nMddD7LulovL+ahfOp7oh+CWHixyH
BcIOef0/G6ZrAq2VqYSbOvB6pcGQEl0c1OBxAe3gUrNjiCxLwtCq/TIoJvGPDcfJhgqTorSaTXgm
GdnyGzzL8Z0JXpiwYTUbIxk9/sVtKHgQeILc6ORV/MIFikvxQP3vrgx8UaedFsHWpDxP/O2QaoQY
mTF7cOjmr/qMjxbVDGVKHIhesgCDtVoQDftmwBkP9jUOMEa35kWI7PUFmcl/Ayq0u532sHfkxkNR
qOgtyjrRfd+O2ZAJjf2g3qHu1UUD6DXD5XIR3oN9Tm1Hs6uoHLJfJBOIzhHf6stpyhiKq/jl7kBE
9a+PtgvjuW9/ggOSHVKbyKR8QFtUigorCYp00CZa0cqOnNf1v7U3cxMnClM9HnHSyMLJ6ZJaRvs9
h39v4h+FNknpEiIDeKSUSiTHmOkHr0ZHBzwV0t4GNZiL1tdr5JES5DpIxpLdnL2O8WhmS1QZ3r66
aSxHpbJ/nVdoDLlbEnnBuUW8hiPVQS4EKkzUT1ZzO08otq2v/PNCSDu3zeJ94m5iDJr4z/ISaSIc
6ojuaEnzgj4sXdRUK3T3fdLEgbq+3vlFPzJ6m4l1CFL75tCOCm0wMQx8bIHhpB+CJpPz5F69H9MT
4m4yDKCNfDGWfViuBKAi5Y1Ol9h9Bg15hziDIrMs9WCthvgn1Ef55X5THpuRlEHLl2VrmJItRVp1
7NSXF683zt6rP+gg8/ufwCSfgsUe386OUO3ahYf7sLu/LR4k4Wwt+ppYTsMOz6JKnF85tIIjvpfZ
OMMDfGuI3sQOkr3YSrPWMo0WKMkyXWFpdcbDlWhUDfSmrVtx4rI+vypkvIKBSVJHB0Tkqnq4Nqab
u4EMH7TvQPCzulyxvzy3AUCWhr4CKEKhN4I+b+oMN3Q6yvTvPj0vXVc4ZxVMLZhd1dCzsTuNK2rC
QZ6srMK1v/+wzW2XHL8KDIiDerWhYK7zoHpUTwh3TA/NwT9WAKzpx1ETp4bHctpiyQbOWGNrRvlo
XZFNOtvTBrNuiIeYIaRXP9xPgg/VX3ZiWcIp6OiX07qQAiU7dPnisFFQStaSoBMbAA6Jg46/5jbu
4JzSORWNjgBbknZYncWGvEJuxvwwO2oFw+Uzyd8FKVqnB7JfJJYpoZLxec5yhqz5W1VJl31Zz12U
xQuIGsk5Qimak4J3hI9rOR1IlPS4Yy1Gc8NTLc8DpY+yzIsIFXMGmOxAJ8XITT/ala5+6dqPB+He
6vilPiWA9DQge8mIn1+Yjth/k5/rFkUOPlww9bSvIHH5PgNcPWwUqNc8gedZ27eheGNR2OJlgcM0
XGQStVTVFGiRk318MpWmpKGNK8eW5PPR3o/nQeROgcUDXYf+GcXGLDZezqDK0I4qE/V+1X/y7X2e
Sdb4gOG1O3EIicxmfhwSANHpbkfMFg3Mk4hA0JkDWcy/ZsPnkOL/OLpZ2qrWH2o57Zwy2+1JKUae
SKdcMNkt62HdJ5YNSdsogsukZ0vJE2qCOfda94DhL34pnDIlyqwlpvmHlnC+w+GCf2+Hq24amvGI
ff2vb1peKgkYjCJ3bPjZ16l3AW8v+bFzUl2mYyprayPaUSM/MIR/K0XtLSxalekWZX6UcmnMmRy7
DCCsOECXQ6S8hVMqnSfPiZW8iDOeVJ/L0tqscUFJP3SVyC7DhHInPi8ZgOuhtSC/adQJuqX9yEBM
U/LmfOz+u2uH5BQ3Uq+3nkj/AtQ76bW9ut6aeZEi8ZCVR4TGVk3xFITYebkMSm5tHFI8wt3QGqd+
W5PHAgs7fO3BFXwYo6gSafyKsIrBX6R1xVgs1fZyT8pHA2yhm90H5FJzfXxN17K5DXdkSgrM2cIr
TjJGRODhO69SfhAlRiZUYAT05qbogVzNw2Lh6bckW+ktkY2Z/lObRRDQyxKAphHJ2m3FJ5fnYB/X
8bbGLZvbgqLz5JOC4QmTF5RELL9bw12p5RdK4Ef9NaNBBNySKQOOjr+xJGpViGZ+gNpIw5KEaTRa
nPv72d89/pJ+B530K7LhUnqYShn80UaPEjOcW4sw/HVtHxsIdJnBVg/bNtjaHcB37opdBB4EIin4
lWcpNi1KSoCRRuFW47h26kQRq3tc6vpVpkovX42wDeKtPZvqoxLB1PThqKbfvk218mgH1+pJodeK
k48jSMSy7NwnFdFlVg1/3gg11lq0MSPPE6cNyJsmeUqqonNgVP1qXxXHLjVEtUCrNaQ9upvMI+j+
TOR5uSluVpwFP1mGf3jfhwJbJgM1xi2242Qfb3MTsvQozJxOBjMsZQEOFbeMbyfV094dd1HgBEZK
3Fxi2XQrXF2NUACrxDiTnZiToAizoseNag28pbz6GCskhsr3p9eUlA8FRbMqDxpnWuyaEA0ithjV
v+TiuXQRliVGgBNuQIli2wuLXZDwdxUcdAZnt2oX8zU5DeoN35KcpJieh1XAgExNnRM1dI6uEZH7
Rd8ab2Uk7pY+kRQOyBlHBDBA9NjlteNVA36aNoREGABZtlA5fXk9AKh1d+r0ve1Bg4CvApbgrZQP
zIpyXpKVYi1Qn/av86GwS02094behacnpZjFPA3m1qDRLlGwyTajyA5T9VL9NPf2ocZY0aynK1XL
56pzMEAPX2o4+KTGVIp91xswxjj9/ash5Wt0YuIga3AoVbTQ9KU2hA/D0LmM++9AoimyVStZTSZ/
Fn21IAMMpWWVaimNBol2pKyqqZVKlE08oPeKGbgmG5sZE9+3J9T1FGH/XJbhqMvV7srxX+aZyHxB
aOT94l2Jth3GZ1HD+PqzwESWJUC8ky20y4RX1N8gkmQ+TIWayXNXLeZSDGtI9WAxmFPTXPKok1CR
Ce2sdYFqjjfV2s0W1JJhwDzo3uoavm7vo+wQPUoDLiu9DrIn0jLb4jqcoxHopDq9+znfBgUbrvun
+ap0WznUxQHWclvCm7ubT8s7HPvziNwoyJ0BQQdvcvqTG2Zu5seGD/Auwb50zoZBDK8A9p0MMD7O
pR/lFGHWe+g2nCItaHbxs/N+V/1TI+5v28rM+gutjesWH2DvwQW0pk8zQ4u/B2hYELxjWBFVw/+e
qfOlWnGejlZXy0rf75+YF3z1tncintpDNzwvGRVRjzKZizL+iHS35eJ7TmtLDyWBUNr0S0/DcO75
RWDJQR3Hs/Q3y83LlsVCatdtpBCkRJbc8VKeyT9C+0d2x8mBgb+8F8BL1rVTeuBL9O/IcJJ5eWou
gCK4cAmzySbjoburseya8sJlgkKqgkYZyNoNPek8X9jmKbqXj6hQly/U8ULnitynp6PfnkdNZg1A
X7A1xzXKJnR2rEevW1qNgwth5r8nU8EvYEDqZryGNJIEWrWaRzfZy6ApI+r7RJ6F40swFqV8nQfu
nTt4qq6MKAPq7DybBrtX4RWp1Kyn0VgSE2QrAFY9JoAVbIRLWIZVVjdYuWw75344CX65+O6ivjEw
vsyJCxx7fneWKJ082XV2orymbAQN5j4ljF+S3uH17Su0PchJCXpwZE4VKgD+dnCImpayCWG7WVte
3zCg1RYpq7QfMeZ7Y40tYMQ3OPFNc+hrB+8GJgrlltKva3sxkvOk4gisG5PTy+zKLEdMR1BJ9yHe
UaGV7ZT+5de6XwgrAG8Fl4O+VjOnZekh+3DoFkueC1a/KDg1TPx4+ke866z8T7HC9QTJbsgLLxYG
uvMRrE6U5yUoQRMYuJQ9rU4yW+qQNNn1ADJX039CYxLuMAkX49pC9Pr8KauGihWEEL/Dv/rF0D27
qxbA5fLIg6VtAn6AS23JZx0RmDxZI0RfJgshcmJqluBfCpiK/Ugv/0BVTaWkUc7quhpern6VkyRv
YF3OpurQck9+jtJD8kfyV5OK8oShqxOOIqfUVZaKxSCPJQw4fJBgVVWIWmXGHW2Qq8egXc+akNTa
3i9bYumLstfJuq/d09PoEc+EbGwRj10+zFvUxv81igX0LYqj1TADk/bGXeX6WMAGdrQ5bXSYn/wF
GffA18IJifu8eMzvrCOdONcUoqR/hCudky0mdUgK+r7XKUgg6sKWD93tnbEBrVnVhPUSPt9LD10n
lZW0FrC4Ygv5Mt9VB/AqtscTiaWpLJy69SqGAgtkC9j53yZeHThdYznlCeKYVAXtAv1MndM0gP8C
QFyhCW/T+GKASsShWpO/YPVFxZnHF0LWe20dgSnAIDh/lPTGyWazsthwoSJaNY6d9XP9daHQsSl1
YQ4FrVH2zkbOTKQNAxlFFCG1rgIaWoBzDzrzcCQ/1dxsjmntRG/BjkdV1eB5DnMWRi6ARTo70qTO
RK13LrTKW7u88sUiH/24FWIPZpdzkUxMXZOkDUHAUW8BolREX6ac33kXq50dho7w97OhDxGciGum
NOXFknMu5SwY8wE2We22SOrZPkwJYZ/nFQqaXipi1PAnFguUs1gHOwGF/1ljwqGFCD7a9aZov/+4
UJVRwAtfuTi7dVOX6Adf2m1her0sBRjyyIrdYa0sy1J/sPLyMpD8e0KEF1o/fdoBE8Yla8bOXzbK
mC3VMsLWmE2JHoWx7lvDAXmwUZ9uJaDjzCBrChrS1LK5XHko5Bv7l1LkoR229UvaJuIin5tHKBEp
bDGtigZIhUIdnJzEPHhIxEhxJloBoMD45zrS4q+peqYpdvCVywaF8L9XBGaAUCJ3N5hQwYKJ1qb7
AWozt31AtlYsPR5vfI4cEYCXxQBcVbXJI5NjZDH0uZHs4bSHkfiCZ5wSyeZ2vJ/npF693cjAtGRr
6f2Dvoza7/rR7L876VeoKPXs7kIXVk3mNkzPSts6zv0IlAXiP1dKvHWjQdazeJToan6hybGFVp4I
u7L2zaLTZO4LV9TpL7qnAgFwZEjhlcyhVI679h8X9k0x51rxKHD1C+hTO9GK1WkZZaDjsaSoXsq4
0MvAuceV696mIhwAOW52ByG/H+DugojHz3rHzwAx64W4IsKfMohbA4XmXgOCsGy7i7bjGzOOKGOV
0TGLseMSL6KqaJ5t4AAC9BsjQlvwG2S5mOSwEWVPZFQzgWbFP0RU8iclqqMRYEwYdN+b0IT8UR5Y
XAPviJ8Qo+aY8naaAJ7w+OpBP2LnN6gIkqfzkLWzXPqRHg4qeSStviDw+mwSQWuSoI01mGRRN4sh
orV5v/qUWkiehp1+NMpAhInvObcflxdL3RL2bQ/7ft5RxwdBN4LwNrTrzvjSvtc+noyk7kVyiILo
wE8bWmVdEOovZwqMq/R0oCfa5F81mBEXd/UTWwiDfY66l8jytYym8onERtLwBS+nZ60CwVBKFaSW
HEChPR+B9+X9w43w89GYDiffR2IqpM0yS/YWwFdcES08VRKC0tgkARoTRhRQiaKkmtJv2iv1jEdR
hSgU3cg+HQwR1KJbOAeXoIau1VS0z14xT6mWGi3DxRCq3gnqZnoPJ1cgkw/Uvd26UabELsmtAfpO
JfNlyJOR59n5bKKF0EnKhw8bnRKzaELJhuAhdRT1IWhhemdB6ErTs4VKAiKJTJWW+8OPRs/cxWdZ
I9zTAVH/C6stxJyAxSJDG38+3WHv1Luzb914Ijzx1llKLMaUe02r6BfLyIm1c9y9lpWSUU6ftJHH
tCbsxZ5MuH+TbyjiNIytfH6dlj/oTb1cL9z//13RX6++RXr/YzDgFJAmbHf3KCVyIOjenQhRHpf/
3XyRNpXkUZhSnn+Amu2p9U2Ou7R6A7FvzaMwg86s31Wv5f2H2CFXmb6exheYKrkq/lWRu/2qX1mW
74n8vMn/42kFhbOVa1a2V8uAGYu16yUm3oSTR3x9Adt3IRvz9A03p3iKhgC1pguzU02S5KHFcYJ9
RWScWGq+hvFjVj97jnBKCQ0X+wjwgb02QDYaaj2iCB6jvvWAxenaeYBGIYfF58yWn3+wRws8YDjH
2ibUklKCUaILYJAMgErrDRz7LwQt/6Zyx+4qM6WQlvDHqgIHLjV+/9XTXykWT/WWyvH1SHrkIzX2
XRsDoI6g78uJCpSpnh9cjltep7VspPmFx68iC9sexpCPBI4BCtLOXV/fWKNvN5Qpy4SgthmDuKec
m1JpAiybK3rn++CAAbPTRkFeKNGU/S55RB7wNIjQdSVakTA2jSmmDVWlbEZYcjoGB4Ve0Lp2F/uZ
TG1/YpNLTHHczH8y1LnJ7OjAd1LhzaYV9B3H3OetLX+Jl8FZbCkPq95TsDpYBfCeOFShAyWuSZkc
TBcapJkL6aq238MLtslX9/Qku79ibouylveqftU/AsQarUSbvVCGq3GUxaDpgpzrnedHNezXCGHD
1zCM78kj2dmpTsAlEPv3zmLxKKBMJAssxRpw9j6ROjy0uwy93xB3PshPecv+xFDT09oxRh3CS76U
BAl6ieAvkOWLPJnPhUC9s+KWC+mocp7m6iCnKSEdcJJrKZrv3zWLsDCmI36Hv+2E94AvJ6TQdysP
/6zh+bx4iwDC7FhsLZG4QVIAa1YtrHDx2oSlcg3tlJ9QlpiW67LMOvbZ8vFL2wes9qZeKHlF9FX3
To2rdNL7ka+foKIh21W+Wj2hoWishIf1QbQaVTMz1KkuEZrdzNX0gbcksZ2gxuHd1LfaoSshYdyS
m/ASXkbEq9l4HKoBgDok5W4bY0vvLDrRv08b5BAD7rnRywQY/1H1WQuBHePBaH8LIRJ9PUA82WIn
DfkHtNak9cEGp+z/UnBC+ael+RgEEIelRo4aOk8y1PcJtrWj7PV98xjnCZ+9y56y1HEZ8uc8gNP0
KPHGqYRGwJnpPVNHePiJhEREOGZTwNf7tTGxvYle2SW3+nJmUEobd7MGox9GEBs2rxhza+q8GOAY
6HV5zltcgl59ph1OqRtZbuNEwx1Jv4CPddPMkVr8jKL+oAc1q9SqF/reS8+Hq6pO08P2msuwJOYS
EUM8OPxAVDAnvPqpRS6oXsR4rDE4cpy8lCheHY1VOOzNhNTFhLiuWZwTFDiiokd2I38k3+Y0gzQl
6RJAd9XIdtAFK4j3IYlUToyq+HGI4bk3TftA0WDosmW0KXImArjNf3dl+tGv3b11CsJk9hdRQSjK
krqQ7fGyH4QcNilUwvj6nc91e2gBvpFXdVg9FAD992S8tS1D9axyD4hmN0Gcq5volwTYkNKUHAGS
Pt5sjiCNJqdcPHUB8R1OEhovchcWlzBamHI61M/MWcNxwuEhaNJ1vqKypMquEQRnxwHZ1wlMYy6t
XErMh+M7jhp9M+PyFWPudoMRafnA5bm/zRRQU0zzTWqDuEYHDdCR0ydP6VVH4o62lgke9rCL2JdP
w3fy6RGASdEqraUkezjTpULlm5vJYsnTy68roWxkCZsayLJwUBWWDLq+jHGraKHpzgP0Sf/hWlo5
klDehRy693mCddPFT0lLychHpfyk5A/VtO+6TPaBHz1X8wpLN+jDjMwLFJ9zYuic7U5iEkUv/nfD
ym21mdO3paOADHkhP1TbxaunBlD6onwWZS0Qx3en/DVn/e4NZ45J4JUged8630Ka+FYAX7uGfBWq
mGWNCO3jmqXz/9P35Tzv2/wMOdxmKOvw3z+fO3GvKOqY0Yt1iDa8fr23Lxd8WMwRZeVd9FvqCf76
gp/qb6b9LOcmHLrG9cdFA7QVJyhlzdo5fkHUU3adc8RHsZxShfEIUO89MhGOkmVE1Uy/af08reWt
lmHigjwqYNKzwvPuAL+JcuVR8JBYFDGYTQV5Q8EMDyInqj1uXhYo7S9D822oUCLvQoLVdQRMChiD
NqnXd7MFa7W4v+tChSFDE9Nd8TqXkwtkaPMynvrf4F5E+rVYN/WUF2IkThEhZFQQdr9+NmtBN+ZO
PLaoqtTVdOgmvmaYBXm/w222BVHS0mqcCf4Xp2Ppix/kHj1laNdpDJKVupnEeuAF7mKGBxKBvXbm
HiyRXseO7ieWiI+VCp2aEkRhRFV4gZVKlSJLwukUnl3cyMmRETQrMoHiZl1jfnxyHBRhcYvAoFak
JZt9ZWPK5rtjO234ticRBN7peyhRb0M1iqIwfH59a9CUCu7iQI9lYgmWMSARel+N2Qb0EqOTfgwm
+UEF+SUNxtSNyoBN+qtkJyNkOZwJ0a88JOGWbODEamZQ0NpNaxe5DNAgAohmMXz6I+iKi7z08q+I
z5mnYw7gS98avtuUg8OzXmYEUDq6BdVXHCd8AhHIrjtzyA7CV53OpqoCXlJ/6SR/G5+z1PQEVl0U
r/5PkfBGYRRPXIqsTEq/3HuRFbnbpFCVPRJkUVc51V5mgVXvcicffggOnDmtc5GdMBY5hsnYap3k
4+UIh8icHF6JTQqkTdb31xBCwA1WCFBz8IT/kXTP4Ax0Ron+4Q4TvvxWD/jIulRiGOpowRSq7qgz
aY9OBv9Cok5HnqVlq3wJEO19MtGQNZScSouWmbIgX4NINnAOt4uPNrCVp3saGpI0ehUC+nhnszC1
egWtQGv3shXmH6Aj9Qo6PTGKCefr2z3VLgcmZ5BCAQT10+9Xlj2P4Utyoa1s47eMqvU7wHIEgL+j
HkH21WYEHzAYoQODj3Ow1hJTkrSoQ2FJ0N86BAYY08Q48cxtGT/GqAdypzKXW8ulmR5Q4ZkZRDZr
nPTz66TIV7bnXTXV8NWSJHPOLZMPWRn4QC2p4g6ANOodXhpAsKgeRKZCVcg/3pBtrutb8kng9DnM
aoJhNHqXj2zm0XfD/Sjnj2UKO/EoDiwivHug9fldHAuTyIxJxpjUbP6jjq9ZEUSgYSQyJcxaizan
q+WwywC+TjR0qy/73scUJzsag/hqKx0MSiy5zO75r9Vbpa33oo0XZ+4/x8/bsF653dkDiCHN7BJw
JCn+KCqU4jEVmBTAF/BhLVytEd6Ge5yL9oCP0/BRmtosl2bpZnj7YupQzmkIC+YEbnTCY6HVViNb
plvzG1/cHpCrwCyoSr2bJ8gytTgA4qmfVZtSxfsNV4nZ6ty8rxeqGdSIP6BzCdOOV1Pd7pgHWfcx
voKWAQ1TuudfFhkzQVd1G4Bz800tob8MvTL/z2WoXtgIdSwL6hrCq9Qzrg1HiecWGiC7AHG30y05
9r8MylApaE/es6sW5dEbcdZZGRqOAM1EaybFjQ7Kee8OM8TVoCZMXAhXWqcnZwTKLLZ7Zi3GZJ4Q
jC1otoyfF+663Go6SXam4PkOiwPQmlOHXXv/1BRt+QaeDd3ukK1FMN6+W9tha97HSIGafPCYRB1C
uKsdjeZWtfiGKqrK12qfxto7+XXXsEWTtPunHVAc8CNdxq6858+2Jo74ojE19ZQ+8peuxm47ptSe
lKGK+FTx9y+82qhuVQT/Gh+wswU5/g8IThr6CKFVicfBhAqpkdsWgX1N+WvQcO0vGS0ItVZRTIgt
vIETR7Xu+A4dz2tT9lO35R+HFW1gk9IBE6t3kkRsGdvxvQGK6lE55OHRIb3hEzZlkioe1L//1OJs
VbI7eFv0HOjNFBtRsSycDfAFcRgAc1B3gM+xdIFWXs7uhC0Y/nCzbJeM1yl4S2cHlbVH7pmxKbum
vxi2sB/pvad6kCZhmWn352+wVwpmj9b+F72ja6QdHxlOm4CkCPHuXRMdJ5SXsGqpntnfrf/Z6GH6
O0dOcaVc3rt6KoH6QVj4whVN2wzG1sDEawOWM3ucBmll72FwD7e+7U8k4d5s/zYQuDtZeBgaYypm
XolKGxrl4TZXjVqepIOScVyJwWHUGMkdPD1AnTE+ZCed/EW83IwsAqmlVJwZ9TF52ipHkfDKqBbQ
PDi1foQVBkuoY9N6IHYZOi+ZnTzv36d2BaLA/n/q3+MmqP8rFXWNl3X393kWzhuHif4vml2UtwcU
uBVSpBIb41nzaYk3Fd4+fB1A3qUAt6RdeZJkhWV394MHLmaWWGYrbtpDUHM2o/qL/nORHsCe034p
6ct7tNVSIBpLCOfGaEw54b4eMSTlHRoG/tbbjx0D1v5U9FD13KStT/aMh3I+COB7yYB8+q1dLU+s
kCj/7zDBA4ecUTda1PmFSrSrINvkFz544Urjc2spnMnm+BmpfcksV9kKi0LWVn1dIVP7SmxaLZi7
bRJ0+FWL87r2hu/uhriDXNVhORW8wl7thpQ+M+XCq7P1BtRpTDY9NyaC9m+3CWbQdmoHuEzSkxkx
QLWg2KbAIykMXKfuAGaLrJ0TcTmX+4J86met1dktUjSi2pYBTfM8QFdgbga3yurCe9n2kLg4ikoG
ZO468Muf9nIVqKjtxNp3mT3DhkRCfuXxY9DpWvYpjzC0ICfx5be3jjtKmFDjU2bEyQFkdSaczkeb
zVUwZbUILbcBUjfegvxCau5DH4heohIWW10YG3xpZ1bDDIfckkMoLI3h0ddiGeikWoCayJEyiQK2
D2xFG63a0aO9t16R/wbTni1aKgG+7ZDlkkxDGGQ6NX/jhjucy4my9NfEICxTyV2rj+5zcsbfvGkE
ENbRPsWK8AnwJiDVVJ/tj54GuaZKmuE2jDVhBf/r3paLkQc2UXsYeCW6hTTfOXz2aT+kuIDQcFKS
3Vy05Ujv+h2iXXVMpbJPkhXEbhlHzbm5uEMPcs9Vi5zAHUhdvjGSaNf29bZERqVDBy0SyuPHWdq2
G8PK5QSB5EUINIyXsD0LQHk9vuqRvT51hHt80CVSaYswk9qpNUMXmv5h0uIhxqMyzWXONey0xlVc
+rMtNOJCpc1gbfL8zc4NYNIRtZGs8GbY/LqN/oqxlEcN9wRaHVS0QlkfXGOgmcmeACkwXIAfS64d
YNSBoB1SXftFq3IfKfshgp+xFjoYOZvYQEH0ULlkNO6nzCpgkfQm8iPIuO5kEJUuMQk9//jLeh1T
aAmYehUH7rIxm7LvBog7GjdbAtKwzRlFCnyt6wgdGyTnAgvx3tQtc8b92KreSWDgJdi24pOoZ2nl
HP+kgMcaDtTvYZZ7cZ35qwDyCkyXiIbThfkLR5+h+40eF9n7ff16NwuXMrtZ5X6+bd/6vlscmDeg
c/h7CiCezOb9SRGyce3Z+HT8gYxjC2WufbPTAuFHc9iGjEZVNbm7TPMnSL9VQ2Ixxyvy9OfqRDWR
4FSjr2FhlktQL7dwYWAxafHb9cV7AntOlsSrOL64plZ2JpycEoitdUn3zspPmgM44Iz8nZqhHYhq
jsCOmocCfxwvChsUSHUvD//QodmZ0jHZauRO0qXIurh0AbHfeABzsGrUS5sGSQ1LnrWZW7/6auR5
yhGLGY2GZfMHH4Oagc8oQRGaM5Bv074SM/0WH+XnLJgkeLWHxgzYQzHhk0R6lL0UMqrLAWPgVbiX
zvn6RRaw3p47aKc2XnB3MGyYo35jOdW9jNXvV/UbJCVnGLRU+dFumL3dSPH9yfSLnQJkK/JrwvPo
5Oi6ftGy6qKwpLc1Iwk0AAXRPJJqdfbwDLH1I+KvMZPZyA/9JCVWqEvAzB0q8GJ/l9uvpVKbZVnk
2Hy+ZDsXQyBZhYEH0OfALLXyfX7dY8NpWOx+uy9+SoAemKOrWPllW9GWAVD0JhjV62ukGG7xA4Gr
8TdieKcHsBvKUWjxeoRSW4C9KwHXoy6FPfDXNDZJMlgETQer7qD75x+o1pGUzqSTtSA4Zs4PeO5n
44EXmqXMVKlGX9pCyOOKcKT/AEh4JuAAywIa4Rc76UZ12OLK5oEUeSv8AhKUUqldl8xd4e/p7maf
cc/5MXT7zTpUF0F3Y1NNiNhlSwWXsQfn0S/rOAECr6svvt1gaSHW8h7b78bimxCJJQZaAo+i+oBZ
nqoM2El0ltUMqycMQseBh2cX/KTelYuLdvNA1jBERZ90FsiiPMOiCYCL9nK0zhacOZtEVDreoPIJ
9XNVbgcPUL883KZU2UijCrjbtFpXKG3nS4wxP7P23R5h8KbCfhgQkRRqw2M1nv3A+noqrvUZUf8X
alGSwBSxuNuvKj0ec29lvmPG1ub8JWULRZeT7sfoQLvlv7CvIWtmm/iEBe4LINBCmX7NXDydelH8
wwMPRw90TZWQxLcqR5MhYfwh4OuC+UUL71+wCLEk/34Aiip0IsPALZz5uFAOk0OJA27OM1y3J0Hk
HKwqAZAbQWtLXi2r8xbuE8XWVXnvlBdnbDA8JxK3tigvFn/t/0t7n7O7igsBcxaGTvBRuI+cjMWC
2mGZiWEWZX3MwkrwaUeSzyVk85dGpSkA3BUSWQqnkG4zfJk4IWzNgiTXCmfvmWgCNQrS4HPJyu0q
H3xzXwohA8Kg4MNNKXfHqBa43i72zEkXg7WPvu1XFWeAdZ77iGlrIy8GGJWHyyTB2NwvFDftamH7
rMyHicClXULBas2QD06r9CQq8VOksAsMC7TJjzsue//NUgxx0GDbPIm9VDYfDh5nr/7yoTgmvwvR
HJ06VnVOlLG70+JTowrTSlpyCKdJNBuVhIW7n7f0ZWMs3+PAMScHkNnLf8rW5JdP/nBd1uc8CjlB
QYg928MNIoLd5cax3mPxIZR8HyDma+0YzhnBh6BB0I/wRrrrPB4MLvVAmWVD6lDbS5xednLgLoTx
7hCKtaYdvWYjV/CahCEqI5hmyNyFrqm6ledTwTz+adaJzRoHSVEvc1yzt9OELubvgdapPpc22Xus
VkoeJpaSAA9iZMZ5NhPssh0jqG5RV5fQVHRyD6X2bnzQMoVTmG+RGTtN5xG1/9O2UXZkvo4sGAau
pfyf9ZR0/ZzERvDTCpl/0pSXE41bvDmqjDdd+Wxit3Q4yKN0qzLcDZ11FYl6yWmEeq8XUIDTLJim
MCbP6jMkEOk+U0lAfkexdM/8oUALII5QGuEnEtUplBuWYsqVFBq0mBKRB6vgqhQiVqSDBFBbmPa4
A9u725FHeDQwVUVOJqJ+YDmOKboN+2A9ia8lNc6bI/cwIAveq5yGJdMZGHmTSy9PS/Umz2NzGtiH
h7gGC5dHqhuM6ph5Ky754WwO1YC/GbpEgDw5K+aEsgfJNC0zn6EYJEA2xXUGjDBm8OU1MYxNEJIZ
oGb+vOnbzIulqbTizdb0IbbIDyyXuz/RHNYM6/z7jO5ro9l98n+Y7wp85vwrQo/gJjGG+ixm5OZ2
UTrzVaNot1hnYELLtpbbIk+so0C+MND3l6PBU1TWlerVxjUMNx1t/xpPlxmETtS90S3rDuDhndi3
2YqhMNpI0oux1SJryrrBAGcrKwglKiLfXstTir752b1jtxWy5h4XjdrM/CS8b4zzqgYfguOFPqBq
dhSTCZXPS7uBkFUPh6i0orvAgtBoSxf3xx2FLWkDgf3OEPaJ7Oyt9so8FbcnAmgs85JXhqVQyi9v
DVsu0E/LhKZ64eJkNaWmpDIKkGpG4AamUs8nxVB+KFpgXWDanuOdFRnpu7zZhIP4rF90pESVeNr4
bTdmUD5x3fA623mfJ27GQ9mo1+ar1cPtSlUGgiI+uCI5IQoJTv2WHExPwStbykyLh5NdW5Nzp7Jg
HVAi15RloHmD2oNZFT/SnOYkO8hvWodyQf4+ltZdEoOHuNATqvDloksJLQkfGSZz7LdAyAwnyoyS
tHT3NJZzqz1peZYur1FE9l3UvZMMK/hv+rlrjf/ID207Kqn3Cw/2RHZgcorlJABJCPA7nKpHcxXf
ZMzL5ypJe0g7FVgrepCzocqNV6nI6vTOLaxzcwSUnckz7MXcZq0Z3gzlamCWSsx42Qki0b5fiDqf
76gMqTsbmW9fgx9T64VR6Znqmybk0HU9JoJeXbzvETzeinC67c1fSexc6QLKxF5C3NIajX6N+bD0
Ww2sfsYeI2Raa64Y4rVpVlRqDsZCZ6E3fmVq303qTXUiAFRu4GzMIvs3jnzp4Vygfl28IgJkOU8X
ra8eRiVS4TGIkQ7wNvMICSUtyRp0691hKIFQxabIN050cUFXt3IXJrFqlFPKShfR5MVBmkZNwA9H
Ena7xP0OJBnR9z0v6bYkW1ZuvX9pom4dkjflNFy4HXmdm/U6Y2v5AVyfLMU/l1LXjSUSIF3R/ITJ
ocBxhe3PzZT3d6n5MxF2TLJmUwIHaBajxqO1XtVXiSVkIct8k3yfd/miI80F0h//ZPH7+jBQLaL6
SwvI3AWXQ3TteKTmmv4FSCzE+KyWKx1tEslzx0tkehXUqEyL+UoReIopXRFdPeXctthv2CCkSgsx
we36faSvn+84gRKCIK80M0o4AnSISLUk1lnkcu70ckIaM6mwqqJ8YkInNOnOvNj4WiVyRHNtCAaf
WuCoEeYK2ECL/BCJI7go9B9E3gqn8cY5vE9m8WAlS9Ny++fWHnanemCFAoT1E55uKfz80cXuQXe6
0wO5qVWB+nzUq5wp6JIEfzthU3fktj6f/mKGxgObJhCpBq+WjJ9ySyWeSdd8KrpLlqrRRTIoR/es
w3iy6aM0Bipzsac7ndJd1oT2gqsIEWpQm1wnJS+dYgFoLRYMvMxhwldk5CP5rSVYIlI7SCW60QgP
7TgWfzE3JAgEBqTR4RvZTl4d5/NB6LQP+XZLYe5fwdMzTirNVkZo4JEKnBP0cexK9qTMozHLBRxC
rmwtGLMeHpZ/VBPYD26lF+CdUAGTqOzC710rSLiOZ8yK3Bk1nGLGy2+E9g60QpabRwEhjvNhi/8r
WDst6+yTWamhoIH0mN0lzmLbfqqaE6LZsWlaa/tjcWCtASOBJir+kVmFYGDOXiZAXevruDuyUFvf
9uCJXrUmJO4KfzkIXRUkIR5O33d8BAkxPTRKatufj6W8ere6+BA7KKktEqheV7B2IhpG+8eMalye
cysUpmNV8mw2F1oEJ1CZqPnz6ByufrpiUcycwxhFMHCtTyaFgfvS5Ypcj4VSTv3M5P7yRe5rKVoz
YH1ufRi+OK4ZQ8etM+p7MnUAYGeDFLIH6A5LJ40q/YZTDS0rb/6PuqI5AzpuTrCFV/w6TR54mttF
8dBr58EYiJgZgaDy0IuaPF2hYx/0ykQ2dnfB/3+BdFH13s6To5u54jq5ng5SYEjDQY3AQK+9wrNc
WxAj9o0bImxB70hSiUFOC9QGe26uPhtteIrHmVBGbafJ7SlKvPzjhOZ9PXPgj+2CRPzPlcqvCj4u
Odlccd37TTLNJG+9QpsxILGkieYPnoqdFnOSFDW7vn+PSsLDs0McRf4NYORWvKg6ngaYllsWUNMU
D7f0YqVU3evAVbAplw5LlkFDHa6spy95rV3BQF3oqAnTn7FSdfklMYBEBMMj5aAWHe5aBACtIQ8c
4fOF6BIyWx1lKKHWWJVVb4FAYxDp8cpupILarJ27nipD8rT5pjV+yWI0+kJYA9oaraLnmg1360rA
uaZxN3o9uuDm64dgLTQlu/mkOqkNm3kHGogEyTmElJhET5G3AJJntd73MwnpcLkcl9d25RdPf7EP
REFWw7lhFl5Ju8DvvFqV/E/wfCLhtXKZjs2MDprSbMkBva/D3CxEPAhI4K0ifbD5teA2Zo5KdXt8
NP6Qx8u3TCyecGAKZtyhOCKkl5wsnc1wPKf2j8o3mgJuCJVRBItrZwz1++flVPxPnuH5N6XB6Pep
rAgp98vnvviiPBOUhw9Qq7+tBEJiCNLUJrcT4qX2SdAhv+ciIJejRA5J8G3flpqW2tKy2wt/opfw
iX0gH0f1Qpnzub3mo4ArQaaifbzAipRCntgapJISrHh2RgUD+SeAWLJMha78oFZINU+47SK8PdT/
g/i+A5p78x94Cw4/5DCeVlM1Q3W4AMG2ifty1En3GZbS4PLq0wh1HEKzknIaz3S4PGFcb0WR5CoD
Qm5Djtu/ZGYE7bOsfGY2hv9AeBFL6OeFvTNyMi6aqLSMYrGtrPNNMFo3+oUsV8xa2evxENRLxW6o
rVOpGGY3wZyl1xqKZQzwzHZWo2/2NxjClTci52U6hTuRIaweDH+EbP4ZgKhOwJgSTKY0/zaEJRwm
a/m3BdUFS7OxWQB9Qq6hHRMFWwXll4CnvIrzV8cDbFgdKmXipmDsJpPS+xhTkNods3TIMJULRlz6
sX8IqcPHhxILDsQpa2lnscaBhqODYkm1sgyNC/t/Ic5Iq+vuosfsY+MIjjsWIhscRlWVY6PwoPny
jv8EPCrAvznvctC7beuGjiVNnQkb7EYgxZbgnkutx2LnnNAeH8wwU/mIKuIg2As7vblCnDIpXv7b
ZyYdIgcPxt0YL1pKQcCq1/Y/QLHAP/kmIcMowrMiRSkO/sKmCkrfsHiMpvZ8xJ0F/VEFHL+xjbdn
Q2mF5t2NSUx7Q+g/ci9Y8xGT1VtCSuEwhCAvLJQIz2JXcNQLypeUtUf7C93b2GVgmouKjEtzCA1A
Q+BRQ+uwkGTNkTsVdk6a5NOIP3N3lS4r1cvrcII2UmTVjQl795jNtkAWahgfAXmbr15HFho8Vqme
LHYsUcTfoQdTwygBSk6GCP8sZDXEWDpilBUUuPM+5Bs7cdShd6ypJ9IPlQqEkjramVEOUysypMqS
AOaECwlM5sop6OCk5fdFXKjhU+2Jv1Z4/GkeBAVdOf80X6iD52Z9l8+ZvQIoUqVfewSCXMrEbOfe
MeXh0gdhAWsqnCGYEyUV3zm02wG9J6VstOZl/a/KMMxKRoB9eplEwOwOoQel0Vt4T45GSxplzDOk
y0v3/I9aBg+CVwp+gCx/oi8tcAn2TB60s/0PxA9y715m7q4JmoiBu0EuIxWjsJQ1DfTfgWrHe42/
QQrrRO3eE4q6ai6lM1wLWcIia8liZ4og1iLOJWvoIA/bRc9Kt/FquggrMKbNhRFlHX2RPHiJ0BUm
Jr6mMJkz3KqLRWMvmNMmdr96GV0lgl/IRTzMhTYLwU1iLx4cJnculaKgD3ZlYL0Epme1OCeueuUo
9BIkZr8h1vaHWF+DXN7I8vj9rylG0Kqzz/rgQ58lEmGwMQSvRL7NZMjPP6hUEToLAZ0LvFPrIqzl
8P9wtdgSKIZmus2dNTNukyWmWnu1QbvE0v//S8JWM+6RH/sEnyQOynPge6oxO63dE5hC5A6iXXwz
M3XUNAH9fconjULF4Uoi1xhNtcOzSquFTnXZjXW/ugtGlVnBGfIfsQxuSLWMnPdgkdABGBmkQuPE
nIII/mq2KwMwh5gzHIcaYJjdwMXOBuXF2k9SZqOuGewyO95OQtSaqEXUSf6CE704jUcKLNs1kV+J
oqZdH4NsjxBrQLmM80vs8uTH+5RfY/SXCDA7YEUNwimVLUWw60JGQvzsb14uOvndMGIouWL0FzLN
fUSczSdkUCWVD0j0Gpvpj3+fj7/SSZD0LIeH7cz9NJ+Jey9RCsodSBKprbC+9G1HfjYgsoDVThFp
XNA3p+DMQFdFD52EJrU1UOX6B5TvE2iTDPC2BgP8MxnwIy5vOlnXddw0gjl8IR8jzkgKSbQq2CyN
1OMCJ+qeojzxLDLbgDR8G9n8pNivHr2msKDDKg59iThoilklzoe4NUHOdDaJMBx/flgpPayzK1Tk
THG0CRRtKUvvkJYOJBeOHzIg20Bz/MMWOx2Rc+O/TeFwtNJM1nZzzpbB+RlGm2FrzdLgJPQyyaIa
IVVHtltEslbmdVuLkCjw7wmXpEjEjBDnHbnHWCk77gmWaC35gqYVeYFehQleoTYt9WYQJg+YeV0a
3j7MfqkYkHffkE+6KzOZe4OhMfRvc5qqeSlVElcou27did0SMhhw85QrHgeGVql/057MSigau1gF
FddmlKHgTw13hO3q9q3lbWtqnfwW25v1Hz/EmUnQZ7V9rhoFRTjmOiHAexg88eAbkNQw/1g1qEKl
mhxEuRCHa+Sr5oH0Qx5Vve9JafhmsZpUQ/gdt9COUrLdqVahzt3yRO3UITWfJM5/TeUuKqlqJc1K
hLiTC0CofgVgrG935vn3HhNfTguck36IV3SyDLHVTnRZmPEjuONWMa+F0Il0T1IH6bhHJYDQoNRA
nJAYvo0Tw+FvXtSomZvQbInOe158QtalQFCfnSmLEa9dpaLTn+x1lj8u5E/5TB18Iu0iwDVJcWds
R75ZwYuOwH3M245iz/DQ1oYu+6HHrrvuuhVO5ZoN6Z/Htr0e14jHCuFFNGxtZhFUoSNJA/yWqR0u
U3glnfzxsEmaSGAhd46n1NtYp5vSUVCDbUnyBmAqakifwrVJyaw7+pyo8M+0SB/q9HLRG8CKTVg8
JB9gRkzp9dLugKe6nfygXeqBruSK5wS515VOEe8XR1qTIdIfmt9PquWY7159veBEvvA2iUerkWSs
kHgVLQqf4nry7eFj2B5hw4bIcUqFnireqdl8e5pjwWrjtgC0D7oH4C/klJxN/z/5Ixw3YJYkkBn2
OP/bl5YoQ9uPsCsMhUDzrVSjrCZRnUu8llpByi878W3IMEGxtUwHwoCYuLnq3WBPazCFG4OI1I3e
OAzH4rVd3tJTl+Xn+mXfzh+At0u3WZKb6L9amWK0cHrZWKjbA7BCbW00Yf2A1fDIqkWWyjR4cLeu
ZCO1rItzjz9SIqLfxV3mYAnmQUi0N8bmnl6n+9ev3BM5CuqFfIzLr0EPAyyRM/YpK/11qG0Ir4wj
FIVWX9D4ugq7u0cZumuxytPVSF34RFY8tK2V6D/08fMFC1M9LpmHWpgl+zuHXaUncXameNfiOt85
wG+a6aOROVr5DH/YXs6rfDenJCBQCqFQDH+6eQCzWtghkiCayrBfsMFFCu0LbOyRIBMDeoY3l+RD
H/xZ2Pr8v3gjXNowgdiEhuOf9vgv8RYycjtdEoGxqqsJ9MYrSTrIYQuLi8GPDzli+08fF2koRgT1
uZ/xwVwjMXBGkh7PidCsD7cQ3dz6iwYmpcj6GWB5InnVvzFatlwn5aF6/makXUAXI8gbiNbZr/7z
3tGUbQpjwqQlY0LkmiioNaOM9764oOdJ/qw1Gt6pacDqFzEXthzaIaYjIncqm+pPKWFkI4MRe4YI
UoZV/QILGWMp08rOzA5ch9IvEGYgeQPc1rv0bTcUcBRCPf3wcjI2m6YuClLVs5FxcKJa5+f367j5
ArsICPl0VIbd8ocyc+xEQ0JIun3EYn+zWDakxmdKWpnIZ1OZflF5UHgw8nwjkZiQxjm+EFzYAwwA
xshZZnlw3e0arWFN3CaUAlsJUE2QFQ1vTEnUai/L7d8xSJrQb7X5LLIQLZ2FezYI6Z44YH0br+o7
YrZGjhY17Hv92MYIINiVwhNwJhYaIqHz2YwjqTnBD2znoK5YIyZ6AdbeVWzKWU3B91oNE33oFHhw
gszcELuvfLJ/0VzQZOmQzqrvYsIhrZs9vVOWAyLBAAxSF1yiXlVWa4N9iOtuLI7Ue6Vf4VdW2oNy
Y9TF/sbIDlW8brPfNCZ9FtIxu5ydqLBlZrye83wPzBXsLxBUbe28pUyfqDYiMaj6ZyOhNA84FNCU
vLhRdZ6NXbBCwaJIAMovlOQJ5YKZ3pomDEslza5Z9vHicn5CMkpNvL45WMXJWw9rtZHAX/iNghso
6DRNo36YiTE+Jk9kusDxTbYo1jgj6RKZSh/BocLhae5PdoLoeosvLFWrKW9fQRBP5c+DwRAepNRg
72FYsaUT4bogKiJHUyK/I0bvGfFV/pp85CzXu2hBC2Xp09OfXtWTYw1bcALeoLkzE+u7vKnYqO6X
245l7k+RIPn2FhrilYxx9SP7qNkNxt4GniSrlkXR54bMLrpfeRucTsfC9zSGN22Nq9RhWunNZfdk
bFG+RJFh0GFRGdZRFBOT0W7SukxKcNraCh4/gTjfgCDEtkKzXdxG5OqTWq9FfSTij/fKHQOGcvRS
jxA+hKP6zFzVqEeFahr/4hTChMjB5SHNrZpEZNYORLHoSCE5Qxmml9CJ2+lO/lBoe+LqMKMLuehZ
2ykfRF05VHbhajkTlUTpfeTYxUk6wPWt3CvHFOqGcuAQYgd0ADFuwYM3xxwF05ZgnzjWOPsgxUaP
98bsTp4afHP2Mrj4IKYO0KsSlWwMswyTesTZaOErzlj0Vgs5Q0az308I1IiDgRQpX8J8Mzf6GBdv
5D0g5hYZPARN/XRcWJ58BHvqDAo/NxMHTNt9H1qmPK0TDcVqXRx/gyv7MLcr8Qz37gTeInEXuPSg
ok/jAaQirCcRe2+Za3SuQ/L5ly5xNc6CyEUap/CubmOURBvXLvAVarcXA0e3Jk2Td9oSADGpz+YK
HWBeACUu6+VtE5RXz93ybB6QktfuVkCbp/cI6PHVzSOrrUrCblHbzzzr8XBHTDtU5C3uOznG2D7B
jZDcVegyWdcu4mTUQa3XBUDxMe5UtAT1zZGUuI5G9H74NwhcY9yst0JsD9vDkGqKzZnca+1dJ17g
qWtk8MT1qdK8iehyhnDLdZpIN5sdk/jR0zLmjJM7YfNbcM1TCyHhdqA+tOshJzOSqcCY+ZA8H6ok
z2dy4k5ZrEYqC4OEqa7ypUoreipN7aAnbm5gZ1XXxnzosuF9R9UfI+5B8W14R4KoKmbAiKCebOnY
ehH0DcVJLBTcTKMo+qEBlZkJAsCFwPT6JBOuU0xagWUni9+aUPebMlTu2E8tO3b3lm4ZJzbuoYtQ
FIgFKXoX6sni+DFOHo2k7V+SyWZBP3ZpoEBvEoFw2s+pu9CHRlEbMAg4ZY0dHaTOpMM82ygT5wCQ
TlKv6/sPRUbc7PdAonBmf4UtZ7En69GZsc4YKmByu5lLv9xysK1zmC15BmmZNbaDITBbDO5Ce3/c
2r5cpm+7mWR/5u+iHwoTRfnElvVdY9rkRIfGK0QKwXzAqgW+Fzl59o3a8JCRKNwN5ZrTwL7tG1V1
5PcppoB2QM/4ocknmclZs33RzKTtntZ/ZZJRBndEVgg/5bXAi8DQT5yhoyasZZpWj9ez3/EZk8pd
Zrcs0YNNyfUZG9qkblGVjFoh5w3mHshCARN58Rh/2eGtNwQOXDHJa1gqB6Pe7mWeTBYnB4x/Xhok
KK4MsFEXn3LENqdgviQ1YNxb+qTbEhwcfcu+jl4jlBbdu5Squbwwg463e8ltG4Ug+vJHuC4ujAhA
0NF/gkpldrrfJYK9BSRMLMMn180Y9VlDGwJFGPJ5/68W5xTpH4z1X1qnQw0J75S1EF+wCgXNlXz2
wQxO70rcUwvqYxw2rIHEvaE9EJ5Nyt08xLWCqS0QBAZLgkhmNLctzidPVspXn1bX6HogYV2yww6+
egwAAt4tZ31bF58OXC5nNZLLFk24qkMQs4yRbo0QzJRCRKyuSqYL1X5tjVEzabMO2JW+deWqfGq5
4IXxdUsfk7obBt+FTdHVcpqWTBG9Y6sXGtoQUxSwuD48jn2KOtv1N0Y4EFlBAeFV+psq8YB2look
16dgDmPEoN2NFZrM41ma1q9QK3kMiPi2GtWeMdqHvB+ckWtjURVErYBSPhymkbPp+yNVQe6nQKFH
VqnsHn0wIgWWT9vHhIbnymGuj7O6+B4PDbhZG1Dg7Zx2Gq8mqDMpos/mX8zuvQ1+jQfHVDEAzYGd
6MAn1j6rKqp1n5pV0QyxXVFM4pnBS3+AHf+/cOYj6vKvk3OD1zRbKiNgLUBOurEB/3v0+NRwfmmr
pygauqLzJ47EKgXPsmJGhqnVTvdppmnmbMjTfwyIKvOOI5BVSS5IQoAS50uC6SZ4X68cpGmE8lzl
Bkc6NX5xYVxBidI+1C/xgh3cPWuKTX3x3kmGDE1xQyIXpXHYhO9D/3kA95pJYs9z1ZAI3u3SpCpo
DMZVRdZ7idZsc1VMwgnTOcmQacKm5PxXkEGjhr55g8utRNiihiMdGFBSK8p1xiPQ6i/6rk/KxxxX
FldaR7m8tzR4qxDtr6fRWUNpVVdoENiKVHuewtyDAw1kvoykEOw3sEbKz41m1ZGpur6kD13B6nvD
C+jxUN3tyw2bysu/s1H7OwqHQUuakzrvKhnSXHvmV4ElkrUB8aHAgcNaMlBi9CGxaxgQa0oEwHZf
27/O0/jYAl6eLj9bqXeihUw+ZqneXrQiVtYwxUUPFnckMYNZbJt1SR1ouqcFORr/FJNm1eN7JQLP
xaWEC0S95pCtMPcEu6oA76nc5sndUEpieli5T/47isr8LQGG41B80sAtOy+ONl1zBxdiFj17oxLq
NseNzrtC9jwXE+aY/7ysQon0Ar6B1IX06bPFbeNA2O7jnscLqRIB0CNOBlwLqTcT+OI3QT3zFaMl
eYebdw+AKjl7SuMaR2+1HwwgI/hGdC9JXEczop6p6V7uLEM8vGjuBO/NU0HvL7B86YtfQqpXaImv
1BxRLEVUV3PqZoevn7ihkpNxgPhyZE6fzfynGFwVRC67IK5SRO4cJoO4tGTr5ko6XdM0ldgGLNFB
eyA4TWAfuG636p7/Ks9h7I2Pl1iDBRbcyafs8U33dD7SGtPwvhu/i3m7ts4uaAjMchq1fOQW7GAl
BwuBtpjY+t4+qqffa/jVEMdq2TnvUthTOGgacno6VnDFk3/PHNje0Mca7ix+CVwpBbrUUUWWcExD
Un9X6wuuD+nezj1nkXiFUwvSX1GEeFX1PUppAaJGgkuWGBFC4OxieKNXFUomQJQpuzDFGm+xtPH/
SWXqmfrgxoTNCeKVMTM4jDzIJlJWrHVUnsEbXKatdEgslt9rWQBRL0OPF1T0n+MSvzRNVKLltbB3
b7W98prMZT9euKZ8RSwfB2AeR8MKmpp/3/a47V7zAhPOrerG7y+bRbDAO30zveFTdppxQG2fbPPG
ti1QxTXzliUnqik9or29Y6YjBlWs+P70f3gU+FlOqhwWz+zqvkWTueOHSJg1eTtr4EnBLXgr5zSY
fvia7Ne0kBdkekvoZdlzODipRE7t/ios8h0TVO5fGc1Fp+rOcGngMIabNOdcN4+dllnJd9A7kipw
wzx2/3VaKM7W8IUIol4vheyqoNR50qHb28Y1QyBGK8P2FoHyRgotAWhRpmGfMZ1gouRLbRzOnnFl
2Rq5YP5iLQMV7lbdzk3gQAlStdX50Imr365H+1SRBjYL0qZMhdcP1f5mq3G/W0ALzJ5kUkjRDJps
WjH2mSq7MwpFs8yhVzi1p3czXE+FfJZYcaY0dZlYSIQlWGC9LgFhgBoi+KJIrO75rNjDktJ+9a8P
1TtUWSBS0r79d/cC3uJb4Mpyvo5XHwcxudqZ4LzOC6NyMW9Gm9TEeo+mP5RRy9NcVWxUvwq13PMY
16svUSzkU0xojEhMTeQu4tdc78vGQUxzFILtcz8vPUiV0L6ksENWa+YFYC2rLEAhKCRnrPuRKUxP
dvEI+NpFum/QjuWo/lLU1+UBlK34SNw4UV6mh6OMEO35cXHgtfzk9YLC53X629TXavxe/jmKG9K5
0GfHJQOrU4++EfOc9m1ad9LnDhX2OJtMdETZMQ/+UHn94jpIvE2VUgb/c9taKgmzWKMq6xhKKAGz
tbvFKvpw/OMXiPfvEAyh48UdEPQiS3lhVCoAaQd+oOQRM4Wv9QxtdpeKPO2WnpwywpP9FbmSxOXp
1F4AyynFtNbGYt2YMdJeaELTKD7UKwaon363fRHhRxsbw00k6Sin5jmNh9caYIeZ7p+/aKzamULg
3xJUnwFiUzIxxiQAU1y4YCz+68YC3Mtj2lijeuYupLYa7vQlj5HlRykGJ65v7yWJZURNvtwx/xnI
EuGGp69vWGEdv3SkMmjr/+IUBfVN32RJuYfbJND6kH/raxoRglxz+GLiX1e7g4mEX/U4n7qQMj29
BGx9lpdjp+M43tF8jyez5rTeGrsLu+NTCLppQYtX5k9gN2uODlzOQ2d7K/RcTsUCPMAc4T31tbU1
XVFFvFt2wL5DbVWgXojE7/0zU/k20ZDIAYYDMN4qSO0xFsdhOLv5N/VNjHTL+uTNjGiW9f2NJya3
GNOds93x4zY+Mzj3yTJRBr6J0zuPxtCYbv2CxjfrHf1+BjoXUrodko4peAom8YDxI25BagAzr3c7
6AcGIWFTmP4UKyHG/RqAKbhlrd6op3Ma8Zx2oTZ4tUtEEWdBVNup00yZrDQeI9bIF4KW0iXE8Q8j
Laj1w934VUZIOFXevmMroGU3w6WrwSWC179yzUiWGokLBbdfYNReJPdn895SL7cTRwzWaqpbkKa8
CgMSrg/2VrjjEECm6LQchUcdQu0JcZs5GkBIinw9t6CaNfVzFKL9Ds6Jgi68H0ZbS5Z6jvsoSnAM
vFv69zY9dP9PsiB2La4AA3qk/GzU5UTRTRKF/842rC+eYFuQ5hXTVtKW31hA9RcRD2bv9Zu9U2Lq
QmEfBj+no6PYSCWyuFixp7rVkzj66bvrC3JVz4496flJ/mqbMDZ62vOraCamNRQOESIgd7tPX+xf
JlDs4AOItAhMatlnCWSy8Z/Jt1bb1+Gn1pRtl5dwgJenQXWTybtztceatMN/RMNXAwLBF5fpsoW8
GYcHGWocpfFQcyEzuh9I9CoB0u/iqAP+KFoTf8yeJE9KkZQcpBzag4cQ8kyMMvcotUvD1kqpBBgx
/WnznRdjjIRPtXadG3KfOq3MLBqZcZ7WjwKH/rSmdPTsFyXZQ7PrU9gBf40SR2iSqIs4IgX9xIs1
6yG110+W863KSYbbXSQvyjg7MJolpyDIXsLVIw06bf5cgEX9LQGaHiNR7Vb5L6grb2bJSIaiRukQ
P/mNbKsaadMJzmfRuwOPWE47xaW1qNSGxBeLamy0x2yoZ9fsFM+jJ7dgs6Qv7euTbFoDhQ6ZN1W0
GvcULmCtoVTMEczpJGfQ745dzQy1kxLCJ3VXY+V0/tPH/LUTe8fiILMIxrZICjft0q/LGZrxNqca
zPmD2NiFe722LHaxtAXDIYi3M70atc+0+rARY3n+SiMPmZl0h+3Zu/kXy5ZTnwSG/BFXNgekO+dq
XR5NJqr6iyWJtKDZxX+unbUaGECpJhxdTdyYEY3nbQ+VfHPLwm5RujI1VWk0thIK+Iis+vP4EhrK
bhj2kVjQ28LbXTG/Ut+2SNJ+3ySpll+vve5SiGaWEjGG1+35s4jRxVU/nuqg/c+NcG6bbaHTwFAH
uB4M6sQp8silHb/QRxHidbLrQvcCSUA1A4fUPhk4xL1s7A/IhxeUw+IPUz1TpZ4SujavtMRMpjhN
DM52GcdgfWBMqVRgga63Wm9CPRW28lvLnUa1lOF4ZkI7oYefYuFrzBpSqP0JJPVX05zOsCM/JLdN
tO0mWAmv1TIhUIz5pIUjlKCyKRpr9yHd1SnHMhlSYjl7A+IWX9DVxxAQQM495FHUeNJCcXCSpIFC
n4FioCUN6eUmiF+c6AgMjp7IC6+VePVl2U/VGbEvAw6JLw5MjLT0dyjm/DwajEJGUJCpug5XoWtZ
UjdV4yGpQ9W7l4qgwRSGcoiOaNU7REokd6Mto4I7TVxgkYaEh0y/fYa4Y+nhklDUg0WgIwFIDpXc
MvXfIuNQ3N2DdKZC/fyOqkCLv7PzxOCr34cUxKc1LX1rFoxppY4kvkUTeWeWM4lC8CpHhV9sTP4w
j8xlWxgnO03cNe/anA1+oVhj3Olyzb8Ai5QygHLFkBCIsvFJcz5ySxhKJ/ZT5PvehENSq8leJ3sJ
xmzhhbzB0YVDlCrH42q1Bliwv8Fuo+zRe+jecoRw4n4qcA0vGCR31C0dIyGE2ckmQpQIIRL8m1Eb
12ihYh3ya8Y8tA10Q0r1k5EB+TsWM8/T1de1tqcrtYDpEV/1JCbUnt3mAAnyDDlF2rBHLSNbjTfH
mYYxrDjDEIE7SDLTUuPko6k9kKyZ4lb1WBrQIVTVMlNc6a1Ll79gmvNQ4VUbcdiCqN2Jx/BT6iGG
f8HxvYrGFEPxBpqsPru0j70upp6MMBNlNioZZ0AiEG9ZGIbOpcT955wnvIW9Yo0bmmnfV2Ef1FdX
DNsFlmY6+CVTSROUdW7VKUSlaB6uTrlqk/D6fblHFxtJBKwa8qmSAnhI1TefhMvDT8FuYIOokjtT
2a2Lp7Ah27mwiGnZbDFfC6+8p5qn7eL4l1Q5GPlcXN0lEOXwZCIHjB99afQ1sDqKUgvJTLf2bJZD
adyZiq4DoQN5GQdJEpyT326talJonC+bEoPNKlV3mkvgWCGYCT8POG4sCDu44tbF9vnJh9Zlj5C8
HVukK9D+zgboebAQChkekC4l0Zg7Tn5yUuYrwUlRJOycxKZxZRk1CrpO88BccrCTLbSn35dJw1PK
Lrdwok4vx837YWIl81BH6Hg60u9u/NBw2m3RKavIIylzsesBokQRKqoW0ro4rzfU10ez6sp8mIUK
Rpx7tGG67Of8jePIDAkLTzjlrlN/1WN+mB+tW9fid1WUbXi6WC5aRxG4VEG2Rgy6yXj2MfO3HqJC
Ju/819wWASNZyHv4WoC/Nv1WemhMT6fq1M168jmMy2kAERKBGCYw2B0Isjk92T+oZsT2jFHlqcFC
BuekpojepWfrqTaqP+rKgRaxTaFf1sPEujVJDewhcE5cIymWCHYuV4/CfcyeTvz1dFVBMe948Ww3
Zdh++SDpRUBhUQ7WHkkriArBU/in6e9grv6JlkvRMfQweOVM8GUC7NMafc4Vr8/t5seA3Cmn8JR6
vdkQMKYo/KlQiuWCjydrh2piD60Kb8UftI6aa7DRT9C9CujNFoEkR7jjxAHuxx/ySDFHcGdPXz9l
VXQo0qrsHjsp6uvggIk9jnKMh0snaudacBTp0WglfTJFrb7la1NjLd4XpifQ1xBApEnQ2BGSJBiM
W6KpQNDp+ixMf2cyvhzdjyrFTFPcFwQG5pPFghWwSMQ8EFiV/HXIDW7Qt+Sc4cRNNRiP9xdexWc2
Gz/UiMl6gzeU3ypb4/iZXXmObsiqROdPGbn4Ra/JChFfbraHQJhm1U/S3WvvLLlgZ7oeo9nO+Lms
IVh18V55H9IQQKCYBOXAGSq7lfxfPAoa26FrVhN5nKO1E4MQaB31U5npWqUqKuGQJ3FNBYk8zRrA
ksWgNKmeyQnjiNjlBOpOSIPk4vFY5aOoufb42GkidKon/tiPW1hlcK9FkSwmWgUPtF3iIp8AAG1m
RC8YTT3azjKEn0W+yi7IRHSqGZBF6vEeb3GlSAPctxayaXaQ6HU0hc3jtgZnoUhQsNDNmbrcfO51
UYVJ4r5XlZiXzsSfVoNLGJJ57TayEQYvgQWXzGXzJ55X/aX9hqTANCogh26ALKp4xEGjqnGb7cZL
auMhSKKYSMbU2jjUClceC/vUO1E75tH7mPR8YpvxqR1Xj1i6sr3h/UTWF/AT1vb2pNC7DLduP2xm
f+WESWesplGnVk7vwqBMbi/XvhylWTZRM3aYFkCjCQRJq+goKZL4zTA8u6mqE44E5GSi8dqq0aFA
JcO/r1Pq52f8/ldlB6UW57SQGXMq7nF8CfZESDbM47rmioB2k2qIT3iYrRVknO7XcizD4C2s5UAD
FuRyeb44ZodozHwq5X6Me+HzDIETDm6DH/RJBcjmoE653s83EMIasV1K9suOXShoCJMBE21vgbgz
sOQd6THusR4Y6Jms0cmughtyn4Nuvn1V7WUQCQm92vcLzdDi6wwlvII7l4fCmtejWLdLfsFcT1e3
T/5kbl0yT++rDKFhgNNFQeQ9L8nWgkmY4Pl3Kuhn/NXdfqCG2pfL6HuY97aUQUMFM5g8CTTPoPXK
OYHMWqcV98bFAis8XcuJeY+DiypU7oTI+sXBKMufj2/4qmWNBnshHKsOeOnShTAs9h42d8nt0qRI
lBlp6RXyRTFAxloArD5w2pbJ+Oylb42y6M854NUI1WWarcdRPBnpDyKaCBGRgNu+N/jx6UVsYXg/
QYLDcZmxiZ5VAtPVma+qEopmQ4pa7Zz3cANeOeJ+S/NpELPy6NSbqbOH9NsGhN8X92mdOo61tCNv
cZfNK1rv2TsOeouxt2d8gSzVPKd9hwH95O3CaPu2JxeEGaphzeaiNHKzOcM1nSVu7+xbXH8a4XtY
RD6CAI6XScmHxVQ6oWzzMaFjOVSWxmMGC+sIiim0CajOxtBDClm/9WhMVjNJj8RVSEOgMqPdwQf2
pMVybealWsCkG4FrNqwimTCXpvNWJAJfkkEBAsVYmJahQcFUy5nqrb5AP23t77g5Ezm5tVlQHPn+
nFDC5gntHpBb3ykefq5lzz1AF4JLv2fYm3sq+8sGIV8ZArEjR3Vl5jQMHI0/FKz23wIH2UIOs3iX
fw2EzgdAqZTL1Yt3jClKog4g8HJPnQljlrUqJHuhWaFdXgqzYVHde6YhX/wdx/keEmAM4xkoYpUn
KrfJ0ZNQ2633PZmaHqFdgkVYSVwGghViR9WkyaUagDClN5q+hFy31Mhoh5fdC8eBmDMztj7rO5OK
dtrWIAuT1cagQC8DXNuDWMoKS7AxuPwZER5iAfT5XLGj6W/yssPmMP9+db7W/qGHfgKILN0NooMw
ZNu5upjRPfPNJ/cBCSGadVycYubYSaKr6sw1+fENhYeEF5Ipw16dqJdEYs1L/qwOzHxcXswz63U/
rscTbTh5RLbCV3r9YjskQgV0opmnRsuMIggLvyD3lvC4rk9Jw9U4T6tyc4zWe8tsMYS4zwHjt0i6
Ut4bdfRk/YA9ovdMUx9cAA7bSHSC56S3cf3TiKFEs6qTox0yHOtLRt5xaZ5iMxtRx759UJWZc/qQ
/H34y/af7d+7RAsGXUjOgK2PIv3IoEVwAYqSh/mw6bwf1jOES9aFG6GbC3yzlfcdvWP8H2RLBw5s
HYxVP3v40zYQGktTtYfN3/tyISAj+B0+yslFLMthiISZZsN7mcKXs7Ok5F31iL3ewz0Yob/YqyW0
hr1+dhcu6lBpXsdF9P4zcHOGO9/gSXXY+YxK4VRZT9uHwDbSTZwLpu4Y7jWINCdIfWVbpQS5MCd0
5xAdYwjra+kIm/PGnovSsXDEALojGz71ICyTVWEw1YlCOV7q/DjPXWZVr0K59H79BwLjkaN7bquT
A6wvWOXSB1bCiehrdnC69QRNZ+xaG/lDBgTYAqmrnmSGlV5uJ4JyDYMxTdbnNolnQ1H7RBfrvYrM
e5Qs40gYYWyC4bDfWO6J/BxmL5gjzae+0bQU8aaX3Tqi7QdeubQ1f94VlN49OWgnAzDErWVsd9K/
Fq0uGPrYJDklkAO1MAvl70/800wmO9LTvt99q3hxyjHsRuvMCYWvZjbX5Do8dMltQdBoOwsrfvcB
3dUSA4QuyxRnah326/KVaE1iN/5KNXqKxVtrltsMp7ZcYskrE2VOLWZazmGDIxGH/2smOHQGwIXS
TiFSz8+BwWnbYuWGMilbRCVqxViNRdQqbol+P9IyRw7uTg0TlLkpx2PYP5vMZle1htsOUR1o7oA1
MhXMriLoL0YaTjQnleMHhU8fPDeAmub1swDMUs31LX1Y1Ekhhu8qS6i4Fvw7mMnZjbUSwcHmXwHp
BYLI5Sr0dVc5Kj4vdUiA4MrlQnIay8jJ5/Adc9iH8nkUZ8J9Cat5XmNVgDZ8d1/+fdyN44qzlKin
rKGHeYhrmZ7lrkBQiKQTMji7R+PfRWP3WwQ71RjjwAHbkt/fSYitlndNFyBqS32nZr4jXxtj2Iz5
sz7SXRX5CcCOmhjC5+AcCe6mjNwDYaIekXQctWKOev97KgzjM6RR1iBc8sxf4nVgFy5kLeq0nD5r
hzIPbgpJQyVP61P4305EfzifDN/fxVjWtaSy0o1w57QKQHqisZy40mr11SZN2lI6VTmb+g8qbIFs
6Er83ZfL+Ko//JuPyCkBaAXBKqD3zeZsLY2IBlGgxykv0S+HurLpAD1vMEh/kZhXMlTvXQmUQDwI
t4NUDzIj72QBOtU28grIi3mNV1FzO8JNIoghpQA/Zwhq/C/rXrfKaRgIUgHlh2B8bkKUTnT31u6C
2X4nG3DMAurJA+mUD1xh74D8Gk1Zv0zammTRp4UYywvKjqQ/bkHPxxJM/y4rT6asZctmyiVEhZdz
h+K6zwpcJzgOE3LiMnp+oncS38PhU17uADGOY4b1wsV8PnRnPuvIk48mk4YcWXsr68190d7Vamgw
XEIr5EvlyuaolzX5UydosZymcKTdTUqYpn5D6mGm1Krj0T0A+zamSqk/hdlHGKlkxmFjxJ5ZUf9a
7N30rFSKCPcS0Nov4Uku/R+RUNkJybQlX2m8UqOsmgwuygKJb3+LPvHIUmSMoEslPAvUIdxs4fED
RkXmpK40b2dBnEGQqu9HgVwLClYFyyrE+1PVcusyPie6jHAxVjeci0yoWJYh60yQWVRlM7F9HmPH
mzC/Lag0POAZVS6ifyOMTZOQ3j+zPpfIQIoxbsx8ddXBVU/XzmCHp2DVwL/RmKRzL0wHRchlfeoY
/U2waI/zoY/o5HyKmXyzmEBbz2JADel/5R+MjLoVED/jHpTIf37JKeSnx7wWg5jVKDc4Y9aZBu8M
AFutqGUZ4cSBHzx0amh9EFzfXxIruHeW3VyFpLKvGI/IZLONe3LLT5Yy+on+wD6Ma/TMCRrOfeWB
DGB7YW4+0nxzmoogAClta1zGBrQYguE0JGPyRcBlucMwkkMegtJ1eaJZK2BVWl6LsiZrMt6aiDYE
Ab9wBx2/oUcdg6zlQ8l6q9/grxZnole3qskQL+EL24gQtnWmEOrQNrEJq9ObYNJxbC8iZMdw/W/M
3bCPOe2t3ymK8WtV+1rm+7T0lK3d+6HIEauxBVoIOaKUQn2sPqVwsI3s8WBYJI6U6UVeooAAqIWj
c2qVqostCoIV2O7NAJevkjQjKV5TOltYDhaEY521M3D3ZlJDB3Fm2O/UosjmwNawfWSrcRJhiUcz
F+FSaOZNQ76ejPcZc9USUcGkXxqEAGEn4XTSW2aU7LALBpXcWDJhdsaFUvQqqEThBhWqra+HStRY
KJn81q4Qg56ttYCmKK/V3k/B0si8pl7+bUra9LH0YXKq1djzsqh72XDrYEzRzIbwJdIdTig/ZllZ
I88uYZTXIU2tOY57vhJfhc2r9Dq+m6sVSv8+CQHpISHqAwQkTJDJJtsIC21P90/YYec7y79cPfks
i+2hqEbRwnCkzXkr7pOOBnWu8KnEYr2iEDX+8IReB9ukPniNMqCocStOVk8E6tzooquDnNhCQB3U
woZRyGt9q7p/FqqnBKHVRwtK4klug3F8xdmZol+HXBU3glCCGRB1IUzWR8YZs/gpAdDeAGj8NouT
/fs+KuKodT3GRohb6YlfNMwwzT4BS1G3Iv16YMnWl7lfF4dZMa1NmxaEWBdeJrH9cBx/KxCQYAtF
vUujjgjpWgVCmPfW9IQ1Ssl93k4QhhdVJ37To0sfRCjT/fK2qo2BuPE01M4w37jYBXz9BJvevvaw
HgG/Fy9LRMAUiQiZyVrdP6LB3H6+H+d9iDfz1F4PX3NVA49ucM+0Oqp5HTNmUGgMjwMnI98ixeqU
hktr7q6xSEdlW+Zu9gYNSlVUJHkdC2jyTxQdY+GqTrwVkl5R/6HaGJjfPYA1VS0Inx85NCzFuw3f
8TEqfmE5kFE4dKTGa7l08T/+6UBgVzCN7dLQrU4a+UUsO/ZHW2qE13Nap2RSKPdaNxfyXcA0PMLo
jfy0ua1PzMSw4Y3msINFFr66Rp7N2z2BbO2WYTR7eFX3b2fRCiDZxEe8DdD1ar6+jK4MPHe2euDI
7/xsz/FVDFIsmmJ8OOl2mIjnmWfa/fD/BJ83rIg7l6b9kOn2oRlYBYFZxSoGUsztuFq9PZahXFPj
xVM8SMxeRpQBcYZzqXuTNZQVD3RAd6gqFQqNJWzA7DMEdJ5w6kuLvf6cUEm1ycik4tK+gDwsjTmI
F8ODHj77foVzIwwPjU5VqFiK27SSYGQURuQzoncWN8RsV5xdnHtBwMJnOD+OdA4m43/N4+h0A3rt
g0yYNoCcGOtV/IcFIIwWL4HCKNlPnOn5qhQRrpGK0owIabrY2ZELgkKGhvADc0pj727YKXAlZvpk
NAhGMPmARhUYZk5pcl0FwH355aQF5y722VX9TNlL+A+B1N3a3yGHEzJm1aB6crjPp59+oMX2JGUk
XFWwT8wwRpovVgdFRNxigaxNsqMJSNyt+fX+hEpnveHwyUkQPMMkzqaz/c8aY/L0WTthE9z3En8b
v4fj56s5WLJRJpk2bAmy30zAxTbwJxI2+UqhUxsQLEur45enZWPGfGhNzHsVqd6rPM0+0JTw9cYm
8ln2JCSeszwn/0qQYJgrrTOLt4n66SCBGGBfSGeBE40BE6f0+tK9Jo0uwS6fiSwA5biEuDkWEG4e
NsLvKpevUrez2KI3rejagiAjpYzKUUUYDURDN2K/74SD/M5zef57s+YB2ZjiUWpyizRfoW0uMX5j
8yv7DwZG290YcZs4toSV1pJ7+ki18cwFzSop+diXaGsTWQ29dFYW4y6Gsozb8vh3loywcU8Vulvf
SKqCK+hEolEu9v3wV2mOO32pMJ+XOY7kWrve3+hNALmOxqroHmZZDlr1PN0b26PMVN6kuE9lArDK
08+MqZapBuHTSxNz3NoAfyWRiewhc0dyxUweS2HwbWfkB2Y6NXHtxh0Hrb2rTvvqNSOtIHKvNNWJ
PJfl13eOESi/FYjmUa530U/WC/LhV24wrr1RsIoVAOasgrMyHqLHFhU4G8K3s2mb86LeTmZgbxun
3Uk5K1o8MOkieLssgN5VigWK5q2bA42s0iZhpDrbTyD1Fk4GNYvPX6ligcYfrY/aEeoqs+f0OoMo
HRQ5eJSy/JvwYW266TSc1AIAMa/gahHxo8i6uTc8aQd/lyyFtkGueKoiKeGVv4ZWZ/w4QpPCr+Qe
DVELj44tLDDpO1JuQQ8mmYnImgvPwh7WC/C0bRZ66ol5V6j1SgtpAqa21mjZ9jUpTz+FgXPr96Xu
wZjxxCo5zXwzH2O9DvNcZpwHoWoB+JPv+xnq2Zk7awGRTfiRUzozhCOKF2AZfiKMWMhedQQIxfQ9
Gf1bajFgQyyNbie6rjHCvw+nEbHWq5kwzrslYXz4Fdsh+m91GZbH4d1Ku6nwvfUqPi0GMRaS/M00
FsByMt/ZhxH1g5fBMRCIQ7GrLlMECbrCNiV9o53bmdHQSoIpHrLU8bjhU8N0D8HCV/iLNlQwNn4P
iUirrIxGQFvS4D0HPEsClMdRYshmQtdxeJuZaq0b9DPHBu7MXx9EDWd4hOXpmYJGYGKZlhx6ckCy
cN1KIGuPv1dSOmtLDbvTbO0H2Ci6L6E/VFgWTQYFO+CDR39p5o6p4TZX+ABebJavyIQ5+FgXZKeR
CuOGrw7r1Uyal2F2W3t8eSbJsU5f/8EOEAa9s8nByZgGFkfjzW2SYVnUf94HcVM9f9XtWoOAhazp
Lrm1eVlhABCm0wLHx9Y4jPshD62iRENhVDdZR4t2y0kMM8MyWuehUQPuSRLOZb+g0aspFm3pz7gG
Dfe8KH0LZQInY80Kf2SVPVO/Z9uZsEgBhfSIuK5tpPC1fJpLdGH8GeXQsrPjRreIaWLkqVU+uSap
Ugn5Qc6kNx8fM0Gn0wNDCSZ6M7hXJRWVZihfMQYbB/OxB6xG4PrrzjAXmdw4gsgT5LxYCC0k4hYu
Y0g70xQw4M1HZk9RbjH2CPXmOh143HFwtWt2v2sFQgSNHhWiB03BQ7CsM0TZVD8j1CnIZ5kvimJx
cBJEPpVwW28XqXF5JE7eXQIIuyJ+pbT9Fld/J/rlL4PCJVVslMZSILJshPauR7R36vmEjt3l6/zy
O7Sntzz78nhzoEFDVZ24NERfmkVL0Q9nb0/N1VjOSmGWXsQUgbcBZtdQKvi3N+5CzZclDjQmikyu
vRxgrf1NaPO03YVRxnMwn6NcASBHM+91tIvBvpaZNUgtqzGp2nFxIIfdaP4PxcvYdjbZ+meQRmrA
gHcXnueB/O+I8MhNcKPw7qCJHvch5YzDYtUq7LG1tgLjHAXwjUQD3gfYm/FYHxj5fiuUeOWM3cJY
i7C5BzVcetHqqTldXV3FsHw/U6KhdjIMaJW64+RcLChUuG/Csea8uoyIz9I/oEJmWP1z7AFwOfi4
zUf//KrIxD7bydl7QxTR3Yo87YpvY/wUutI53SR1v+lMZwwu8re3RX3aUJOH6MpljSdhi0gr1f9H
tOqPBJKZTcNWeF0ITO0H1UEwEuKh7JP+99v0Y/CxTLwGhFmUPG44GpF4PEcAkZPZFmGQJxZ2gvvQ
a+s9XQcNHl+AmrwGvlBi7gmmio34acgz9P+qGdquYNKoespgCGP8svl8aIZ2Nrgx2jtEXmpf1pd4
M2l93H0feSI3qeVqCxZzSMtEdBegEn4wewfT97C3mBTYSS+HB+kPl0BLy0cAWNdu3D/vGRZqcfss
qu/KsScjpMl/LMpzxauyQKUxKz1ls0IxMxIrWpXBGRQivdMGg+YhfjybabIXNVkXBITJcjbBJAfq
wPwBg/n/+CNbgynpcHBK8nKWD906xXeMWwx0QKs8dA6gOD8VdhSeUqpGSoIpehFQkWrHMBqrXdzj
bG4pVMh+mpswIABwmTLfW/GXj6nmOSjI+6Krgth4NE4M8SivHhk15sfsDnF1zEse01QVoMoDAjcT
q4P62jm8SYzaNCcKZIrT7ozHjpp+RqffKN3Cr76JfYilpD1+gngu1xFjD/6xqfFe4LyLNkwairLj
faly/giQPl/WmsX1K4jpzCc8+SIV9OUmIdU+PFejZOAUfWifKAXC5FhEubI7XPYdnr/Ff2UPkTtg
BEPlcR/dUy1CksBXllrSuCKPV+HnWtU8IOlP2XriZSensou4ajgC7+N5YzaVv6m+kUBwfs38h7Ab
WYGZxmjU5tv8Htz+pE5S5jik+BrCSMDqFiTI3+3yiqm6hei4ENtrKhXGDyLFV3WzCG277QkPKAJv
PHxygBUATRCy3ULJ6B1UBU6RQuaq+PYwf9dH3YCo+v34LH7t2VVZFrcA8MzdayMzqUraRVN9yYK/
Z7WbaatiEOBXp9A/L21sSdVewyy/S+DtBncnt0vTzrauizvjZ81MBuTqvCL2+hbMCUH6vkjugMcw
bUySetjTiDxFg1qemejkr6h/LFJAoLghnKcsOUFp/kY2TDV1EqnMTCFFPWaTl63r+mD69sqHwJvl
Tx0VfTk2/5nSFnde332kHRvO94MZ0QkVzsLkUZK1q7EW3TQfexOKxV2npjfe8EgJaIAqTwfVBepK
VNKPGeO7wtcU77yCrRklKqHofyEzeXSCxKHm+pST62tlCunrQczQB+n9QJt6pGJB10rl/AmbtmOY
EIA31pEVZcCxgAiOU5hrN0a61c76f1vrCGlQzbmf0Fz5D30Fpjv7oiFSuW5qLC6v1UWUseRIw6nz
CndCZuQrryJBrzCA0FlggwVG5HHAATMUk0aThHi/VvRjoP/rHI4tit6uEmFdnmQB5JSAv6XiVPHk
v6yWgnX+r8fjBHSHnCOYJZ0ABkit49v8/ib0qycf+Sezwkh1zJGBMUrl09waHyNBZ3lnio1T6wuk
hpQq7xEdukSVeeiAttZ2IcBc1aJUya9zNJTtHKAgcjAFtZas5s0xBUK8sp3DeBt501lLqg7v31WU
YJNi19cFerY1tdOl/Mli0DQb+e8wRpArltR9j20WnHeGBcgrZcm7ep8x9WlJZPIMVTOiSJN112re
NJQPJlzvlQ2VfFBnIkT5+q8A78exAaJAdOHDQVMdYbTSBw/EcH9aV0C/XPnALKAYm7ed/vsuNsbX
dTMjcL4PK/V8pNaBhn5IdT5I+vOlFj3kCFkX7r9Imb7PDTAUuW7ri6RFjVfDC6ZW39XfB9G6+1/h
kW9fz/JDz6b86UnRfRP6hB2FnVBtiEQyrRtXrRkYDmtuRzL+WqamHiH1bVUpsnyJwDlb16ba+R2i
ZYLQ0YLmKnPT2U0bmIwdAT/ahf253HCXpDDsiiBydKhfyLxlpqU8v10A7SUCwVGyxiGwBYM0IaD2
DeouK0a4PPn2LHi5+TLBCuvzO4qfENA24a0eABPm47kbJd9Vw09GjhJ824cS+GXxt3UXeKkjYw7y
H+or1bbIjvjhXy9Ku+PcQBUNRAlnSZWvp18IUu/KIbRgp0OlQF4FQbKwmqHRCxmA+1mOxAQ9NTG0
c3v4PT7zgfOq3y1XncVRltp7LawzyZ28Pd6YPPKazi8RAxeKjAxOtthHKm8TZKYSQOVv8i6XlnFN
43PxoIILkAXa95ceaHcKoQmiutcG3kXo2M+RB/SLpcHSQ/2nfyb2r+7kQfV8FTw6fEtGsqAxOnmX
t4Him+SaHmGZU+lTb2j7IHmraxoSDiMCw4G8YFRFQpVk8C5Mr4hNvnnUZPAqNu+y9pp77PUvjxm5
HEn4fBz0mGLKXyzaYbf8P807xI11JqgjmHwqnaTFgxiUxzcca8DVC/7Ylm6e5gHpW1k3GVej5IzJ
mMjR3YJkaeB8jp+E9LaSdDR2aEoyZJnpOLIpy0MxOOBvc4YchtKstPVqfv5UJK7vpYca2X7XFXEq
9P6YolLC/Cjoe6797MKTYlJK9ZHbvcd2970f1kRYWrMR1wu07m2qmN/x4ZJaGzAkonBtZU3HBaNI
EecuB7xNlgNFa2aPHA5YG1OfLLUykarkEvZEkAjXi8yhOoSxTHXtiAcd/ufy8/+NbjZkp3uP5BU3
x2KpqlmY5yyZXlaguCPVwcFAzW61NDa+/pVFEFIRk0yHXXXEZESAcvb8BS5iHmD5x8tar0J0bLDM
EdA/A1r/sHuMtct1I9AyWr9wUL8gRAhnXZVmawCKEx6HXSWu718u0rMNERv+/cB5Vf11Y+ioxUSS
5nUaqY5H/74SA09mgvCgFg4IX5XVOTKqi14DyoClwJcTwAU52AwrcuZjMgk2dGby3rjzeDbCvJ5M
dNMq4gUnL9DXnrJPfzlouTRI7U1qdewK77yAW4z2DMDkby2pWlgW9AyF1b1x5hkxcBb8yf/NhZsY
VNlLEDANMevGLXt64wabq2dYnLsS/QPLwz3EgkavQcgVoXFXEPxPVuE4TJ2vn/qasy9XHrxDAXOh
nCgYdlQcM8T5UQ/9cZTr70Qnx+z2cVEUCnsxug8CjgnbsT3OifsrWbXu+QheZuHsXKwH+UbYr5AQ
KsVQwtF+tUxNQ5iq+uqo+vWkm7xci+/swnMwh94Vln7VPboWEwqIlQr5oz7VOjMdHGrKw5KjmNDg
gs9kDdZy/LuGRhE1mneWrF8jDt9xchHS8isM6UyUlvCfb9u93CWArBJ5GYzi2Mmmg4scY+3OPTMs
hA7LHxquvXXjjRnFmeZmIp4Hq1CDnCRY5Zuq0jlc3GYHa3tIjpQP5JemF8MfiNJm/LUG7gC5Exp5
U8dk3rZXRz26B2VxJBQ7uAx90uQci0bqZ+G5xmG3e560t3nKHlUYQnxyvoN+5JV5/ydLXNngraYp
+CDCvkslPuBnzx7q4U7yBniiJ1FNmCYARrVrBeMTQ7qRJs8wiKLKjZfIYBe5wrPdOaG/Xeo+Ttak
NuH0r+agE6pAVwnlvvmZJsP7Q02MasAnn80yw2b3SliCXdSt+K2cQJdKUJpSWOrWXO238VKFfDvV
pgNUdUZIR3um6f4iMacS1sncVjjRy4SSJmPw2CIbHTgKKLxSCFBSGgM41oFb7Iu+PTbtXU2fm85q
rbjT7LdaC2IuiteKI5TsNwVuR7cl/5NMZYs+2r1ztJRrcVf7Gk6PE1tjBbGwDVy1za17d8y8W08S
TFPWj9qMY5pLtYi+6PrItjcUbPLlUBgGIY5Iv9UwUsrditJVIeb7JfXGDEjHuSlYN7TYFfByCSMz
9ymoO2IIHBrgE5QzYd5wzvl10k8fF4ipq+Bkpg08+ZmYHlAwyrIBy8ucxj23IxB2Elia49kx5ErZ
NVX7TEuKzoefNT0iqKgfOsmve3MUfJu/sgNIriKYBQ0ZWeyO9igS9vXPBxrAyZAcYqTIg/cHzbby
WE5e+x+YZ181s/KpPrnXP2gzVWH/sSpoKXfpLaNg1Ms9LUtxos1Z8O8x8J8S/ZwJzWnDnVAqk2s7
Y6VRCYQOhSORj+SpGeQCf+q32sM0nMrtY89MNcQ8gdAcicOmYgm3y6f8CEvZG9uVuZZplyuIjp50
F4OkZ+VwOzsp5NlU4X7ud1OygP3qhEBQjaX/Qm0wdRk5KcKrHL4RMXO2FCuhdbjGt0zhr5lNeSyo
iqwMN0XFXDNDopeEQtXQc2W+MvpfEkSgtrtJ4ih2N9BX1vdaN3G3fzHcGjKcazGBL3P3mHEYd/n8
ZytJN1PrOc6EXnfqII7JqUe8nfyxuRSGf1CKNhixrmlgiDWz6WnGKTmgNFFQEr8q3/mkPEk12dtv
dyBMMIXm5fgdScpSvk4N+ep25IkjZbOm2hH8WuMtEKAMVmUFWH9RtKmInGMKKCwdjNmw2su5qAv+
UlSYmXZbiGbS4mYiYKMBo5/x6Bdmu4d2dxFQaUvtQ+H0vejWpV8D6UabyYvHY20bVnm1KKKIMwpz
C75/DiC7kRilQKoiDxjzX62TfASIMk12mHELUTc33DtFkwQH8mZ/H8RpQGQjXOzR6Dmo4pZpQSfP
Nb2H6LiPckmMw2yQCUmwtNYZIt++mfyUItzWG+yGqxegaftX406GEOBPD1nWW1ugZnNjk7kxqMb3
vQ7dlmq5tlu6x+cnMBzm90b/9LfOZB3QjOBrygSJPi+eb8XMqHcBj3SqC+lIVc++FrHsnLZUxNKO
4ouVcGzbfM8O2T1YEtdA8feBWmaDzx8IpYMB1EclcVnaVUVl3WY2EjvPuz0RdIzSP5VvHPsSzdxp
V/4pM2Cp5Txopdd15K4ebK1jVK5bbCp121i6JtvmmDlNYRMzfxgkTuSjXFwrtHQHbwlBMc/+MdGC
pu2+mmHlhPfPHo+H7sT3hLhE7wSWNGvS2B62EDpV7oBk4tyKG1gAZJ/REb7Qa+RItswuyaR1OMC3
o4Bx2XrdcoQhfdGUPnWc8GFBbdqWZHtn4uRjO8pl5pb/+2XURmVY7kSbhKXU2NOlxOI+6zNBVUPa
YuOmVpPSgvkG/7LlUxnx4N3ajGMs4V3Zbx8nlXHTnFpC7wlAJO6j+sDP4fphdGfe8F9b3dmB5ld5
3EbPUTpOP6LmN4dPBy/ODbI6C6mQCOa5OI3pfme4HF+LaikdSnI6ZLe7qNfgw55C6TtWpxCJNMmX
poC7nD+ZynPO+UoGNxgOW1BxbSpSafqOZOYHh81/7OCnImoNQIrZy78wp5ywmAtyijWtajoZvn6K
hyrYcoimS8z7ySsGPKI42ybXvqlfVoZKOmZYDCYPFsYzCJp0lvqMURyK088M9kUrukiVFCaP6FFu
5vmYNW8WlYqxkiBXiA8WPiRc73ZHKzlt4+yDrkN9amK6cLLegqTmgmD+BLW922JFiNJ24HMWkzxg
eNUe9ub+i+wRr9AqxwnI5pYw8EFjFFk6jDwm8W5mbWC96R3r12MiS6QnXBs8UkBQQltJrMlNtZrS
GZalJJ/4WtgnHOKtSSVyhofO/umtdhQKI4IoeF8CMD2Q2kssku4y3egsxDfw7gTw7/eJ6QE4VJ2o
Yx05E48xzNHgnxzx+TXe4/0qM+ZCcJMee4n+3xrvXwra3D9NXfLjMLEo/7LVbD2g5jHfbirA55N2
32YzYGZoKiwxs0hDZg1AIz+S1W0X8T/M78GT87q+Nn0za2uUGzYR23e5Icf/ORBxCrd3yvFdN+F8
dP61RAjuRh0jLt4ylCWPDlaTQWZed98+nATu+V1mNQYpDeDWjBuiot/M2j8EcS5SsBSPauQcUqCS
vsIotBSoeTqbDdgxmmp85hxaBThk1fH+hYGL2mgGmntXLCQoNX1fbB6dQpd/gWBrW/uDJEkr827v
nH4rdyZbX1YppDCemnbP96L7GdHnszAl50rlmmWwIFvuI4weLCDgWgJyp1dFu2i2wvBUkjb94l0U
uE8Lldb6ZxzkJlfLZhKE9U0lzD8HlsfP7yVXwyQOnTbRhKWBIgF54k4S0N5y+FAVLEJO8aIF2zUZ
bv0Q3a+skywk+kRVv9voRMPyMMC2pn8MQlK3Nn7PlfW4B4ujH9A3Sno7+D/ewlxfEVtDA2hFV6V/
PJsaP0MltpXaC7RHaedg82jB3IDCHEGb3IGWc6WswCdi4/l2+NJzNwJT4a02y8hgdxCke1aGaTOw
UWaxa56buN7k9mX7np9UEuq9RywgOgYE9jxHo57ZV/vsTTpo3Lee5Dr9Qbb8GhzGUtof/w2bvni2
lbsKZ/EGAHDyqGYQjq0hQjT7b2xtmMfaH0VToKfTIh+BNjsoefRot2EgtEcG5EVPmoF4QQwfovpi
OgjtH9vg2LNpp6cIej8W5S+rgqm7/w08S1cNGl+S1PUuWrFV0BJlmNlOpuvMvvxbVTHD60fC2BuW
7dWdcDolWZTjghSSCly9Rxyr/QqCba53sr78EiAJW6LijsslEtsWEoWnHxnxbzVSikRJLRrtk8uz
30igyHCtVP6+k9hGeFCpqUTcO6Ty3j6qfvq+c2LyipAIVg7PGL6MnxBYo/svFGQb6qH9sRPh93lL
Vuh+LZUkuIiHUBgIi2ZY93nTxndHFqE4aQxGVqyPkI8JkbjLz9JM/KOu3DftYiZRxrFDdl+on+Km
2wHDGJMHegDQPzr4DZiQjIGtSuOLxh/erKF41IVolftvlfNcpjH7knA10z2v7w2WqhbNikGlUeiI
I981hXRllucmzZj1PzAJRJDAnUx7xds6xgFlFdq25IPT1eygcLhOiN3BrNwBNedgvUarLnT73p1E
l61W1MnY0OrZy1MOLu6/q67JrPNtNmN6Mw5yn1Emf5ypt1oPhzYJZkZzQ+45yEag9opgJ9AsFt3H
8Zw+cxx6GI7h8+oHnKDW3KlRtnOjEwOi2TD+HfugoHqhcFXu+eWb3OJCPBDGrFoVLIvqWbU7o9w+
1wGtEJ9kUMTetJDbIQJPKern5GIejbti8m/bVYhC+L03HjqjRb1XbTwqEPR030G+tskG890ICBSr
PtWk2GA0buXE/52iYYl6XT3pQk30eRM9CREYlloEnOWkeZ78OW+zrwna9QyLbh+2CSy8yemLJENA
bPPBMWoyRhdY1QIqpYm/bXhH8NWnDfdR7zA/9JdQA1dqnu7/X2w/4jOYRWMqfyQ3zNdK5ZOa8V1E
xJAlP5Ri1icQOFzlquEY44BqR9Ma8iUzAhZZbAXHMcjdoBGGQ3aKi4PBeK5Xh6B8h7ecs9pbxOBN
WGMp42aIFN+h+kCYvkPLC1S7LQVzO2Vzs536SN9dnZGLMx1QWwFa4KxtW03abfKWMvLW6s+xmowC
wBuontAtmRrCdoLSrw8Fji6o73nWUSc5XZGpYhUy3KQQQ17ELGFuF+g/8MwZAoMX76fggJ90defG
QGQFYxvcfeM/bqauUF+yiN7gq2VcqxF5jQiPhGk+LEs1T/GG4Q3DoAoPMNyWRiFmP2iUql9UAKgM
q8rTSgm6uAc7OcNVcUQr8KGOVhqGtUoE/IzBPCR4wF+gzrZSVk4wbOMdBk7Hoy4QtrP0Kb2jjveg
Ra4JZALHQtJEQgdSVe9Q0WaB0arZiHLPEx+koW7lYtsqdZFOO1UpXIY7qdVQOfJ/N73eSz63sp9x
IXiHSE9F7GqXgheoPTUWGqwWwH0f+iBrt01Ai55k6tIM9Wy2yOij5/f4zwAqbpjGp6d3ilYXnoT9
sd6hmdhP9TJQojJl5QG4RMF86lRY3g1ohbtUWkY0Uc5qkonJLTRr228gPjhRsh3sumvnPoITbbUU
eHzjX4rFAOoWg101kmxrtIQeMp5wtNszccVuqBcp9y3TZlL+jiTEaM+p0iYzsBKo92vvsfeivBTr
VK69p/GOMUvTsDx//0Yyi/1wLBARR9IUKMyqr0c2iCrEkoqoY94dkFXMNC9eJ8ENG9rw7T2hFIql
/GFX7YYXgaFd5QiprGSci7vZLZP081U9SXjsBtUj4awKGeLK3D1k0+XBV82xuG6xxlK+jF4dfpDJ
BQCMbeJgia3zX9+L03JyzN1JgTkjIzvtrC9+P1xfV2n19v2sxDE4vLWGS8Iqak3L/lhEA0P1GI/E
RqUHOYZQo1RLLyPa9kpR2WBXGo2A6+osOicYgGmF64Cq/T7B8VlvZUh/tBhvd5khjvjqCmhZK1tP
UuV9yc9Yl7DZC8Ev3Wbu3N/MfTO+/KARX/Eff7LB8kZcptZdLed6rZpt+mszb6wadQBIZGIz2LqT
csAD8+k80SrDS9Rtc7CJUmOcsEo6Urtl5tU4tLgzSxVWzhAUOMoJKY2XMFgpWBPHnO12/aNaG9aJ
x3PhsYbhBHwIiF4xWfQu1CrsimT75Gb5e+whp9Sz/7Chg3ueIjTYI9DQ+YSz2681sTDBII8RNLcr
IrbqwrWX/eEOpO7UUHGXj069Fvmp90FDYkHX7+Ao8Xo/bRq1Yrjqmk5+Hu/DgHuwwwzCjVUS8bOf
I3mgMIoYDXL/yVLb/6sxVirmYvPUe/Lp5P0JYHb3BiJ73Z5uXIziQZ9/fb3z2xepAuebFNjiXMFN
/ksbWju3ZSF2IG67QIwmtFDnPnznqN/JgjmUw22gXjdAaREXsZNsGKrf2KprHO4r8qtT/WXJq1rZ
My5CT+vTe+sn/Q4AwyHeZHQ/l1CMnMHD2Q0xZdnYcUVFsbXd9AovQKZ3AqMXYfe3YaHY+j6KjE3Z
hz8fWnDY8lZPeKzeJAdj9FaRLWuaclU3/Om9EjewiuBuPkTfC5z1WPu3ivcD+1HuVYUj1iTK4oyi
TtkZ3UYXGV7XZvjaeOm/SB6RtVZwcLQ+i/eASHdHNuUpC0j1TnpEFAbnf0lKv22w/HzRkB3v2ZEw
qdzzeKvTUF63N5W6RXWh4mOJyti7cNbN6wZXHNuPkNKnRu85iHpZ7yRtwQJgH/izZ/WIBrX/F5zc
acSfYJUSU0Wd0M669C7Ks9ew6PesshNSf0gQ00Xc2kcFuER4PVIliAJVQi9WA3mj/NviSDm9ZzrN
p3HmqF4MICYqNfa3/sRXFSiC/AnOgUZ4DyAl93FZT3ZqzmPQljTd2xTe5qPloGXynLMETxlcR8RD
+OCdaEJ3rC7qWvEAr/aWcoz8eWrOEidvrgXuNa1otbxJ7UecBb9hheOLxqS/MnSpD4C17hLr/WdN
cjA4x6ivPRtS2pkXX5T9R7glIEgyXM6TbjopwZzLYJ/+xDmeomsIWDgM10VO2RsuNJEQf83mzo7J
6IqI8sUfDwrsp+1Q6jCc2IXQVNDs5bo+NYvp1ujoX0Jg2vNFdy1CpX34qJBS00PW4x6r32IOTlc7
ln9MQyVMOdg7c0vonQxHpRuVn35+X0fkSVaOmVtm0M4Y587YUXNUK0mlvwwBq/hnch3xKRkIjgbn
fH0/Ckguxonjd+t5iXkV2DyH2KlgC9ubeAk1Q0l0QMb8CG6GvGRify/wyOxc9bM5WO/iPPuVFtEK
MxKMiO7k/T7aKcQ/eO11q5WXJeaQ6CCSG3W5e4v2iWOUuQD3yiDfzYHzBJ1hpgdIkjvxdUCIdnM4
Jk3+t0oiGWGnJ23QdNTY0hrc3ivfEZRe5zjtlnQXL50rSEeF+DAXDpx61K96U0TdqSi82RpPlbF5
hCZtlna9BmBawJGPZtfP1Du6TLRq4T95PmK/KpMQP0Jv0nAPwdnghIJ6PIYdoTSRO0qDU/+kzW6h
N3B7af45O4H5/Z57eZz2qEvLTKMwMRBvhfdWO1igXPlSCfDgUqHdbtdC9e0T7WvE3OM/nBkSNRfc
SFGxTgj14xe6QhGEULgSOHKidjEjeVCU0ymMJ2LrIqTrzCAtsKqiQGyELzphZdrXHNqTZEjpd47x
s9BnImBRl31tBub96DYtSsNFg4ibj21lrdZzekoWCLNk6mwPD4cz7KIFjsqyOSUobyiNUc1xBK90
T0eXRFneeas36ODOGhHVBdgvq2/yLc1djRK7s0ZTgkx6+paoHbjkvnpOYbRhwF1zBqrW7Xxi2XMs
rGWhghNwuhxuDgD1frqXo+yBvoTacE/BCb2Hz+biHVhsfeSbSXgSH6CCN/1bSSpfqvF7OLiwr3/m
w5cc28dvingByt2uP8Vj8OgyvoFw0e0IcTdsBU9bDkX5EneUtu1WKRRz8YHDaIoPULyQhPTQbaqv
W5d6Artl8sz2NYsD2xAyC2nfvJSTZxGs9p0WESMQsgg6imB8LxaAFEzGWaBrwfofnGL6mX55B1vy
tK0EkoAuekynkCw0N4ch6xgO5nUMhsfSLxv7kvPRZuV6Wx9CHL5kgd+PlRg1NxOxPFJfh+joHDwQ
hs9xxfpVEgX465DPzLp5yroc5XntVahGowfo/pm++5FIpiYvt6CnqPLLvrok9E0EomaFi87Wbds2
Yc+PKIHB3haAZF62IlTFPylIYUDpowyE4MptXZaLZ7A5KMDixIztxnfG4r0ICNzRcF6qo3CFXk4H
KXyIlqB4enSfbGiO+/Fivd7PNJZu9gIoE6EDTe/L73dWpi5ou0uZ+MEhXeqr0ASN014EoXz/urtm
400cIYC0nB8IWEjqn/9Z70bCA/qT4QM0OeDWoD6HV3gx/7v1oN9E7cZtWbJcLsqPCI5+hagwzH1d
IRB2Wkly+gXi1Z2ajS1zeFldEOHwitjexo/ZRvbAEPIu0MIJdIrDMJIbqcaJMj74KK/CltY446M6
zUl07qHXiaVhdjOAwg4NHvNE2DMVGVr/7/YPYePVoHALoaZBcVwlWibILVd7EBXQMbunJaZBI1xD
cwKKoS1dnN69X4ayRaPgdCe9xX3rtSPrfvrCb5IsiZIU/pIB97ABxN/QWaurp3howS7zBVFdvYw7
FXZpJS8+xu+Pdbb+lnREDUuJqnCZh1vG5ItocCgnuXKNkPIa4S5gGGO4YM9U/FupNxHXptXSmGng
Ta16OP0Dgfk2PCLPPdp7xTvcswqGeRKFqNtVQFPz7FYsD/IYay01kpkvHUP4eI+/qUn6UnyivWD1
VZYSp3ReaW0zQLG2qmrftYwfWM7xd+X7J5dyY6otpBws9Au7sW/TxM1A9jUwL0aWJDFGKg40Uhm0
y3ZGqZAAXMVXJZ32KMehoAY6BXY5Hpr4BfkdpOGMD/pTQLh8Wv9RDnIuriX4eYHbBJs8DHqkVGtg
Y6KoIs8Y/0vQyqz+vAUr8XUy3WlHZ069pxAf6dZZJPgjgn71nSHbUNO8XuHxPTqwxpXuulHBAvJ6
SkhLWVO93777P61rnIXDLRIPtPtI+b+iatYjEsaI7qVmbycWb3suj7KEYKRZgmWvzDqgmBqBrhmV
AsR82G9EDdU5yMQlcFTC/LFNqg/f+tr4Jv6tfCxQ8hgudixgk/8cd+JLKmAeWE4NGz0QTZ2cv7SV
/OmNNDP3tMlKH49WPwWxmYS4M0D087xXKjlfTT6TqHpVMi3nYo84Tdc9vz7ehs2KMXxLwXTxpf0Z
R6IsH/LbXwSxvO2EqxcPM/VizI/jfibqgRYTUo/48/E0K0IF/RaEhO8G/1Y5SdEg6+3I7ZjchXCR
tyBqKQeZYtMbbHAGNQODcQGm9PMeL+2iGU4yxEoNqCNZ5osrv/p6BmzughQ2i5yZlgCQiVCbA8wX
kK7oB7L2OMg9I9yB8mdoBnmnm3AwGUNlsg6Tiudf7IePfj8K5cFMM0ssrLzbfI75NeUCPXRV87HJ
peB6DsbvkGRURPF3ZwkehqDjv+ENMApyNJ31FUym3/glLM/z4vEr02KTckAka1g+RY6GY2h1ztre
0I1BSSdKvZkSvYFf6JfOxTYNaFIpABThh8MhxFWRUcxUq+/8VbDuLcuzA2D1ysZtvT0FexBxOBd7
fHFmOR5WViUWXcx4e3YTOa3gcJpGyXylwsDhy57DH2jj1sATwVI+IDPEZf4xTO0DxCuf5JYcEb1b
JRww/tam/f9SA8dPWITleewUFWsSt0SGxcIF5keobJpLvMFJqbpnqDnKV7m2kSlXTX6PVyeRSBMY
rsqjvwWuKmohCkVVxBn2FA+W3vDbeRf+EmLFvnpVY7h9c1cbQ2UUERKjMobFsXKuE04nE24+Wx+E
XLBxdaqowvS3PMInqyBIygYZFeB7QVuWumNTI1gRFOf7UY7DcyKK9Su9DrZwh18vDzvRPkrrCRLw
HdGIOKUp0GkxkTaspX+Hqx70703BV1C4W/nbRFGFk9JDHDT0LC3kFVfe2g5C5sSO5btdx/jxGgQQ
7CgYeSDA6YQaPYECMDuJI61yqXrjHWBaBZbPJsGdi/GY7odtojOlxZAiww603PmkqtuGTOR8/zG4
ieeoAClWjCoc7YAx5jkBd56WzA/Or6la0BK9wNruBu2toorOJ/wA2pVZ3ri9UCbHt5mfd/Kc2/6b
z/SIVRQT0EdSVcwgpMa8638gajpgd57GOEDuqEIsZ0bQH5sXXsN3aE3VuynS42FgizmnZO6LJ6h8
X+QmzEPyqBj4RfXfrzNMq39+iSaHDytbUcG4QFYw2nimTKNVU+P46HyG+8tgWdfTcrLT6HmJ6V4P
kGIItbfEuaC1drX2jF/DFum7PsL33NKBkqtEo99p9mKBwpevGhWEI44iH1lV/kz/uZDtFAl5ziYn
72JnTSyH8EzKMH7O3OBdEMWXxXr26xisfFUPfJi9ztLsH11kTmuNIdZMFRKY/8j6T3Sh4r64VUFh
hxBLZkG0Wzlcr7+sC1MEAFCASf74W7/TpgRgyO2NnYWhVpfAqxfL8fHOztUB14gDfNuk/FVRe9ao
BwJpbKXoxft7ULokqnm3r4GelDUeiL0/O7JonyUoEOyQAglUeCcKu50Ej/u0YIBELbwof5tiaDA3
kzqwjCxYhIuGA3z7yRRX1QUP3P8V7jGd7/VmSdaQq0+wst3uH2hoF+wBEyzAYSde7URjmZwGFB8Q
w+ni0jbYd3BuLQyUnWLKR+H1JF6rRvzJCVtLba3evJ0wamkxe2x2muNNklORva+cQs0vHjoJMh0v
1YliRrk1ncT6M+ARBEF3FQBKuB26Pbqo8Ag7BNTzar29A6dwNbMeWnpNT29xJ5+v9cNwckbIIMVN
MP4pfLf+q1SNvkhIE/zH+oB4yZgzkmCRYpaVLoVJrYKJgFhsecA6fVeq+dwiSjSJuCIlFP97SuWS
7SOPWPQ5wV4/tOjzuVyy2l9BfT58E4RdD6J4W6CTyjVamJJuHzMJOU18gTSVunh91FI15vEuUSwf
YYPPI3FRlvufNnwiPoHZNepHavlNIQJqrMtn0c8fK7F35DrysX9cPaeEpjQNg7y+2h2CeVOXxIvp
/eh7WtgczHws8FbJTOJhRn1+uH7nqTLPHtKczdiNHAx4d59JxINitVMcZhuRxi1RZLXDQm/Dr/uy
FCGog/toHFidqF+DWp9TIUGmwW4CcF7ausYyiN5c90ejbCcZQdTy9v4JE2js1aS4Io6dqLYggflA
oev3TSuESyqdjcaHJCmeUevhgcyknRPNu3ehcLOpFefpwbmw+W3doRHMPP65JyODQkuNaYRN+5d0
baugP/a/zikkuY7rpeYKmLcaID8/935OiGrCTVcSSbiO6B9PRySGUS7UmjpPEOIu7J01oROL8edu
JCJpfsvCtJzpnBf2tyMrZk3iJd3C3Y7MPrBLRiai3MdDfrMfhEVQKON0l34TK0QHWr3pdTYXKu0N
1XmI5HFwKgoVOhX26/kxb1qPk6JDYe/BXMQnVkvbrtZ/PWquJw9fACnBZuReAF9SYf2M3/3yofcO
q9AK9sHmj7o5YYR7+Rr87HaWNCA7CD3VrWYINmX1myQIEGCFAJEyf5znC+K4ZFWKqHlgZ3MVVzmf
9GnNaY1YnbQVmDDbrU+ARZEStMfr0qSqfd73GzXRdrX72LOHJIYMDIjPFTzjFlXcFNsgpqEUUxgf
ocCQJ/bJDTWbe+xah85LQEI2OXnShOuT2CULE0RxbkS8lMyg0uppN3r92u3j/57zoMb8p0LyNpDZ
ojqMS5nn8GXIGjLTSZgwp1qF1yM8c1M8vDmrYB7vs1P305aJsFYimjF9gVDlK3DMA8IIyHzvuVia
KKoqk3OjL1oGYGepEH1o5KiVDgnRGDfmnNfHkcoWnNH5WKykUmIVL4YY+RDumyOIEsDx27vjN/zK
X7FSTpw3oj95NtvvUHzgGUftzgy9VPB7Stm5YKq8mFx3RQC2QTGZlfYpfHMacAnUmKg77+V2NcMv
WjUuUaxBumlOVelsuyxC8v73gkGY1pk2xm/VLPsERXhsHlleZIOAt2FTnJujKHQ0YlB3+8rheuIQ
aTfQsW43cGqH2JWZ9SUcWTl39nV0WfTfJ2BVUYKBM6WMhNIgWeURTNLkQKeytxNSWTBJRCtZd1sa
8cKN5AfjzC9VpYhUQxkecSRg/wybEmw3Nz7mcT7XhnIDnBoHVSWNu3c9Q9o132hRa5NFoCFlXnyi
taojvfrsaANejJIWGxdTCznAwllfOOPS6oCi9iyb4IkCaHfBhUo9srJIzLmL93YbSTFqadInIOcA
cJ0N5q7Gj8RQa1pfC+xw0P5xVqdiwt6aDkP4tzkNyWI6ZQay1E71dgF4fgeQ6FDi1eLVHau4q3qK
uSwwmQ3FAojsKy8nOmJzOi4KGOTNWkCSu/CO5mfQ0MRYv0sXso3gRsbSnGYF4PKp6ydBfy/J7+4O
qqsTpfkKfQxaUZ0m6D3poG8cW5KRTjF4TSPAvKrH1dRCxKGdVo8U8fTZTHQ15uf3F38t7TfJGIdV
hmvaQhbvAuQ0ZRx9i+zRAZaSvojop9YZ8G30JxcHEe43qRGzqXtg1Kjj7gn5Dn0X+ddo+/xeUMFg
KJ1ex4d/mN4jN8maHrTW0wKr06MF+gdKMRjnIxR1XtxDUoV9tc6Z0UKx6mmV2G7tH8ahpkI8GHnM
C2okdK1GhdUE7RD5uhxON4q122XoZrwT22siJa+BbEdyxSqa4ZNPNbgQecFj7C9ESG+7DZPdC7Wm
lngmXNekGjgg5l5pexiCpnv7goelSPX3HTDQL+9KWSFSYBCuks1h1Bph8Cmpi0rGUJNB5adHG19E
U0UKb09c17JeHzLuk5rD+1AwE4XC1uHuNgj1IPA0JWdpkGHgX7NfcFIgd6zzuU/q2d1VOoZel/jE
rh3SDlsxMmkdOPUFG9HIaq2w1Tn5F6zyGUis21Du0wWC8/ckuttWR3Q4aZKIsS0BxCWF0s4aci9i
agpZzxqZcltHxp2+4OkmGXbZhHuXF9OWsN1CrhWfi/hmLi+rn9Js0sPRvvQaUkoDlWIL7f7gSIL0
Iem1kpEAqWMjaG12j/MzdW5zt2RAe0Fzfv6OfgoukEqHzvnT4+knC1qrhllNOksYQIU3Tu3RYpvT
ycJ1h7HXAcu7PVp8ZHjJluUSDxW4wXfQbRp/F51U/djOGdilYxC1pZRJHIrjKz1MVUl0XYQXFpAX
9E+cXbFCzxtF9+Fz4HCv2X+ddmU2688bySEJpPf35LHTnsZUkUp1JniQyO+VDpGrnDajiEcOmuGC
8o+R1KAGaTJxdMRoLQmhF/vIExk/FWrtj7aRfDGDL1lFojcQzHKDiKMSDNQAsiysAo45zl6y7IqJ
S9sow7Z2hnVSem/cJZoLJIvABH+cYWCgthJmOI3kTx3NoaFgQZQLaaREy6YXve9+7qHj9D2pGVX7
aiT1I1S3dIMdfsVymgQlioFF7jV5GNvBzVq0T5cYClac/Hc2et2xq7dDUk311piSG7CHRUW+L8qa
0UgjujK/OTEChuwHJW5nTJ34udqzWl99+z+6QKnPQn76noEyE0aO2oj1Si0rE69tBqf1T1z5+Q78
/bqmjLlnKxf+XXnSdHUR5ckHDA7586HbxKseOLfK34xvtATmsxq+2Vi043dZsJwjOdoYrGF5qpVD
Sw1KyTK+wDG0pcC5GCV6GMj1+z9JKDW0d6NjCrdarke8MbOfITlo5j/pO6xxIhowcl5geBjjM8JX
wSalHwtKoBRdB74lMT3UGKsPsag9ruyeKo7GJNWgAgEaZstNOlfMA06W8kNXLOmtS7HO1/4RTTsq
SJYJA+y4rgJVlJ4UiIorcOCc5X+va72aiv+40aDy17OUV5dpGFaybS/OJuEVigHWyL6NSuGQX/Gq
PlT9u53RzgnPfaCXAw5wQZ3ttwMQN/d3VzjbcKeXXvMdaWHMIgb8UUiLwOfA7TCY/h7AtzWiag3z
m3rPMdFFcygqFHF7QXIgi7DNpgQwOn8zLC1i9C06iCjX+lseUEoMpIRli3jwyqVxGqVF1E19vbe1
vYSQZyjenn18pA8Nd3OFyG7uPTqDqU2eC+eQAUa+g+6OHIGAKYxvTHsgzf9m3N5sXfPqJAMQrMAq
OZ8p4aRn6KnfPtahB1w00yLcpkWh2VjikuKzMcjZK2VkjUQbP84YBasexBgDEo9xth4OPIWH+P1b
XkIFt50+DHuFvNcrnyJSmHXZYUPqlOjkQt4ejp3PXGVBBXfwzvTkbV3DymqO3Xr5X66XJ1hyw2Eb
7bPGndaF6iP2yFGwg6cPkTId0QbKnB15/bvhcF6FauvboiRD/GnHYxWQCWI/Tf41nU+TTSGIE8c1
yrCn6QZll7i94ShJv/7RpYJmuDId0B/EjWjAkZc8rKm+EZbebqBAkglbDUSy+u3CrsPNs0cndL96
wdgzMZaEityxRnE7jNpbnI42nW6SHCBETSTcz5D3OtM3vYyOID5ACyLiSpaPsk8mnBZ2jzkWAnaI
2tR0kIMWeGDyvQG2UGwNExcJ4HxrxmUEnj8cMV48uw9NG/QGp/bJMaSalmj6+40aBrDvwN7/x4kX
18nqbedk2lztuRJEjS5TT/566Y89D4DIjX1wU1GA/4iylmFKu77TIZs1yltMTC4JYG/sBJ/MilMq
61bQ1SAoU0DQLlXzmPVti13+ImYzdbR4WYpYKgU1XtnNvycUbQVyCr/+10Wnam+P4MsAkWfi3GIz
ZKZ2W5jeo3G4Hz+R7d2yqY6CwhxdEuNzIOn7O7uWFHwleWsy6hQnoF+UVhBY0otFWcAkXWPiD+kz
49puGHEYIl/OAmprFK4nyUZV/ZpRn8QOmzlrj/+cs4PDf8BKhGb44+xU0XmMPHO8n5AJjBzWYo5M
ACN2CsYyggt37dAX3YpdUMfOKtplNTAyjXuRixLpT+DbrBmWhbiABnLQ6bR19UKQKHl8oKNmicr5
uefkyGQ/+a4DByKt5HTrySeKuLUaGyDupXOf8Lafn0dg4PIV69Ke8hpBiiyu22ZHzyjZB/aIlJtH
6GLtZwNrx8urKOPqmWklxSaqlOT+1Q8fvpbfjmbyUb8Cpdk95yHQcDhSXkh9QVUMOuFOUdE74XG2
2RWH3RGmyJc1d+xah07HXI1Xunjgs5+IpQ98bhZw4d8415Wm5+11SNgQbsjAFZggWO5B9ZQEm/la
2y3fTWoWpDSy6MLKgogTqFID4tgD3LmSuGx8kp+7eJfEX12ND8RYZ1fvjCV2j07KM8z+dJHb26zS
FSMy/nTO6JRZSeHxgQB78ytK/9kPKRTVGsZBkR28K6AUzlNPkljWMMMDl5GUHrYFGBjlnBY5tO9j
nkglhaNDzZeAfrWh+LWQxaIznlDqkAwkHv3hivBpYmdqH+GYZ/nmFAny1NqvpgX2FgFdSmHtbSf7
069dBj/8wyHw9rIG/4NBJNuB7qWaAy7NQjmdXp965bH3kf824TQttg91vZ/EFzThpTvgH3x3U+NQ
uzUjqcmivveBbSdEnNJ5GAVsXjsuERhOWzykTHrm/6+mDAEBrUsY/QEeMknHSgqTHbHKMkuf9xly
TUJwsXGSwkYIq6OPgL035OjR3VRyFCeSPnV1it2erOCJHy4WLYxpWVgKu2PLm9GS0ceMp0hBv1i7
pJAnVSl/Nfv9X62vg4bPUF/rDzsssBXeVkpTNDu5qmXJR41UhMCYK7O8OhK3ZVwS8mn9isVhMLVM
FvombkDRjhVBzf76TaXGt7u8jPg/AO5CWbvtwUYypEJRGDI7zZwiLzSlA1ZGHTblaGL1fqEJpPy1
RuKKHUbdPOxualxwfQ0eLxAk87cn2JLgbCe91Y/Mcl22pxlDbZkwXmaWBsM0nhYxgeoOTQ74fBHa
11b7BZGC+U4bcda1saODXo7Sj1Nrfm7s5ja/UZDccsF8g5DFRRwc+SNAGPFNocvYmDWto8toBZYB
l9xo7PLepI4MOuupAanBmd9erLQ95uKzF8h9MFd6EyqJUMf/uiDk2goieoL58lqtSRib8RUoVX3L
BnYI1rx9D7kLEtNF4uON2gp8XqX7lTpdJU1kxsOSUQLA3nBB1EKwu1YGv1jPoXi05NJ2/Q4XGyiN
0Yb7fDH1xTfwOgN+eaIEVEhjdnOdFASe4BbFkqLx6xMScpnNMYhIh05oDEZY7yfwPqmvgYMg1ymk
DB/lZYvh/9c2H5q7Lrx8mODPx4JQB+sww22VTRRQISqZYysnVy0LuO24SXNBsDBKJqXX6WYPXjgO
xHagp6eIoqDwrKSRZcXKd75TJs4OrqcGSzgcaBwWpQApzYosGnLYr0VvbcDwm6jUtTlOTuJHrI3d
4ypI4FyIN1iXgvCetSaF9yMRXfV3iEmNISa3MphT8PFxLitftWbwbvU2o9+I1KDxlES8/gppOSfZ
vxa8w0T2uHU3d2eNzkI6KFAUY4rb/yuon9Qesdkenq7NlCP8ak9bdISsPJV8ZrFO6MD3le207+px
LrZR5RcFZjz1oIfI26EDW2G37KWK6bletnj58TYxPh/kp7TWyNwVKtTaua/CfG9nigA3zWhJHDLf
+LtO0GVLQ2djIzexY9VEbUiJN9kK+6rU8MMuP2e1xbUe0L0gg06wIUWdG2oU06ZTOlILp8T+iD4T
WQWJanVyvy8yM1bKAVM5klBDt7xto6dD2mGfXCJkm0ObxktZmmei6uJNZXrAGHDlv29hjE1R6Mnf
BUYBU1ybH5pRKiK3FHNNQ/r5veV8m3dKovP9h1SlP9OlM5xrmmfnLMke67jggI76GwhIReOM7B0c
jl+oBASjGYctoN7YXaaeWylFFVSIiZ/Ynoi695I1RAEG/PX6RYTmjF1jnDaacfgEcrm144zX21Ed
3en0QRjrStYAfcL/lUOB8gxIlrZpGMUDwCQZ9wcgmbc2e10VMkcj7KT9+cw22hCZjn2v/Y4OpYN6
PaNtj+Ce8K2pB3Oq6E4XKnS4AAftlsILm3umrT3xptXVOvyAyfqsJRntPucp1e5zWtCOp1IOuUyT
7niwCyZ4LszOvZmEOkm5zMtsoY9TpxrdQuJBv7ik31oWEX/GAf6zrnoNdE0IFKnRNrn8msy4C6xC
EG47fTw1uAl2wxMjqD2ZFtVn5B325nd8boajJR21RNYsRIcr/2uDu0uUNxwnlCeY1c7FUIeAW+7P
uZejn50GJ33sKGzeofBzTLQPcsjf0/6xlOTKPsZfqXk6NjMa+J+E0OTRmYmA6AI3siDEiRcMHSCv
cndtxmAcxLoCMdiinoUD2wUePDf0jaB0dbp5PpGDiDPm38N5DjHeffW6yOuHPxrZIdVBBd6XUl2F
UfokxUKMyS+PrDnW8XdW032pLVO/i9IA91Ujh2dgkaI6QcJ2rCKtRZx51/jMRSRaNxDPKk6DrQw1
lbfKYHrEaQvZ/Dgbd7YLCnN3AigLInOSKMcaDS1Um2GYUaSi/TnJ+3pq4A5zQmrHhLbhlFjCV+gY
InzUnR7XEnxZcPVgc7Erm3qRwzLgeitaAFMDe8I7rzg9oZ/XXWYUko7M3xIPQHXvKPHmDprDU2Ou
s0vvA4G1TM8y0zBrw4X6Bu8X2/eospTiuT+gCcQareVexLnMCAXUsX99WBh7ZfQZRG4Rgz1AOP+B
8Yv0Jcl0fs1RDSzQZfaCw6+nd/MgMgwt3mIXP/RkRw0QN5DmFwhFUOX+ZAu/KZvg0GdW7wqu0EZo
UfFVKc/Srn9uq51NBbwSLabwnmdQy8fcdks7GQ8xsMPAPgPEPhk3f/YELvjx2dPJrIoi99oc+qEj
5SsC9AuMvZdyvpr5LYt+EheTbdknVZcokayS7FuZ192gsixeWOT6XPiVsWuJ8AQ3OohAUVRR08Aj
1L5niPhyLljM9asSCZMk/+KsV7hMsHGFQRjpBG3ggXoXzKXzM+oAKdWiyxwbqlcvMfbU6GWOA0C1
HfMbBwVzXXuXtDR7J8eyc1fNWjeoFxnDM8AtC9WaRjOB7tWoZBQBLpmu1sRtz48MwY6PPVm+vKeV
QZgyvmsZiwhgEwqenxyxWTkFPApKT5u0ANy9E138w859wgt91wW7gdHYOuOjhHU8wZJzCuuuCMVm
ivBFIk4hSB0d8Sed6J1RWp1ITiZOHydvmLapmqrIZ8t+MjfX0QTbjQoCFG3s2XgB7jJa32qxmpoJ
/SjJAN5YtcLpsQGcm4c7OV2zcZnFyJ2EW849Ldc+hbVKjp26m/hzdIy9JKJrUvcOJb5QCneY3RpE
9u1uQlmeHtx0dA0vwzppZwqq6KZkmOh8UGxRAUHIHwZ5HKurGDeornAXbWjcBMM4vjmwe247qQI0
5OSpcYM/1OLHCd+UZsGRXPwr/4DwQRY7woVcIc6XRdTXImgNGvMou+LJXJt4qp+6mZSaJfvnCuh/
mJtQEK0PuYFBuxLePWy6OD9bSXB87pLpuif+kbEXfLVk+6rz2mG2e09G5grQnQ1fQhWCBJ3sHQc+
+zEN3mev9lqSK7BzohIgzXqU9vV+hWzx0qzINOxkLskqN2v+G9znoWWwcgMDY3/Ty1+IZ7/eIpVu
Allm5EaxP5ZVnU8FuvqraNlHTfxSKTynavyjC/DHFNB+O1S9CCcKRivH8LMPIzlAtaeSJlTBf8jE
0pifRaRWrzBGAHmj5/x7HmJpv4+LcHPfQyZgakqO90hggwzxegYJ3b9e/bAjMv3xKMg4QlIHspkD
K0+B5W64Xc5s65c0mQL4WTpzPmSzY9MlJmdFSgj/qBJ937kvgDRnATzm6kyN/tpRGK/+zfRy9ypJ
w8W6nWJz/8CWRULGFsV/BnLNDa5REcFTwf6bfgPFoDiGWvvZ2tKSXms9xv6qcpGdmTcLWjt9EynV
rve1BNH6X+SC/DcidBjw2HacyFkxLly3H+i6Vu4t1FbtcrFrdNnyWMH/T3vHh9Mp9yav32iYv+aI
ZZc3+KG2k5zunxyhyl+nu/sgT7bBfIX/D46Aofk8sYy3EdKpYDxQmexXAffVoZzsMThepd8qgKzc
0T8Wd0J8viLkFRwc40znug1ju7U1e/MgyejtPBqeJpl1ilY2j53ebvEJGlYTSb/E7GL1ABE05nnh
Wk4eJ0Kv1SDcZpZWw1fx864gJVXPLFlZiETa+81K/z96kny3gcN0QPryA/lE2U8mg1Lguk1mAbnN
L2y5ovCUpMPh5LM4wLc1qZWqtCTo8igSs2VmbwnHrPdEDuMd9gxsJBRRnU2JSaFFk7knJPr2GV50
uf0FVXfTvvwfHHmP5r7NDRqnTgdczZONVkf6Xm0hfbtxG1l9vx1jDlSra/b9bl39yhRjFCdnI07u
y7vZAyvOzKzCoAQNNjUJMegvnizrLe5pRitnqLJLXa5JXJZ//w4poSL+JyWoOLcnpjZASdjulq/T
+8UfZP/Q3/uXVfwujXI7GnRWltCJGGpyq0mMTN+U/3eDfwF8E3NXWbVPNHxPpa46mx0h2j0RSyF2
Rqq1zd/w+dKFG8RBhBwFbR7E3NeufAXkea+gb1jGZ4Xb1ixaM8bYZwH0Wc9WildPxQUqum/hF0tI
PT0x72m9zL0bNcSZX/jZ6lxhxGonFa7S57yzSE0DRVuLYU50SNROUkGwEU0hq87f/pGo7CtgAiF/
ZVZiTsqhFpJXDfYOitEPXLi6DUt49zDD7RCnhXtAYSWM7PNLW5OAI6/KBDDEQLLl5x+DEeWurSM5
PYoQ7+d/YxuNfiYEkfTOFbJ/SnxCmmdXRqJrElJn/ZCr3zvEE7Pt5s6X11xNYu1YXiouZOOgidNz
37b69eAuhp2CEE8uG/t2ZJVxnxGzWm17DRnDOMAZcXm9qXsxqz/03LZLOtiKCxqB6Ql9XsJnHm51
uhQ3j27SZQD6U5TLlUIhKKuIVA25+PIhE6nWeA14JmesDmkv1MUESVGKnCQB+1b+XIRnBJpW2Bcb
Ox48WhW64Yiw3gwf719LbIsF8cszqz2UQ+9mCXD7aeUtOGrKOjBIzbfz3QIivxSUnfhEvoUsrVPB
OqHUy2HYLB0b5DX2ShFK4zbeBvgnBsHRd0UFXa7a/H6tv4GOXoW2rF0nugTUjPl/uZOotO0aWMDU
YgIR6Q7y3as6WszAEC0OexpynRekItzqdU7rDclvygUk+2KGHQewqrdbHcMTo0gCQl6uQiZ5i8iK
26spr4kfvEFE6Ga3SzcahT62vAsWe84DcQvBS0zo3rHOLmqdQa6ZpOas8O9txtbzczu5vpvgFH+U
E11Qjhgu2nZuzelzqCQc5SaMP7oXROhPBvn5yIKMA/xx2Y46stAPzncfzTH4yA4b1voH9gqvE0eU
aoICfJxB22ThENEi6pgA5+y0bpRFASwiKduGw8X2Xm3XxO2IHMoRO0/FwNcp/rZu+t8T7BNbAlvB
x1+ZXzf3AxGkay+6QVlC49RHI5jB+q60Wt+BdEsOPHzGgFXU3DY6GQIekM219bHqa96Stoh9y9fC
GHLf4SMafb2m18lXuyvx3momD80JsoS/NqzjbsMxU75iJIT60X9prrwBw9sUGFYTOEDe9fGqiIfo
qq8YZJh1LNcO3SlGPAj8x4WFtRjkyx2h5NzrOEecsDL3Si+6MlcOxO7Cpt5mnWWhDfME4bmMA7oM
ye/51I8FGbaQ9iRtse8SQdj5SKFCKPHL+JAFZ8ozpeYOLejrYrL1pPFTcwG/Yo+mE4JPNcioczCz
TESUt4x2wXbWEgw7cNhYGU2V04Lo2/tWfvRY5tVNfOQjeOY3+m5dVNrFhSFx/0T8NhvZklWoLXnb
nWAA7HhRnlK0bAlJYeCfWGaeE1lkPyWkhodNIiGDQgN4YId3Fu7nNX5f69iiRzR5WpHKzM3mU8XI
txkJZ7U85Hgi8g5pK7kWiK0Fz5XB6TZFD7/1EOwzqVzWWpb4fs8guflx5QTb9l4EAhjkInG13UBB
P/LrtyITkNtv8zq+PaxWc/up/yH9oCTY2z0vlHsINsKt/VmvfRC3F1I+HAvbxj20gdTwLwFQ1jpU
aIM4ECJKKtrauwRKyxWCqgdPskWEFK0N4JsWsKEpAqQdK0BHIFv24NpjVsjviMBhbIzxiaF8Vgd0
7Dzi5ZAyidFW0kGmAlEin/4/ExbhQDQJDXzBizXjhWnmgkrcXUBjc4qIyfM6pZQU6zEpeh7Fubqc
H+p7zQfQ7eCVKjDQkdBNppNsgEcRXxothBTCQ6vjCRbIf6/8eu2c8VmOFvq1HSvFWasHdWuHuFDO
t/OtFcEfnfOldP7Hx8gGYEHjbBK3k+Cnv7u2BY14GfE12Gu2WwnP2oqErGZigN6g/0lw1PqGygV0
t8hzHCAAU/9yuiMAZnoS7HRaB5m4hWAeRgSA2zkm8KejnWHs9YYQQApMRQhvuwxWv/9+GfZtEdXR
vByNSdoOm0d6VEQY+GT+orPZI7qzOqISfwVIpSnKykTZ+rCkZYtYmgdGOz8zjFSozjFXCtv6nnx9
qLrQBZv53nvP3MGKHd92TORe5G1fqVgqYb55+Iq+lwJtda9x9SRUtXoTBjr6Cq3PgOj1Dhv1ZQE0
n0vh8580ABG5/ISsvhF/i3BWTtJ6wDURisu+SVZBAIxRk/otbJiOnnLFeBx7u+MdIZh0MzN3bauA
qeH/2hPca++WvtmvF2BbLGNAPpnLNnZ4KPFnJOhbXdVLckJUsnTaVGIBI1vwq0qzMcWV/frOagKA
WpTbvcGNIH2XONISKYunUBG9av4s7EXQa/UgPy3xuUj73/906o1xW+NPK84bnu+hv06rokqjSwY8
PFyg1voSZ1xZHk1VB9M320D1VU710KG+n2MFtf6+lCXOAx4pg/bb+aBQy4Sdc1JgaeGLL/oQRgHx
CEBJS0N9wQleMiu5aPKDWu4KVyfVDK7FrS/QuUSrFHMTUhcwC7N4kiv4QuUSAlQ/1/jUEsxbo5Ne
r1NxpNDGTUFGN6ikTHvWxtLrhLeYIUjkeEVeD9WGFjrI5xOSkomAalfhEBz3eZ7jMUuhnh28FYac
YbTzFTQEy1dSaHcvs7I8rDgi9uFDDdmjY9dStfJW20+48aq5V+6ra9izoFIMvPnNT4ULWdIpvshZ
dQrtOIvqrcYNfcBtHOD+WCOi7q+1pusAucRzBJXh7D4zDJQML6586Os6I5KbPRbQnyt7pao2u59p
wwxSXGzfJWnqtOSfAsMozL7o3Sk3vHi39paY4rGbqPFBxTbLAR+VeQL97C3ZZw6I4fdRWtJviSkx
95Fxjb0O/vooE1GPp1VlO1pPQod3AtBlEkMZqBwMDfQugL9Kc4Twcnr2WMPP920DZC7U8uOOQZdz
bqX4a7wb55BDTxnLEzBn4YK0HgvK/z79xKvunyFdRLbRbKKUZFthMWDM+3SpPmQgiHm+twS5RCxa
5zAYMcqn9phEHFFoFT7WaFv/q0sUutxcNv2CCml0vDiakyhayGftyE6NbqxZgwj/Idnc2zHrpsQB
ukig31HOZYEb/ibCiqgOAdEQxJKdh1V9P2tzQa/Ar4ApyBracNjaDWfUr4+talxgd+clXbg66VRg
zT8/mvsAlPSLzu9sg4l0M1KSUtxoWXBV0egL4b6z2xLpT+FxyLHexs0Tm7l0X/4TWx1W1kVB7aml
55i/UocP2De+d55ainXZlLx1WXcNwbmmymFW8g4QHWD3wEbrjpdxWMLV65hv1r2h9TYyi+fIy9QY
PN4ArbBzDN2hF5uaL9gKiv4NuHjpAVqqP7RiW0NZ66k83xsf4vPYXP8Czj7z2xIoliXLh2JkgxUu
miCFOsWRVjjRDBdDue/osCP9c9t0mHZlJqOLM46lqWzqa8fxDtkMDjP+g0soRo/P9i4KIOt1PMnC
YoEdVebek7d6kwAgtoQj3xdnq5mkXfnK+W8YX0/5wNpMr3A+fIfihn86+rc1kwOAFCtZE3BAubW5
UC8rFRXEO5cX6OkzE0NGDPhYr07RPVhFhPgJLahPTBHbrt7gLESFovqhOTOHFai0IE4mX/GqcNeo
B6QZIi1dr+34qqREUj/mBtB1xvZ5jCj5pUhBeQZtw2DNO42e+h9EZQhITRnJnrzbUaTQ4EIoZemw
ipID0W7aHEX9xAsK8cioKGyofeLxba1srpBZCABgh2XSMMh3uygsFKDvLJxj2DE4XbdREYmg1HVz
TCIVqFQlyezYcX2V2YtLHS8OrnslBdGj4dH+fPLxNt2qGW89qTt9/KI7R/KLpT67MwfdEyRMkXw+
EfFWayv79VOo0gXmq+Kg7rn0jy9ABOAojVe+QB3aqUd1OkkBTdY8AN6KObe0Ja16ukdeU9L8gPaV
7FKqKzrq0MayPzlQl1zhzeXXB1+wT9mCOGPeWKPHn/C/QUxYzNZA+tp2yjcrMQvFHa3XsaACqVUA
jrJHlPj2KhKFbHCDSbYADiOQi1B24VICgqs05+iaHGf6xi5vlBXEHWkluxsU53OUqbEme37nVA1J
mbo6lrkTqC/v0l+1vjdZskdLkojaXNTTet9/KMeD9p9Dg0me9eknxlnH6Nf/fsrOWTlMLBGXNdEK
LKRLtrJxRJtCLaM8Hl1VEKDPUTqgUbFYIEUUQSbM0mVkHSh5Bj+2MYuX/w8DNEmK7FF/GpdBZFO+
XwT0gORd8qsFrhKANSdpwnpbvhlhGB0GvfbWYrD7719hYJ+JEPGvACWqFfNJtDLSQxjc0xgpFd4H
RQouDyLKYqZ1SKfVCDpvP3PQZaLeddgwjjLKTrGjseW9kvQjsh6cLHOn7QO3nS5m95BViVUOfCjv
P2bw60eAdIC280QBl/AZm+l4QH6AjkciCz4FLxnZ6B871d8ETSImMEAHq/l9eyfQLxGqNs1tSj/X
+qkP6GW0tUoGVKo1eaaMWFtlCoPTJRXz9tcKNyBCF5d8NUgQht4CYSP+DAGfDCkVxgDVkxZHI5JI
B3LbbzR7IAz6kmVD/W3bK4NmNXN/HE4omIAOaVhh0aK1ee9S9v39wDz7bAr//ZZe5H+Nu0Oyme+J
IbdsWVYFw1UhePJ+9fndSV7ZVnWnU+zO4N70tP9Bb3uG5mvWu4hVvGLneojbwTSYXQcxoKnSmxuP
mLGQs7pzi7xm7wnBJxIIDXZVicExfEQAJ4vCx//Ygpks/EjOg4fxXV2c+0nt4CNiiMAkYti4ZPnQ
WNwbh3s5k6othk1KigGF4PaCSZ36n5KYlAcmBoEqSp/N8CGPjor2Ja4S01warGIZmLg0vXeYSy0S
V2qercpeF9H4X9nNb3MKYI87gkxVOPTB+l6oKeAHl/S2Z/gCXHmrEeGPAMKTbVuXiCWMFrzNbW8O
o+6onztIIS6Ffdkj2Ww0tUd2rT9Cw/NiZHruRQomOh7aYtvR8BlwZkXopjZRwx9C1bMF0gfG6zuG
W4murpTA3w7XiVVqUxvSMr39Zo8A6OWoQTsVJuVcyoEP5cKvJ7D0USYHtlvEPEB6FgwdNKqZobsq
e8S482H26dJX2u22+HdV86i0pr/Px8fVv2NjCI+F4b7uDGfpr7APjwUOZ/wY1Kez+kWWicEhpq3H
2buVm0byUDD8Ni01osO4i6dXZbRSq/K5iKn0vBzXz+mZZgcHgvX5zvui+KXOqKYvcZ78MQ8flfpy
1DoyxIz7ZsXII0WqsSocCs0bsCXOw/9LkJvxrqIhFZF/qZc6XeGz02glqaT5P3eWp512liiVGMH0
ZFLF+XM45o9KCTgk2R6uUENEbw5uk0KKuK6XyORB41RgFMlAcav5nuzaXAD+5iZHm95KkBWiWJku
Q8gDbqu1JdNX1y7F87uouXiv8wqVex8L/DNJKQGO8s7cQnqwE+yXLUqpB+ui6C8jlmzczaTSfzEX
BcyiWsPReuIqE6DuJaNwaSChh1I0exJ4+8C/tgcoSGqPNfh+BDHSxUVceiGnM98TXuXKD+GKuChu
GK+dri6EAELkKcK+ZvCRfp09ld2p7M42Ys4gVuPax/SQcbTlLEAWc3cx2SGTecjhCBLohWuJhHfX
cxrv1N9Odd3xip6nYP3H8Moukb0FUkIsO7i3azNKLaSLIWCA2FRgKYYWg9Q0OvUXkFZcQJj9z8N1
OLH4Jt1KwnyrJa36E1J7TKfBQQJoMgCMRDfUOV22RuCtM156NP2MmygRlSYbXySStS7UvxTeipT8
k7JJJbB8VBpBZWJ1yd6SiAgVX5SR+bhgSuLUvo2AniisnWp+dL4hxf/czH3r4JfnQOC1+TJlY1Yg
SWHRJZaCLyHakt8YRuQ9rdNkghgtvaf2jNZhZyH6q5Cti47HRAIVEcuds3bN4vLFV7CiG/SLExvj
flFF90BIdXdGvCXgzU7LtsGQ1/gvq1v/9nSWsbXonS6BfbJ5FP74Odshx+izl92/AuJ+SVVTCmnO
dTKHXmFx99AWLQzhhe0pxOrHO7lyHlbI82ZMeTeSx47bZBt1GmKIGQzP8HTwqz1moicj//iAnrZS
P+96rKSIoINtC3VXmNqPXIZwaAZjCINYBiO4b9LPRNcyqRSa5G6iaV8PiDd/O3S0U9oNmNjfJWLP
a7WASWKN2Lq96ym8T3cVAbHGOrS3rpaBOglTi9AoM9xNKOC2du0cP0frTTjOwZg3GQ8Cq1p6wkgr
nkTzoWUeAMEY3OeJLIGZq2+rkeUhBma+3KwFz7tJ3N1yU9upUD8TE6+l4jfWG9txvIckTfnZnoT6
WRl5Hizq5OPe+6XaQ3nJId6aJwpKv5hOeeAPrFOqvCjfSCNAgMPB70gkRjA6CXRcRfpQ5/ph6gRG
5xMAYii9OYE0LH8pAtLZUPdvYRiE9A8lhOmLvkWUO9kLNW/8wstShs1gKkqmvXSIegPcibjvG8O+
8a8ZyWHh37LbGhFQxA2IYs84gZCFOgvDzAGUkQGfh+Mbuoit9vXBNV2IWuYdYTfaTxuIAulHkZL+
q3lFPTwQIpwh7Dho1OTQlhMqnULuPx/+YB0kVSti2Tt0yAHVCJhfq0+djolSFSwbmRF9WfCV2r7S
9Uy1w0BAJvWIQVLsYzQFFE9+Fy2sVqAR2mgv1fD660CCRe7BCzOg19idqVgu9Z0TwM9eZGrzdmyM
ZxOiKeOlpOHWve1SU44K4VtC6OvWcJxla53gqkKbWJbrOaeVY7EgGjB7tGOZzz552H7C0o7d/+Rs
cueBIUcJVi4E2Xu4lFwHBvO3fUKTHxcdosADiy/SE/yJ2vEb7T3qho4lCpPiRyEip0e3K5FwXIYk
if8ovxUiqqFiUBxV0wUSN2P0KSRhEsDbC+HwXt3LvOXk7v8zXmpdTWmwCudYfQi4J3fz9JnnBFM+
swQi+OTd9oepg6OS6mUcOS5JPEpuQSIaljbV5pqjfGjfLZrmMqK4F+Bw9ey1Z8hM9ABIa/YJMesj
wx0hhQz/QqIt7hUTE5/w0ZY8hIEHVF4uW3CbmJ9nOflKCQ/1n2JHEV92yRCFO9K3d5fYIWGa0IUU
3SXTGDuF2IBfIpi6v1n4LZKNs9PrgMKVhsOfAnMxkfL8dDYJo5fbYHFLjmMARYHte6jc1ztpKjEv
6FOS6RTaDxsHh+0+k+rJLMEndA/R9XyY+lin49JRDG8u/rJTlOUE8bkLY0u/ZX1Nq0Ll+hfWCeHu
mtEFj9ze8Y9e7MgRMGwhRRzD/pwvWEP2FJ93yHWEA2YNNNdwjjdXS7NGd5m+hdbuaOwMryok73dE
ju5WP9SjIpp8qj1e8GMqdBPoWNhbcRE8Tgf/5rmNMg/18dN0rlb7EVCtBgFed3fj1EcsVH9gjTXH
8SsB2W6RLov7xx8tPxSmIMnk902k50bj3rbkzpWqPU5Z5ILEqOH8MTtmSvFtmKdB90dPImF+ML2c
sIHfedQaMQuOv2Fcr2uFoAI4YJ9kkduCQxiBmo/HFHp/N4OBpeECnAmMjA5YItTN7R4hCTwPs4M3
hLZopPL6Vhp7KbnnTTbVxx5M6FcuRWkuGLAm3eK/EHCArGHm4ON7GQK6OtPuwOjmqThY1PD2JW00
rNcBsUxTpWlb8hJB80C8bsYzN/pUgpijc2WAoyXooeAqb2KdhCD64uqdwPy4hLuRKydd+CAfsuEM
xfoquB0Tva1xzSUcvgJ+NfciuduQrhtiZd9ohNsFlmkWJlFqqO+SddQXJudz9AQFBcVKCBg4A+kQ
0d+iHV1HRHjP51CoILM2pG3DhwUK9YzT+8cTco/LXums0G/iyMt1WIen14hlpE8lsw76tcsY6Y9K
lHlvIedb3p1nGM8Wn5jy8eM+zzQkqgHL5CfLdh1TcMnpYdhyv3uIh0HCrTMm6r0/5M4KUhCCBwh8
rCw7nAZmMvTDtwuEZvT/cdJDQuihry6aIMemXzMs9K8rG1UW3h1NMcPnNQ46ggms6jrrlQM6zFHT
tIP0VG6etsHhoeVApFd7lSxm3/Ayx795W3Z2aaXDgEP49GJryvE3Td9wxbFDVTozTO3NgiEtNejw
RkDooCbkX+0+GFo83Tj2ROyAK+oj/f2ZmWVqiZPREZffQaADdqxR7nq+v0lGG3yCSo3Gal5laQ2T
l8Z842tmcLnB2+jpcLizxA9JLcdeGAqlldR4EdDOhszocNmfzxwQhCxz2vIeu7OZ8N30V2rF9q6l
US4ueqv714C3pdCciBgwcq35jKi4NNqQ3W3HKxxjE53YSc4+lZWJWwB1SoX3dZcvOI3Lk5CGMR5a
5dxwyCeOirqeyHswWCyUz30rWV6ithXWQPT0JdBAB/HzdmhyCVnjpNB791FyPa9C5qdKOWrn0GLb
PN0eZzJto39WjrY93J2tNOFJduYPaf9Z3WbXs9bPOTpvN+IMj1j5uiWkHlaGsTVuTEMNg1IoSRKr
e+9BFg7IFR8Nnxtifi7EXd0lhZBBuTU9FHLhDcd8VUiT/RzZYGeEQMcLQyMPZhOrnpoSGpJfasIe
3LRQUWlq9FXEa7O/iHqXmpWHvx3GWc4pojshs9xVe4Pvu2eb4QbmbD7nk4B4w7WNFrDEumThEQhw
ozv34dD/3DiMSscMqLl+s45RdP22kgadskZVbiDdkd012cPiWzZM3IihP3ZCfgCQ7JZPHLIR/2i6
lIyJVm5hBhvOg5EzZj0VdTDCqRM2FObWqfukzlYuZjD6/Vm0GlXQJeCUc8zXZSxGVIZ8CYR/Ztsl
xHutc/KI5tCmaGMQ4WQ2o6KfA6/IwbwZUcGoyfT6+aT35IZtstF9zG3m1Zo/kqangsJogfgHXro5
ojbLqfJRfr3s9lVmB5wgKUy1rydhOZIykzxA0AfTcZCm8lYRXqAKbaBJmG1CGp5hAGwaFjKICeU5
iEDQv4mSQetuOAIXDp2+bwHeNGrHa98ywGVB2563qVCf6sk16gNiFp92ykekmeIGl+wdODRjliT5
TfVaWJDDRAWC3zoNlSvRyMfkb0VaGm0qGvTfudd1DhsvvwxjcBF3qc7JYzUV8w5ZAqOvJq7UyaWW
j/bDM+6UaEk7pnX58Y4A7AyYbLbmLrUn4UHARCGHe/kwPSfKTMBjP+Q5puUE1oRvj6oFNWiOX/8h
Qwk7+5dbPRWCwJNdS72npBUzBQfAOkaYyPlikhYDlKwavgK1BKLVDR/13DnNbQc1Y/09IpI1CvDb
nFxuCAx0Alfv0erl97GRXqyYwN4UTeGnqpO8Hi4LFYit64hNRWIr4PSGQN38JmqMHVKXKwmovYiO
C9/mH9qEMM9US4NUFDTiWSYIIfEEZ8SvKmbLv+nRxB77Gt9LJR97sCL6Gry4Cts/lr7nSxGlpSkW
cUUXZrzOoGL+QPjBUEC0b1BnRx6R4xk7x7aaKE5/19FwCOfw6aozzFyqnmWwrLWdbfaYwowT2T8J
ca5zkaYPmpGI2QpxXpUAe7KkOg+R/KmuBnrRCiCN0c2zLrIYUK713/bn9xYXkh2VfMz7iz6pSGhN
ZuqNhAUtSfco7bAHqeXEm4PRmRmmyVbJ5iXIAQB2lvgS7lHCDvHQ0ftaStHFgjo6uUUHDMxsJ6oS
DPHDs+DGQxHV3DVvkk4AW8aXgVy3rUfrL+jyaszvFZvOjwTP+wqkzkeJePZT5gCg3uEebZMx+Kz9
q9K0eub6zPS4Ja6lydhag/2dBrIsO3PtF9Gr/HwRvY2Y3qw3thK4gHeBs8fBN2QyXOOx48aS0MI9
2XXhlqURtneKCxp0uJOGRmW3kAg/GON/ar/Y4jcz9eDno2NVv79bZlmWrFGp8jP3wi2JOK3+G/eB
bUYvZ1Ccg+q5hq6fWz2lkYpPe2YKFpZFfwxR14iNEot50c3eM83MihKIH/lruyDXWxbiokOsJNrU
zgx/eXUEmeD3tjExEiRpmUggGijXzUoH7+K7HQo+zsPRK7zMHmCU+nJXJ52AUat6cFMNP30JX+mx
oZHFO4rOK8dqoeaLx1j4MooMSP7kgqstMkdTlCslSizmoaehSs98mymz4QVdMRcIIFZYMFyKERRO
CnbjSbZ/owU+tAWsAS4+JZ8tXF/sPC3DBpRNOMhc32Qb51fCZF7/IUh8bpC1QDo8yXzh9nbfuPFw
DiAjd36ISIuB9ktcKsxZL7PB5lgNiK1vbNa6EfK5AbxSkqY2lYePwHYBwnLFqDXSxOamz3E0LGgy
WiEvu/fzxf/9ZDLHehPz6SaSU8G2/XiFmpNTx0r8EfHqA7FJGJkyaoZNQ4agENMqr2ajaEsKap7G
B27dmUcA1EnEKNoHzvalH9E7X+krwLvCgot9G9uoxpsbAPkAWwKMjwa0LjBIAXm5NuzmJDExgtkE
KMKYUuUVtRvYoEbbVuJbToDf8yHbuHLZM3qqUTzQ5+tW5qfIsBPesmU7zpM+FLR2xkc7VecwjAD3
ozYM2Cekp/lMmlwvazrdywi6/AJEOIIPX6ONZ7eOoEunR9mF/v6BvyhrvUsK3q9XATlgD0xVxcDw
rMIheyLjAv81WABSwc1oVwECtMtunkCI0hJefMogz2x7JRsGZQPPOkHvEKof5Z3UHBg+QwXoc8e5
YTRgmMHWLNcStmgPOt3ut+U8T8hVGgFMSJzCwTJ9pgetm905Gprn2tqj8uU1W/+uFUKyupCxg1y3
+0py8UprKFjTu+wsFAdCz17VQWPKs7+OvQE/ovgjVg5chOGgwFIB8BcvdUOnEelDikfvFDtzf5st
O3MXokfR5bqagDJ7LiWoRS4/hR7SNoTES7zxG5jBdioLq/qivscYUVaWYcw7qHg1eKVRxw//K11u
k5hjcqXDD057pDn0EdsgHvfftZr0M8MZ5Y5hvJ0HevK9gxfiwFoFUPLM6Ew7/mivMpFU4QOaCTmb
KUsbr/zFdMoh+UjDTqyr+MSqdMg2wx8nm+LPPU2ONEfqxcNYtw4wWKl8Y6VTP2ZhfXjCGawllnMl
m1C94Ne8/OMbF3KMbO3TPwWLAm//a9t9wjsWbnx4RWjaeqyiEjiTHMCVQSMlOBlTT8+sf63nJE+k
j7y4F/XKEOudMItJkazPEHuz6FAvy8hIeGIWuM5hwFu39epkgUOTSRdQOVZIykaC87K7Y43DI+5T
tkZsYH4lkHEAeOjew8sl3XnRYjtnw2kcCiQKI/e4/UNyufUYP2e+UsCvzxBj43j8XN4xoEw2Bzyh
0shHl2nz5eY3BGTRncVyReP2EeVx4ujZraHXnVDrDSt+pjpWbsdd3ykIwlnRdva1OpLkB4JsxfCV
fz7wylCODkGTcRTrrfqOxc5btuTjKd3bRsT85ysn71N1YVgxZvZMeHCzbd981oiQYU3PN6psbdgy
EOOKKA5qhNfGeZRYTY6tXTBoH2ghrj1Eo8lris2GqUi2dF2CYeULeeVwYOizg2I3px+sCh65X2SS
Kbph6/zwI/UzT7EvXBj4wm+2P6/gYMsSOJGfsu382C8L+s8spf9hU1ZlHdL2SWPefQ3dBAzgEo8i
yih1qmFBKwvVKSM5647nKa6iC1bqNzMfo98NUEPaPAO5JUCYHbT7FVO4reF84KDsKAHoyY0/AuQF
tV7OTq1SMiW0J3zxqiQ0fkBuZhUjlebvKVfp0Yt/C7eAC+0DRayDyy/X9SmBls/2Kfr0nEuXroB3
SgkDJRQ6SVKLruNI0jQctSjMw7qP+34anuXblpJxWwjSQ+MkV5QazaEQ3GuV4yHQTa0tD7arXVp9
OQs7DKwEk3evAPkQr2IZIM3GPtRdMFEKczgxZC8Qn143ykDobS/BrtYOKDQAJS+Ny/ja1tyWyMM2
VUnuuFNsxAnWSwvqLqj2praBMDvXT42tVpBD8/HiuWJc7GSp5OuC2Om7qugQ0wvkoWVzQN2OfZkj
IeTnzHscYBTUrRDnKbOKwBycnWzNejFDBjvAwccN6SeIPR4tM3CJ/1J9/J3cdGkA59h9rJ3yMbn+
JzpxgIxaGdvdZO2cDkQa0hQg/ofLV0NTlRG8nyQWPOkv9Yz6ygVSPc4Zb97z3yYYdeMC/MN63y0E
P1SGqDggilMFqwVKoMf4ar+sUvrYjLfZSn/ASG3A4Q8IX2fv96JT7Buu93agq1gqM7vAViPEjinH
FF6Uut7ocs+ZI3Jw3s2bmjYcwxMi8wmSZK4yH0QokoMMZNXvGxhZHGj743Fe3aQP+B5BIChDKtCf
GNRjTKCmSILCTHJTFQLJCB0UyNNkR5UCtQrXe+vmSKKEGHKX8KOl9uOY/5vrms9xYJyR3KqB91kS
CAqbgQ0Qwim9wq4/fq5lUZH6t2GER0uhW4hXxJEgEC0sLgzBBzYX3J9aYaqpJSquvwgIZAW1eHQB
5hib4TxJIPUi4eNTiO/vczQNoJhIeF8M92DmVTEAuCc2YVrY7YO9iaOmNRBV/OuPhdJ/C4+b1niI
AgokcWyJnmOn6OKu/CTR0EGV5LPKllvzk2wcbl7CdQonlu4DM79lE6e58FLLttmEUoddqJMAk/I9
A69HaT6dcngokTkFA5TfogGMl8aqpUQjagJJXf/se1VLMLa2vVUKEWsDt7Ye/+LUj5Z0gGGZl96u
Sn3HeRcEpp9foaA/30B/93+3BKli76CTvqFNb5llCU+5ADjXKi1QnxhzCmVzWThFAcL0pv6VhPmo
xVrMgMMvjC9bUPg3PSerzrLmAQXBKbhBFsvQTanAZn5R4EIcgkPgPvDEXOSFtcE6rFXJQ0d2iKTF
Yc+ywn42Lv4xcrbUS+2v2TwL+1Vh5lXDne21b6Cx1CWC3p6fwO8BsQDCJs+dvojIfrIl/pT8iHlO
LMScHLzzvxVjoQuRW/rFeME7AMnvwQatlNw+v0Xoz2SJqEP/nbgYC0DYSEa/Au8bvvB9RGWqEO6b
4ZSWYhU131plC2soZnEJHMy6+P5fOwyqF8N4eRoeRJxfpJQX/jHgpZfhoKIp6Z3TWa3uxjZjbjsQ
R4zFCGJBD9bgoUFZDQyqsQSLBqEVyjJmFmhXoMEK2nPnTfZblYYPlYSXFC8q4IQAfqPu+iilQmvU
lEquecDqT3t7Ecmynrh7y07VB+6pfMwqviiDp0crH3/R+xWrV8Riwg9XFEkf3ZNmESDg8hK+690r
o/xQLTKPZzzIbMqEZYF0rbhOZCkRP8/ViEfvk/tzMdjbFhKAAJgd9k015k/9zfIjJraM+S0QSqee
VFZYUuVdgu865Xcks44Oj5pG0IpGIMY4yiOlEzmaumuBZ0hZ0q4szpRvOAbZ7DBIi9D/WOVj1205
iewtntj01Y3vFXuynufHCOvXC39DQtOcTj8mSemRk4NVDayc9BposNxs9SOOHeGHyoopUdhYSHQb
dIeKHMML/YXi7NcyPpPG5NvA7mbAAhFSWON5p0D3HSXo4Bk91Ip0aduxgFus+VzwhHJJkGGFKrba
58Hdo7dQ61c6pb/RoDjn4N6o6hJZH7/UtWQbQlL5S3A5QfPydhSO/VacV3wyCwgZDuKjbBoQ5eTb
fU38fRsEMJiV9g17J9mVrNEjMh2kaMg4ypZ8agC7jb5SkhFN865ENW75gwCySmhtcmJpAtdM5gAb
FyXTDyDKlpsfSneet7pTwVSnfRdujN/ZvDb0UwXUYw/t5mQelgPXaIIHG9u21FfyWWO/r9QGrZlX
G9HOVf5+ccEkYfzZZ8BoC8h9n/teAaTFn/lTGA0WjykG3idgg32TIPCoDv8JOXzug04kacATUQRF
G/En3x2yyMxjjlNGTO62oR97LJwAR7gGoOsq5jUd8BZvY/XAPKCEYgeE7TIjcv/a0zbNG2Nt7418
P88LkcLsEQ9tCKpGH4yFFpOscn+hb85so3xxK7YJ4JZa3oJgaD8Ms+ESXn/2CUpZzpJfdYuBCmre
Hr0PExbg2ID6V2WPVZdcKHurJklll6KoKSlsnNYp7SXZ6oUyluKVqp6QUQMPoXTPMnYKMj+1oTQC
x7kt5VxXN3KAPdOmhIFeX07XajYkqZHDqC4sZC0X9fajY3yrYpNwrjaomXboZByKNIZVtVDZWRcY
rqYGDW5lJVEUDVCCnhwOvzIswqrdAalTLp2stkb+aDBXtGNEVS4LZ1WelbMHXr2sZ/kVIPgmnxmd
CmumEHQWxNMZi8orlZt9W5Ky9e33FL7WPw0okcXVebaJyyQiYNWD7IJbkoDdOdFwjO60PpO+SghR
RMXnH+wnmyBQm3M4BxwDhq9Fp56s9gt1jxFUyIvMOHhA6qhlSIxUDQOhNDTP0FjoAJqv4gwoq+fi
gsAf/CEZomWUpJJAr6I1T2TKPg3By+qVzzMoIKY+6081o913/c1FGId5wOWWqUMHQxrmVH3nakTz
l6OzbLyTunIVAI0cHOzypXd3QwzqzX/Dw0KGjc4nBHJcoC5V1WR38+w352KXDjnz4xD63luF06Zb
EFe7WNCjcY9+V2d3dcN63BCHsY8ypHIx3dTIirhf7Jwp2y7curafz6qcrfsqMGuclmNPjo4n52s3
FUd2igeisn9U2PPJZduLCw/qlFO0aZs2IyXAm7SFGuZIy5NvGggBP+0YgA4Q2KYdsFelLBwLit7e
hV9rrY6QIrlUUlW/DzNwqtt6MUZUcGrkv7imeGmHm8/5M5XCffDmGZnCwH1ULmeusArlGlBQMFe2
7TMqftbxlMbqjVYT0aFbtJgxsyqZ/zfoY8xp+ICBMIeXOZG7HpgrjDoXMj5NRBPyQjOvWKJHyRFd
Y0zZrRCvGOcFE2BzlEK4TFSj81PYhP/Fbmu6D9n4bgYEX12h8Y0WEu2AGGFPTNEgYWq9Vu57EOeh
OIeVYzrOZ7yn146vR1kAEruf4VC1YMbVTSZDqx8emAyyrsXk+9/5QooHSk9Ntx97XIva/BqiaHQo
vIEWBYjHaj28SN3heTcJE+EwRCw8WhMWYJr4TwTawVtOQy02iqEsT6AJpQxsKRu0klwG3xL5Gnu4
p7AIU58KuvWnSGZ8eaZEaF8vBWrvPbYslTnK7eZAid5Tk5EboQUuxqT6wry93+r0h3aPTinqhgsC
2UyVoIFRkD8AP7b4MBsZgorTrr0vaigT+u0xKglZSZK1fXdujRwoZUKZPL15RfzoQWvrVtvp0bHu
/cBRozx5PKgG08l8gfRaBZNHMBFOUaXc6ohaf8BuYU6SgiVEUct7Xwp6NVGeGVtT28PAnzF8rGAy
6QZ9q9vrgTuDhGEsA1dBO5TdobPu0L5Whegv37v8ne9Qb7Zq0Y3b/yItiKdbuK7zXwcI9fsUitR/
k2P2CNxPtgVN79HXrsudImjntkJh3wIR9zw2jqScBz7JwHdzOwWYvPchOMwYvJ4ZwxwMXxAGoEBT
BAZq+zP8WvNOcpRvz9lvQgPZd+MMGaiJ6uPpCJmcrEnQtq1CYbt272Lu/5suYBmjgnvhhg4DuOoA
3ZzFDlL5LMN8DjN1LGYa5ms0grfi+X8FgInt7PDHnKXL9XXiWwjpGmZ4w1Aj7Bjz+zEMB+cx7ECe
dGipUw0bgRxETAAVsa8ozN9EnsiRDJZ7xXoVQSNuyugzichz3TTy4l0V4lgnlAy9PufTZQU5XfSx
6wY1nti+Cz+QvkpKhOUGXF1emdIuyWJe2xzRTLr6rXsDNCoiKSa5mEZl1h+vOsJBN+icHwECkOTs
j/pEaaBFRBbGJRqIssp+a4aGLfzlRfScre+yKhoVkzapmywmAXHAwKf/x+sUnkBlYlcDHJoQzs84
utT1SMQRHJ3eQuCTCDQdll7sdXmKEBj9e/ArHwYeulZaA7Ps69JxS9cd5T/bPFAcrlPsHz4u+X7K
HEwZK0CbLwFBVqW2Axb49puW+vhI6NNNGHnr+aIrHAjaGcr1hYKEd70z7c8v2efayjdb25SKNP9o
9m49Md7eIFTYua+HxauX6EJRuS7OasAJYUV2FW4Mvf9TuG0ceEaLYn2X0ErfbPRCwc9zSQZXiHre
5ajg0WK7q5DCq4O1q3UTMyqitZe7InGIeHzBHks13S91z/2aW595Y5m4ss+cEnyWkIrAsS0z4uPc
tbSrb5LS+EjJPLXRbt8pi4gHEiN2epU+buDNhNrXmjCD41+1DP6D5MDbHMwXYV9pJRkSDnI4C2cV
9tN7QjlPOpSS03i/mKC3F8OxBMDLFqRPnvkA2UrvaZhD+o0btdkeJL8Oqpg3c6TKz3zSiG1ay2sK
T48Msu4ffnv3MmvBS8dVBDuYNwB/77TVN9ZHFIOtWf71Ud1gpVP8OoHU3ONtPwIJEXhDAvGt360W
uP2ZBgAceKT0Ix58kM0n/+NHI4iuw7+n4ip0D+boUAx+LFF3VlAP9NtLyeo/STBdq0LMZ6iPRhSY
yM4IfRjSN8SElSkjzATP/J8oYuadubBRFZRrK4hBJnaz4eVV30tRpzBmEQiRGhMZ0tMKT0fHBFMK
uuKY+BMPg15tmigK7RiR4PgZaxSN4GQ78t6b+PP4EOAP5QSytFay5OqXHfyKUvz90jlj8B1WPswJ
ckAs+gKuKof/lwQv2h/DmMiilLE80PM+0b+0vpS5bx9icxZYjW4AZx+Ya2GiCxcd5ZYGrfAja9N5
frLKso5OAarRwM8CDGoLQTycWgDG0HP8Qr1XPNz9jUNBI/XYeV1pc3Jmub7KvUZgaJ5uZSAGtmfk
k/JCNHNXJlQ/4JwdRG5IMJxAW1tOE3qexgaH6tsl6knmjtQLUlyfPXYPgmG6Siag2a+OA3e/tofv
0jsX8qzsp8t58As2opR6chSvrOUnFSkm+4PIX0A+xb1IcxWEkLefzvXpd3GXqQHBsW1cMdIpmRrW
LXh+lk6/sgYJxypAKB8aYeOTLIrt1CGJc8dN3LdOw5VLk225FFsXMPLqkI9B7FjMTNIKflRp7erW
yNLDAcdXpy1AHo3QLOvi6aGwUebG25x66zA6CCj1PG7U3AgozsAm34wosflFE1/DlWw4iFwTs9UZ
AItFdmwNM/x9fvbExTsl7PJDhuyFTFdrdV/gQn6Zei2k8WOBef12r48TBC1OHp5g+7e37Wfd8IsO
h2AfwTjUl732svicv3udmpki9F/nRTYcf+KTRrsYehupJdNUcUgd8GhDbrH/phhyDSNT9Rnufufg
T9V68Q46Bnw4yRmpE+2rklEJzuZywOaImggBHicMNlv85RgfrMR1zDrUX6Ylqyh30qcezGc3at8I
+DD1j4aye2uGGJaOhFA8VhCGz+rJRDc7UxDFbREunl4MWg9c64tIuocaZhovwAfdb5kp8kg+jDCu
8OxtO+LcWTJi7jPCjsuWh9Lortz87JfbVMwypSS4UDFzsaaM+obPDKkUEnVZA3ftF5qh3vP3X9Am
gOZ5zGWO4eMxp7W6vi7sF0klk4xZIV1qg3Kd1wO8578RryY6n5EJv4btKv/bKfkzuZ/Tc+Vm/Hbs
xHgzOMwJEFT4LLCpLX47V/oEFeIMhBF+IXVVK2XGZGM8y7BcKY4mALTI0C+qHs/bUcpWb6rt/5rv
eDZbCD/d0tvxf6TEirLg6v87AETiNEaRwKxELCCmfX/P0EdgJeRpASceIyssYB5vgo0P/ZwpOfM+
VBrr51sr4QYx8ZmqbW58FKdssEaQXFof1ktjltoQR54fHb9vgvV5rCAcKDTfVmgK5Eb84seVm6gS
fYoBJNAVhMRMpoUQuVMz2JZ9MjZpMzH4Vu52ApvyQ7ODuujH2BssIlbAf+Vtbhq5hSuOFpxX0r4H
iPg+src+UanTBl/pd/ap5O/MG33iEZOstV4yPu2pDBBeQXIuBNZ0LoDda7ROLfSWlMkT9s3J+aua
CMry/JW/Bt6nCsRvkCiPiFCshLc/MG+DvzA7OUBIQQPK8QZhJWgYknWzFPfkv5KCD9oM2CCQ2PBK
/BG+b+aDNx6uiWl+QG5Pucwhi6lReWIzO8POfV35mVY3SwNgcTdsmddNSpwz8zQnCFh2+WkD8SYw
qVRt2oLaWIjPVZo0x4/PPb/AmZHZtwlnhOYqO52ScCNqmS5MHgSeb2pGAg9uXs2mjC5S5LcTMikC
2HezPUBhop2EAlhc5ohMWObL2+pvZxibHviFvToqyoNyAc+Ba95okieMYr3R0chJ3oXLUGM5T2PV
6xxY37/JBfkrCEIpArbtuz6Cwt3q3Ngwe2dLlPiyc+Pprzn0fVx6Eq+DhU+VeVRr1Jbto4nM1dE/
EzcVFNG5XwEjndHLulHLqHemkhow7oq166lsctX0yGg+bZbensaZX65fxoHyp6mY6cRWGJbOLHtD
aRpg9w6+tBE3xNJYvXkJi9ig8E24njR5mmbIWx0D4ORjztnMJaT1jiuKXlqUpe3lCWKi/8oRdj2u
c6VG1XbcQqkbwzhjki9NQMXHrnqFpDbwvi0AaomEIKDXl1DawFkDbxrwIV/KMtecENY/qheK9Xvu
rDnPhB0hSS/kHEErkn+yCeWRa4vFzS6mb7GkNltCWOrchZcf689x4sF+x9DjrXBddGURirPdyonw
ikTSjcNI+7yCbnOInhPEfA1POFjFHtY6AWdXyJk5l7UCMpIJhQjshzZOi0/BcVPT26EpGJ6ZIIre
aftWbko8uykawpBiQTXzzjoGGYMTna0cWg5mS5guEtweJolIgPg5K/O/FRuNjCjJvF0yySGyr37U
LJxlXd/w/GXR65k4R/EmetLSkafIJ8GS1fRYgQRlpEw6ZwFo5C4bvqMiX73PX9IL9EMIbWKdopq3
6PFAQaj2gjlXUtVK87Q1PbjGQ2MPfev1xnLwUS3hypdOEnxuITJe8MWpZZDqCnY8kpvvW8l2ONeF
MJpBylFDnooNUETXpWyCoHsUJkroqzX34n59xbFBcd9OpYCAe5t5XBd0pXGKzfmrMkJJGyRfo7wJ
MxExz0fZirzkWuctRstmCwzYm441sNHKrICfh/hJXO1ElqiwKWUZSheRU6Df34Czf9fLPszNcuR0
neyaAQPpfpCgUM3kffUCCU0kZvoeuEo+6bv2SybUtEhlZhUsQ/BelIubY5kWs+TMievC+GoiFR7+
6fYIYsID8zkpqbfFgjD1dIe8ZfvxqCNQ6332/cADUiksjNYZ9OKAcxEK0XXo6mkWROELNZqoNDa5
AAVfO+zBoQsn4mHgtl85AzYIc/05ZKlYcp71rvmMhjt07qJdtkI8PQd1ajOrlQj9WlFXmxOnXgTS
1GYRggRG8CK8OeMBQPQmCi+NGXCWbI0q9r7OlJq+1ZSwgQRs7UAa8C5hlaatFwi8Ub6TWuzIzCnr
4fvBx/Uj6Nj64dbMnt00MHpLdkKjJ6ZPusbtOuFKHRPTF1c2liSeVPh/nRKN0vYTHg2itVTbL1LC
g49WQrch32QFNksRBE8n1jCFbch6nGbilaz3Wsa/xe9jn80Bgi6l7xZImrIChmiQ2yZvtehZi310
VTNf/3WGOSfxkw3oTh7djtzJs7f5+Ll11+SqOM9HgndccjKNAYaJLjSZbLx766K0RvxceVVG6lG3
nXaovu/EmPVcWj2X0ZxSp+Wy8pO8OJeOh+Y0qR7DWoKaOrrquzp9A7lBSkOHi4m2fr/HtYcc7EIE
9QImE9CCwekU9ZxFM3tiiYp6e1PtT4Y88nxVhtcpT9BgzLQVpMVp7WX4Ac1o/Y43MpP0z3klycI9
aSJ3ZOZBCCpsfRAQO+EJncd2fjx+dcaLo795oUs3hPTGPw+P5r9/tyRb07gfcUS0nhZFJZvhwyaK
qempoLxrI7aCfsNzHz3dXpwlPduLTkEdTCUFbwFKh53GqNax0JyMESMbVx7x02iVmGpl4nBCRVGR
PRdDACLRbtI7tWRqPWuJxtVSMR5/TQxCcD0Di1wP2VI4YBFiqjL7vdVWHWckhbgw02ii9LvWk7yP
d5vRn7TqFdW+yn68VvBbXnZnOIVfGd7wKKypKxMKsOVZ0f4JCsB2fKoy2FwU1ZfFgtKKRP2fXwfb
i9/cMctz7Hf1uAhPV1Q2iGNlxmDOa5EnU4voLGj+P42qGxbVb82lVmWHAxYVCi4fkv7QkuD2eYXW
jupK7HCvb1ZlDyQi0926B9odoKNtVVN3UR0LCO73z/Y73YNYZDkK1D1wBljgzDuQuvoinNbIuhix
laktPCT8RKO/LSBK8p5IlSkvqLNUbjgq5UPUsePsWhiA2r22EWy50Fp+9exCCvbWBM/y01A/TcDR
0xej5lWBZXF6xYef+dhcJ7IZbp0Y64xsA3qvkeIDqytmaUCkq9Lnx5n15WFmy9Am5A5K4cq9N4Xt
ymfjXXLfwAbmYQuxZRm1H498CkmyxFo3NN3eF7ITHr0yutftUp0ilYSKV6tEbliG923cjN9sSlR+
D9mhFVHewkGNtspfIhlzNnCs076HHFYyZGjvLWjZWaU4y4sOAHQLo3KDiS21bDIpdxhYt4Jgbgun
9h9o/DS9B7eU6owrNIpHBO+qm9BbMsQCp0FxUHcOhmpu0SvwTgDxUaOrKDEOug9gSmK5IGy2vYAG
C8sHO85elp5RnBr2n7W0+nCYcxm8rrG5bDdiibODxiJbi2iwRhrfYckZisHxSx6dEEKktwyd0wFE
tFmriPvlxVKaklFubyvgbLkPDT5elJsvfWhaChiumYKjut4eg7mOqmntEy6M2wbfXg8XV3JkuS3f
5I+prbCDU6Rvder/FmvK8mEW6nqwJOIzyITFomzEtxwUvrfKpbQ4y7UVc5UU70HqxUO4mPkGQDdz
zmVMaMOK7q3YDTgg1k7xAPUtlZpEXz2U5TVVjrtWhGusGMmoPa+ZZpzIm6p5+Oh/QHtMo7fV8m50
lytBYPU2CPrXjtmnz4nK34CnRjiTs8x0/61L9LWnvQoNeAj2SPmI6q/qL2S04p8EOy+jyeT56s20
SVbY8rRnqqnrsmFP6YJHmpNNRvvKzzps1VmP7I7XNBm8jEmk7l7dlvLWIJorVD0h1HR+COzaqGFS
K38KlnEm9AI14aKNH3YKkZBpfYfzOb4qhj0QwjpWY+WUNl5g+MwLh9q+rZritpa613Ib0Z/Qlz/T
yG4Q2SlPlzEpLNLaZ7p8Pa+Dci2TGu+/Oa1xmb8dCnVrzyqhWNdGsL8Prr767q2lN4CVZvJGYvYB
Gp3Tut2btv8/7L0jpT8AoYomQ5ZwT5ADBhaYd6J4wBkAlAKGNpzDUMRzhC15e9iED0gDT6ZPtJsY
7klnfyu5suCZBYxoC75BfoMOGHMWy/SJQbgqWZ15lREFEjamS3Momncje2mGDk1qHz+ekWKnTfHB
UKyRoyPKwM5c1bXBQmWvVSSAS42yddDIGp6IUtrlagikITTUbsEnsPVejGMM9copTcKXOWGQRG8S
+4Zqz16uwThBwkOvbgBrBdc/Zs/jMou8H74Ky5vC58H+Dnhj51iTtUS0lMCpOF677xigbkNnTIgd
BIPHVnCbL+pgo3fAlZu1JkTRwaCM8aat8H+FzU8L4QyWrbRH/7xZAwyZOLsk9QIi6rR8SGbl0oyE
ERvqdzKN+lH7d10RT1h5mNI4OyH+yOhSNvjLbCrt51nYY4+K6puPJf7jqV4QfihYSovP1uqfN56G
NlZqVo2PjDCXv1Tn95p293pvWlngQCc8YJxhNsj2MKz404SJJCsvEfo5RYcOPBxUVEqMj3Fu+mUQ
lQmurePbbdAZLZYgJ9EAA5iLq78yNu1m6Q2ZtCgNPxKjALJCEO1GDUhtlGipORMsZx+eRwQ0mkY4
2o0w6FHZnLPmDNSDWSJ956cQE0Vqm6vlh1w2V6lDD6yMgHVJhO093xXASchUuAMRjN7JA2p8r4+v
jnnNXl4uz12ZojqeTS3J+SyK9SUXUaIyEYoo7bveU1UhqqZ7NeTTWgsoBPTlMWVUEjUaiVPIvwL+
i6tvblDu+ynnK6yW5BIppcKx34pI50h78Bq+YSCgdpsoHJTWksefkYqmF8IwqEFSSAJISzlUXT/Q
jtR/u23evNR2BZrTl4tiLVHnyRbNCkjl+ChOma0YNGgbAD3DfHlW5Gbx2VnoK7XnKxCelpDQWACK
PmLdMkZSA+fOO1gg0ZARDfwyInhjVWiftov2Z80VpjCyE32MpfY3yv9HY4UfKr2U263/XXBM16iy
huTyhf5RVb1TB28v77VKAIIhVCWzFZ3xmr8dGal0dmpK65g/t2vwaTFea4Np1BrYqkTkJFfuTxVG
/WPxWHe0UgJToAenYHwqvc0b5QdisnyAa1F/6LDzJNJ37HgxVkDP611TVF6cTo1dCI/Ya22iTAzU
bQzlV3bTRYkkOxcreNVFcVgqZJFbCsk0YiiovCFQ0Yss3cNqPlg2FfjxJIS5WNOviSJszAL0V/gK
GreQkRYaNpUxFnF7xrqhGMaC3edQODYUalP8LzH3QXFlWPmb+OYI5Hht0TsoAR6JT1XPL6kI1tQn
SO0pCHDha3GZ2lxxULL1NuHNy2938oM4kycUBYb+Odbwj4euH7Fe9rZdrXUwbMMnOHIH3XD77WWw
3nkBnTqhgPCEO2F2J+w7If2tD7ZfFVVNDh2j0r59F6brc8aPZywjGIhRe/+y8gUF819FOphWSswn
DzMpJ92zr7l5uHQXu4QwKECsTsWPui8wjbYWbf5UcZraGMDZGf3+2HQ28jeo5sKz3aY+U5VG48nB
8WehUrRFcpwWYIqPlhlRef5UHf8PILfObmBtL/w04C1/UuAbr3YC9KFZWpGh7LArYoP3s2DUqLjl
3Nr1YYDb7Pbs7bVPFIDZ2NVgFhKi4rzN3ATXQOWnrdSbKL01j182/zc99QDNmmSvjQcDBhtAp+og
b/Z2Kupt4CFgkOnJToarSn2Eua+LeSve5+lgTeG9Y0qM58c964z2czYTkWZlxdeeQk/wFBOUcL+V
lB5HkI/rWXTS0g+cKQ8ckPfvwHn3SpHxP+08JpU1E5u4RZA8fLP371iqnYcX52v05uJiFBLOkRjM
uvQUY6uw2lo227tyVXUxuuxe1OqUDo6feJrOlVSox1h9NiqAlyKwEhx8GqhEbJFRvXCyzqnucgVp
hXeeupfvQlmh6RyRTkSTuWzwJGw9hS4WeaRWODNr/axYhLPgQDzx82aQ5Zg7QhidRS9bXonN4R+W
gTeokLojP7vuaQk2aIFZaAy9hpnt/H0y15xlXLvf8Eqxpb26iheCZAjPARWM8S+jfHFhm+XlFFju
Vnt2lX4EY66qOv3gVojaBOhngDar5D/GPoQjVW+lu4UIjxO1ET4XI14EEGA8QKNtyKprCLzJPap6
6ZQdOOxabNqqi/sC7GDJog7hZN+dM7JxYJuwDvsr5ciy6NYNw8uFLrldU64JSPqDc49pMG7759R/
JrytMhOz/9PABfoD3H1u0zHFT/HUlUp9SWyhm3lOYbj2ZC52O8Z/6jzz7QiqmyQ0RHzm+9n8fgPL
yGA9JD+CZhQeZxYuwPwuhQxnStF95DTkzPp+h2aTJP7u67YJu82ICUTzFh63oFJCoCgcfg5tC2tN
SIlWknxwVXOMYJghxxNQkKosYWMGNLWPaVxrkbp55/H3nuBCFq37ASQNqKkbH+w+6QHwkDffDAM2
vWyMBzH1JjT8oEP8BJEOysdfSu2hterXbhWmu6fyfhCVUwxUvI4zGvsHh1G/9ELgmDn951Fg0uV+
vhG7/E88rKAgHhQqLxinMk9fcw5DznmCgTO45boDB8/MYHkaEYzwOoO91otTtlVm0fGJG206gEju
o9cTkT7YfnzMEGcSCyoLKVTJIu+9SoWIzRuYaYyvQ4KMo4DdVqTm7AHP1Te14zHRSVF2oJ1WuT5u
6AyNjuFH12WW4yCJeIbxBf9kGEJh7aBItyOr2El4v6Vd6EOlACzYvtleF2NVYvKofJJO5Fb9HS2c
jhO1AQPCuRCHfOKCJ9OX2eMzDtzgcNCdfPNmjaU2EChEujIPuzq0fJj56D5tBjMNxAzckduORikJ
Z+/2EBrGKYe6IbJY1qwGmMBOyc0K95yPsJ1KbFQuBIT2wiCTV96hfFjrCGhaQqygG64GVH9QWZ9L
7UmAKu6l3u/iQumIAI5ABoxxtC3dltCjG0EmQ7f/s5MX2D//a4HX4qMoNyL1a7ucDTHLWozd6FE/
3mk5080MpTHBujGvcjcZvDJPJTVRxrGC26NVHS1d/JBfuqomXQmeBdIUbPxeKRo9gWp/ULNmHjE5
saJ2PURsLbB1bekRvARCnduC2A9svKW/D2r/dxMEV6LIWnmdD41z4jlQl9fxJAX9M6gfb5GYOgbG
xBHnC2ifCisX4iMBNxUZHWao6xGl+wLLKtsHuDl4zFPgaR+UXdjPenRoQenjAUBySp4cMY/pcdka
U9xHnI7H7kBa5u9Rujnh7RBfE+FKbr+4xaGkAwfOhPyTOahFUBiGOO31bbdzvhDU/5as6YwdAuwU
w9ETXbtwofQ281iWdjKUxwOj0xQiIxMvXgWDceyB9Oi3eqeNGI/PlTL78emRteigd8SkY82L0lQQ
y1zWpyThV0rkKkPC58J3lTvKA7+wFhiNxcjFfc59UfQfWcYrYqyhTBUJdQBoj+Ld7C5yrW/xzro1
gpFUvrx9nbX1b8U4u/C/u+HRa1clb9S0BrJ36mZLoyNlQO3DFk/VxQAxHO1A67vo6+mE7wiWimhG
KTLzK81Wb0d6S8FIB/E/wRV71AFf6coI0Aqo0Y7hfSXEiC/Z5NX7x+Mai1LjCupUmUvoJ/rmR+eW
JcCwYEY8QbwFhf4G+F2wHgWlwXi0LVk6FC7fyKPe70k7tQo9xc9fW0+o1ChRwtpUq1+6+Lxb6llS
9WlZAWh4GN3tOFM/YPtk+NHWEiWLGoD1HFJKDTUvY1TAnZJEeTQiPO7PtuPIxFjYRQGXDyllh30y
1JY8gJbCaBO/vsUpQAVTbuGvUIWR/7vULe6/T5mAncF3XHJTiissBDxD6ccm9A3Y3ekOALoCXGMC
W0SM1BAT/YoyOGPv7mDKK18N5RWgvhkrgx589livLjBRxXpqNsAvWzN80pZ9l+0QpM44gcaT34uU
v3gLWqjHG7Ta/yRfEoQP/Ioj4Ac8ajqPb+D/sJEPfMW8Bk0YwdLPMs6OoHCP2JXOWL9ot51HfR0L
D+le1JDuqjfHkJbfjJC3jf2VTLkrLnowkUFFLsuQ73HGyiXe/zRw0aSd0bNcaSw9Xk6wJmx9FLuP
h63RoU4otUvFRBf3llogVCXwp5NOywmQbIQnVDoMnnJeCleWGwvRX/SL4CtL9YuT9hx6vCDtlmme
h3xwDtF6KFyPT7uNgBg6OUj+VtzjzE5Yi2XSPEKA0KZtsj4KJq5e4dlLWWL95u5kmCh75R57SdGQ
eQDLm0kxD+z0Jrb4opz9aotrNGYzV7wjHpAomo8POrXo7Lqo2BzMYa/Gm3d8ytgoaqUrRJp+BfrV
zuZJlrPILy6lVHj24XgV8E82rCIU4b38jtP2A/Pa1s5l5PDitayqWsxKpeuTs5/fxXWoQ++w8+t6
XCSv0HTYpzQ4KGKhjbfKJA49TmRKMGm1Y7UdQCdXCXKnJtY4YlN+lRWQSs+pmAxzSf640jG1bTpZ
0IdnFrDooCZEh0/2sgosl+NkZC5l9cIG6LCo0jb7kybAWebbremmQKEKeNTAyWL5kjcbhJ6HkpqM
WUxIw6A0ggVEzLXv7xsSMtEFGb9cEYeeBCSWblc+GVlJXS8FVswOFYAlWLMRvZS6JYE+N/5cdYyU
GJvr2GMWRPhkIAB2tEH00aLrPkBKkq09oy2d4UxsiZbh9cNgrwQrXUBDxOPNQPXEreMrWLLCGTZx
KT2Bgh6RNZFDw+N247QLug5VQHpdT9IeIUGKZn+bsdRddRpqfLD6w26hS20a/UE3qXXo2RIYQvOv
9ae8gzdlZ+d7HDpR6oY79nbXwnXr8zAORnK0B9E/hbD8QO533tfD9iVeWa5PBPnXacQcKsN+Lev4
nPOkPomkL6BbFrq7e0AF4qglmUctGRPsN8fGfIYbZbR6UM2uyycA6JpNIfdXbv30dbwA7/slt0Us
YAZHbC2M1K/nbBM4PTkFcNVHfxBqJtAzBSPGqTn0utSXxbi1cKglg46k59ijW/pWQgGp8VLZJX2D
wCUg//Irg6N9ZA23bPt3YFKJwoH/wWA9QZg3PkFAF1dRC3GmSsWZ71JMfB2+ZPhD473HpWfs/oNf
qqbJTzJ8jCFLWUgLrWvssh3aTI/UL31GpY3AMLIJyWEG4hgEbGu022WJGvdPaLYtC4+gAwf/uwE9
2lbyX/RuUm3rGmcoyJ0i+KhU2s7hr8YSHjRhHBSVViDWFoFw5bEeH451meA+HHdN2IrmxHG/Ckev
1XZdz8lG6nwXDTRon28ufGKxlX6JH4eYnpTAaCAMhkL/u+57PpQsrDJRv/jb0s8udwVsYsmfmCFn
ZKSVColOcyX8nUwb3zULxTG0kM3jkK2QocGtHY4rW5xbFgMBZZmwLMaSR8ZS3egfLl0zIaIcBZjQ
6r3WrHeqIfnCUdsg2ZTyl7qpj5+dB0uihtcJg+6TSkjcM79QUgSv+nAjHOhL53jx08WJrVuJAr99
Jg/7cS2QtXSgosszMMc8rM54PttO2PVJqUL7V9qY0yB+E8FuO7J9a1bwzTMF4cHHAYLwDgL1g22V
5+f5U9Ycy6x53UFP5fH7CzYd50izipM+9U8OKSWBZGLEZrAOgE5VtKgk+K4KMXQHvLJnAFumShcN
CuRAE9kCg3+r26W3Vz5D1u8k/t9sbb9V4fmsi9hoDeLNxXg6Ush5fHHECJEcC/So33zaMNB0brx7
+/7+3ej/al6JzNi4WNRDTJHq1N+Swhl6m+SMclxy9R+tTXDe7V43stqadLeJdgonLAjlMAxhUheN
5yZ/mWdGpfNLKUe/HnUqIz6NzSkqkdfcqyQ8cF6GM+yUTzK1YLeRH9YWM3gV7Qznb7MnR3esPXJv
9IqithCepVKSL4If82vbkrQn4Etk3AmUqa0BxrCelYekmkl2ouBfKz2DKsBSaHLI1w5ka2nHfB0l
xQ7TWdU7/7gQMtZA0P+T6JnMk6+P50dce0MsqvHlXFD7PMG0oMR+iTmZL3jzSNCOzPAAfyy9LVBj
FpzoyKkm7Gwgdt174HbuZlABOGmzJIpatG0o1d+90ssApPvy9NRWIKctjilTDtz1u13L/Xecz5cH
/SpO35WYsVlITUXPy6V4RwfBjdGkVoy/DOKsAGN/HNKmC2pJg7vQHra2DvHNmaTM1qfNObg2xFJs
mBtfWsx/M9LwG4Nthiv3xk9b/GKF0gvZyqNhfjniMejYbOa5k/0ILtvO2igSguJQtV+5abVmO1Sa
sWX1AIfALVi9JqTCVz+tIxrbNRvKMYNQRXnllL1Eoa6hW8TvE23aJQspUOOfX8fEuunfyHWnHd/L
REDOT98o9jkjlMSUku8SAXk3SHIJjnb0wgA9zs1NAoNOznvv3ddnTCM5rUYVNB3sD4xXJxx/83gU
LfiJgw/JxSiLGjFqBZviWZ1MHFrUX1q9MFFYvYqPVQ3irHt5WMXV5Wl5kQq1CaWciBDo+VrgiOwV
Ljmg/yjx6xGWd1n1li48swLmfZemqdnHhHSGdcw7euoSI+k6oX1kNsnzmcemFoU4nuV+cIOo4TYa
eHgi36TVnWhjkr7hCmeuuvEolRKJQM0pKzLy369u10aLrVZ4DE2RdPZGKC6yGzCXInLT/A1uTDir
ex50f91qf9Aa1nJgDeUkDW/8O6MgpSny+H6HGbKlXmz+alQxLhKZe4cipVDPJXDkfRRIx8HdAVt2
YKGh4vVDHvNwLoujHX3X2aG0nySbKzYtFCv48FPOt2y5rYfzx6Y36OZlsZZx+ohUyiREkad+Xmlo
yETdegqoo0YR6Otrf134DEW5UqaIApOwCozR0JoM24+KNhCSaPCWmriZkgEw6HJezof13oZ0ibMe
f0QfRKwEaSXKBdvd4o8xC5Yv/EarVDPUCZCgMiSh+3ci4K5kZQ9PqoZcYFoCJEG8B+NG+LNT7HJF
BI3T0OIlDtLmdUnX4hMtzLTel+A6RZhGSWNUT7uz/3ocknxzSXaK4Z7N1w0rBulDTxluSMrHZHfe
ADfaQSjtB8loQaY+sUZMwLOMuBT82LMjrTu9fIriobDzNULuTpQsHb7wZw5LjKuxLAuPeg5Qn2ji
5V7g6IbaTqMSipl9otQCSv/G+mjtMU5oyziunxsFoGxqBLsnJIwrVffEzs8hom4wRpR0s4CPkXhI
13w526MMtvIcxRNqkOXnPztvr6Ez9Kro6LI5hFkWtmIm8gty/quEU/UR2a26L99Ln6HfxN7u26z/
la29pq4D8IbWyJVwmUyt+yguAmHX6kP0jHznMueK42lzm4geYe99kexuMtc86HAKlV0hBwPbh2Tn
NKAbXTXs/5mANVgxkxZnuIZzC4FCkVw8y6WCeWgyDKzAag91BnqbPE++igG2HmxPsxi0Oq9fRIfY
zwzAkm09vxxZfEu7J+t2QXcCp/qun6f5EnqbhG0ka00q6IyiRmQ2jmzNPwdtzfx69TPrDb5z/tPR
i71MhgaHAJUN+KOaTu2gQmuQoUWo/JMMSCG6Yo1Po1LfrgtlEaPG6cstMCF2iH458KNztS854fWB
oEDm12QG9YPl7GjAfQmOKbivO3YW997isFumNtKynXaqMLWoGBjT3hZLwCuvfjCaua4Ekj6T4H4K
kyEl5cKpLpl57sIOFPfolmaHUpcLXTYLlEBa0v1wwVrvl0fyzrZM7Ia1ankAfCw2yKI9gIUj65+e
I/Gk8pSZ5a37RkBO0LcZnubW+Bj5chczVQpHNT6EgTeqcbKOWi/kQtrE3oXmlol6B5hr14g1RCmI
Udoz3QnkhHGJMbKY0XXIOhhx8QyPqKiOViMen8Q2RgJBL0ljt09wR5YZ7PFX9On0nNi/lyQDa9aJ
Y4zU8XvWuNpLbGGBNB9iyac95rfg6PbWDjtcdwz0Uii/oMS0p/GBCtS0OadK3audZU9WFMmoRnz2
8HB6aNTXSST9U5UNHv5n1sKQ9Kjr/QqRlsiF++/2vrAqu/9XP4E7IQ8rlO0NTeWazaWbA60oim1i
kusIxBsEdhL6GE13f5poRjQRD4LaN+pyXfbA4U0z5Cj3JMLLEe+7I/i/OqefyKxzBmAAgfrs50vE
lQifLrpzYmr/QCLwxq488afqkxWhGWKRtNBh9RM4iFge+3ekHM0RqisLFQKA6qgth6b9Qzh9L+/F
T+6WQWRAMIsV9/0eZvYZIMEO1T8whAbGdskPp3lz57BoQuk01OWJMdYc31NtGtltHvsfOYNSOW33
v96Q/fgP4kh4bMi3nxfxpwBggHuzNDK1GT9LYRhMuJq1UrHtKmp1ugVJquL6YbD0NstQ6+7lrwA5
wSUcpfQpkNRQwUeTwut4RMgNVvQSrE0oGUH5S0rXkb8fWhCRE0UegFRo+GAQJv9ufc3Lz91Sss9t
eMYKebssjeyqtq2yUJ7cdLJxiTGJIkOXbt0b/IfhITI9UruspFl82KdIen7C1oHeqKyYiYp/pcAu
yL6TjD2u/Gn8WfQv8k2DS8PrRdW9eczz34F9OIFm11wpqI3mNtLUltR9MzMnQaOEQ3a9rR+L/yaB
Ji4I/WzRLzpVCcYJ0YQejl5oB4ebWgPvTTaYlEg+ItPPxnaBQPKemNaAXZYbzndtDVakvZt3vGDa
dULIZ5S5/b1vLW4cyR+JTNZmhs3BD3pAtBO21En4uwhkANPmuOxDq5pX6q9bV7iEEbjSsCQWfJTm
i4m9OzAW8xfFX6QRCoyJ+ampGtbtbm+3VZna0vOq+jhI8zSoRyjnU8biDqdqDynklXbKKpDcSDQ6
UUCkGrLrW5m7lw4+tNWvWATeEaytk7VwjUZybnekyWacu6y5dcqLIg2Hy8Aqzj04Lh9aGL9gRdiK
wF+O214Sgv2EydeA+rM05eb/4fIAWj3Zp7xA4xXR/2liIbfwN2wIJR5GUpeReZIEtOfbqpdsNLp4
UnDhvoeTEx54XmjMkZ2q4/fX69IFiXtjIqQ3dB0qUSVPLXdIs3Fgcy3UjOk1u8dUNy1YZ2gzGdCv
6VemKUUQlL6hfcmPWa01GmvnnfBrn+cOQ0N0c5kvkIocXRGV+mbHKoDvWAboWGeBlLsY9jFLxiGm
PCcWWt8e8D97BGJMzVk5PPWUrO2Kge1qfGTTf93658JIh6eMqbdzEOK9an/wTG4xXLh5lbDvYz/s
mUAq2+tL0YUSau3P9HfrMxTFQ9638wX2JSjTmhIJcv4f7IRIBZa/87TWH72T6mrkcNayyIRPFVul
2vgxiAH7fij5HxYwZL199c6ukGBaRtDPrT6rVSeze1udkZ99DXEa2vPCvcwpo3JDpCplkZMnFrV8
wUiQPaWMG81/KNjhyP2Mw1QVu1fZGQtKxkG9d0Ja2zc/djaTTOMnSK74LXqmVSgtTH4sN5eqebYE
mKe7OvvcVR4Gtu2TFvNmDbrlY6YWih+5QT4I5bfXFuqTtzDvPqfOT3dAwQbuPV+JUvMicoSNxI2U
o6KR2OG+eKSPzmrQ8PAFXmuqel/sX8h8ljmiSN6Khl8/grRr247ngnrrSpcuJ/bPDtBmRXpXkLFJ
uujo5hPgKp+H/bRgJeU1v8kcvoOxGQ8DYtStC/7CAeou1f41bRA+12EomljTweoOw95zQ1zvR1bw
6kCH9KynRXxlstuiYkGBsnZqaUqevfAd26X1pIhIiD3kwL3nmH5yR2Mne04ztQcwdHqI/LH3C7wN
QpNj1fm2litsXFoGvDupXn+goMe3wKlmtw2EF/3UciDk/5LmYjM3Ep1GgGVxSHn6rinTOF6yuAEE
uelZPmzGnUA0SHfYUOw5SbupDvKXZHPYBgDkAnwoACHFq8Eee7kurv8HlbqvKQNQ/uMaARTv2frm
OW9N03oYYZu5DOv3ymqQJPVHTOtRfIKDdTQWZHgk93XThgYo+FCIg4ZLLwIWM3j2M+tXYN0L1Iio
akIg3cwnSMAPNUktN+KbLjlSpUeLPC+4SKYEMpCJClNKhQLSMiEtRLrmvQYS+qf4tpmS6mIE3pUg
A6xkMRMpWrBM3mY4N0vJsjFQuUIuC95g7vW3kRFuSxcr+Rqa+Gi8B90lGlqJVXiVbnq7AXh7ZHPA
+caxiC38en6BuQunAd5BlMHBlnHa7SdK4eCffNvhPlEZh2c7h9gTqi27sxCc9kG76ufNO9PHas7G
H4c27n4VYkATdCosGiGC4V59EyoNgj8iC8Nqp3QTqukllcRqTXsx+nFfOmY7OjqSVTYKAk/zL3Yy
jexFDP8vtRHziRFcx3sW8yrzIbLzEw7yrkJ356qwae68TdHR0W7NHdjEz6WskNHWFysDNVP689/s
XWL18ECd6NXDllDvnYsa052VjNMcoDRKghwY8uRdLbNSy/BPRDYc+cwGJx3AMmPw5FiRZD1R4Zlw
zV/+X38yi1BCmqKLv6kKfPUOVA+5FLWs4VTcjtiJWIsTJSzxqpnqVmVxM7LfOlUKANq83RyApcc1
LIE8oLIrGRm2U/nEXZM7mhu/dlW8DLGzT3vDXBTwkkGi6Nw6z+ak5DHsl45IoMnsNf5gDkqSAjQU
G50tQJRpG9PVTENQfVDntUbAQ0X3pF4lkYL4RJjouViKYm7nNu5L6XyjTnfXCbh/Vn0HcKGwJdv4
4DrquxuMa2NhSNyKmMjDfeDRN74kqe+H2yhULYNcyKO+nzxRFxEk9XOijq6lN2F4AWmzxWWHZfco
aga8AINre/ahDKVrfRqMFpe/jtwG9pdAQJDUvLgNxcgU8K1WiD6/quYyMhPlohHiNi1oU3pLDos2
1ZI1xlrPLxc6Csvy2pVERt/m8ee3DJt/LsEKR728Di0ux8gzEBiPa5cHxwtrJPTxDYil3ikZYmZG
wlwNOmAb8yCouqnmE0NMo9kG58XCzVD6LAY6GxCd1C7j0THq+9GeAIKUke3mWdT7syxBIIzVigTQ
SEWjng7ItzGUANycV75bn/+c2SNGn+MEOV92LtNNdATdDMNa6JB6OpgdBAXI6HVo6zZUNJ78iC1e
+fxQgIvolq7FU7injt7ED5belxIXRooBdPpMU8I5zmD6P9k1tFpAA9ieiml/RVSvYEY1ZSOtEKXW
rgBUCgo0zXYEJhh4F/nusbTGXZRRswAKNN02PisS6VTJl1Idi20ziBiU6ppPoHYshjZiRfqyrwef
urm9uK+0VK8nkko5bsmmgfCakHAlH1kQXe19TuYRWQEe8Fh/cImyGrukf6aImJwQwsN/sTW0nopt
lw+yzrFDU+b5trxXfWEqSAoAHZOONiS8T8IB4PZWFfG3uInWElDbszgnYKGNAiNwiZme8Hu4jf5p
vp+qJvPxrtIRsjTisMehNI5iGbuGc4SQ7ZTBizPMnW0e+0d3I3jiXEMK1jmqaHOl1Hef8ZtFGUNj
8wW+xFD/DJaBCqkGozjiipvMIapZX+GyAaIpDme0cxDIO5f42/0GFx2y0ixqFdRczZGIPmNWJTco
2g2dZdfc904pxXO0sTjWCV9u/FTJ9AaI13I8PPYZP+2S1u97+h6IwGgUfMHxltYwY3QYuHCPYaZo
Hy1u2zOUYDLwxz9nuhKH3rQK/VfNbqZ30xVR+SdvEXd/N8+z6wv8UK+3n7hCsDTJAoaAjSritp5H
Yi9BU6kf2GjCexaK2vA39MA6OMD8hj4D0PgV+tpFHlNS+EpTMXPb79JZB8rJV88Rkn5xacprdnJN
0gAjD0Ua9PzUloxN2nL2e7Fv36wq4Pc22jzqlVn4/P6AQv1/I9G624n6IWL7burHe65zOOcbszm3
nN7b92VEwE+MA7DmqP9Jn2+2xFxzB43ZP1CLECfGiHnTF/dEgINTaGpo4AlzFtTBvTYml2di0P+P
zyUo74P2sqFK5YrSXQE6VMGCvfvox5teGn/uzmLzaMBZxn+kdQ00CPf93OkoOhm1Q31gOe1oQKW6
Fn5UB/EEOeim3T8KtLDZvG3Kp38qhMmnkKKhisXesWn4pru2cjtBepghqDlbWV0fG4CUtJlUmJ8y
Kg7kCLqyl6OGIoZQbZy7cFLEqjY5FKn73Dbqy9cNY0NWz0NnNpgRtv7dlBzBHFYHsFGur1lpvHJ3
7IMW8uA9vZ+AOha3G9CYMMIbF/qCiJtCPBA50iWE4rXnjxFMOFM1EPIZA/66nT8MtLS7566oB6o7
2nE5slzGFVnhjGjNmRXOpX88xKTLRQ2U3Uyx/POZYIpZBkSOSGAmpim8uWmbdTg99QX5HhwdPfI7
Ou97dfLIbruAgAOcjat1mOWLVsKy6rhjSYgRtu8FObVFOhLnKd+/BUAj3TkDChvz2Bt6otVABiX0
ZlqGHkc6PGIuCCEHuP4+YvvaHwQ4UuYcRIzLmMhKuZYeOJMSIfVRg3t4B8NKEzMwDjirK/qqALYF
sfCzpxnPgLrWP54mbGKG0T3FyLEjD/hRWau2UgPomIz83NjYToliAeGJ6vbAlC8BKSqJH8retzQj
10C86QNZgWqWhjPeOX/ooVGSI+V3/9S5o377NbcOkFYetlp+cs9SeNMkuMQU5ByPPnCCaVMZZAQJ
PT9iORvxwPaWqL8wEEAfBK6bT23oabLJFvo0lJ+MY7Zd+H6tK3YAclj8c7V1P4y58H4k86BH2rg+
cS8YyLbFNomqyONIgD/36W2zQa+WVl1ndR9zy/8tkDg1QBSRuwRWsi+5YC13JlddcgHSYIBaRQKq
zU+sjf4fyQOCCnM5H2AAOLEk4DeroNUSQuZjIaSw+RNn19DuXY5Vz4lcllgHqdD/glUvhEmFEHdq
WsejOeWG6m+lY50OXaiY/dY10zcytNugN6G/xMP2hGeTx8I7UkpR2F6XNPvtgawOSnfJIEnxeuXE
ZB/Fa5Dkq2cM7/mOHK1LXk65dy74FySZI0fd/j46KPv/Bl/yN9MkuCafzxYTA+/wvXee8SbkHfKh
bNId5uOS5w4Pw6aB8phMt3s9/BJOWzsTon0xtQRWEcKStL8GtC0WCJB62l4COmPZW9Z91ikMgPDu
YTcGQXp7q/VD3HS5sT2RYg9kGyE3oQRC6DhZ3zBx1IcJYNvgrJkk9pzzqZFM0vQGKkkmmZWV81+G
mgkRg7Hf5zXVC7X0W6jhBJx5Nyl/wn2gNWMhkaA+Slhs+EatZqOR7y1sWGc8aNWlffLHPRubAAS9
0r4nCBPwbSuTip6UhrjcwpJoSaFt4hYaZam1dWsB3fxrSokf+2ZPD6kLQ8OsG+rknRb4bOULb3Rz
HRRidtyFcPg+XZx4uBnHLyTnF1AvuSgtqXeRlNuI935KHKANcsHY1fDd9qoKz0sqBnmJN5S1Y211
BOSm8Avoa4FrioHzneKYK4GhPh43armREHnDwmR+VTfG/qY4p0vvstpyEFxqfBsk6U6k5lzxHJe9
AFQDiXUGRWR3JYGA6tob6mX4ccLLEYxyILlbLuOUjva8thEStMZRpGgtYrf52n9BHqcnpgp0gWHx
VZcI8ou+qlbqqjcmDSk/JKwkt/yHT5kpUmrb9Z2SiQj0eEjhdJqBWvdC9qxbm4r4LxzCo84MI71d
Hsec17Vqurx3tbgHH8kHcOX3NGn8gnNunKr0nSXprbRQiMhYMQIDDluEiOGR1PiCDenFNCy67faD
QtZ7tvvQ4kWr8Z2epkB3Du6tMgAUubuPbxKOWDYYdpT7AuSaCWKahm50KaGzFvnBbFDFJk9360ie
m+wMvgB84QMammEDlqeG6u7jxfLcRzgFjfKwkXzvmQVolzBx6b7poxqP0NDXOZjR/kUTf0YFB9vr
XzeHAXH8BX7Lsea5jMrppfVFwtM6XBvRtACUkSgj3g70fOMEjLKaP7SX3lFKnHK5LC8PralmUg0x
THjxavMI8i6TuyZ687DoSKXWVzpzIORL+i5OHW4wvw/OcXtQFwD9peCfBvCNRUYvJctWmEjty1rg
2SYHQE+44yPyPzM1G5RHoNuYj6kDUva3Y3w+1Cf4puPmf/bAvQH5ybO8FLVqhFPJrxtjdp6bBBZ2
TcqvUQ2INGa3XLlnfcstd0nNt0kn1pcGACbACeVBqq/mhbSHrrFy5fF3U1wg1dXqLxUMI4F0X21/
9ODw/9GL3ngQqU7O4VqtR+vleceu7LFnNMTPaeBoaQdPfb//gVktQlKgqImwSYqi5wIlp8f0uNGB
CDuyXlHXgwxSaTtiX4eiireBNoNWcT8AD0RRbZfyx79EeSAFAmjNMJmDFPT9ILBtODXPhgp21aEh
8odisVn2vdXrSXg/aQEW2gfEPIJM4pm/+yD38S3XkB0UM/EvBC1fCbeMsUtqAo183GXcaPLHjtyH
NmkIHxScHKsVc/wUtpU55noc1YKEvM1Lp/OSqQ9quidR0g/kQzoJp55kQaDCldx5gjAesRjvze3j
bN5966674veKx5AVVF2eXM07EFQXZ5numzWpvS+Hwx19vyuG2Pht4ylMn0Xs/iqeHmMTND3pNzz7
eA/rf13Is4Wuk9H1WR9cP+/XX8CNapIxPsvpubI6FIblohieHluW2JU+A84EcgcP1Jo+EaQTv3eS
Y2AWxjlBRMUM/e40QlKpq8XH95yQWrkJkavqeBqfjKoVUrVY1I0iagTyDeJYn6XanWm7UOYjuwyL
7InsdZXwvvopQcBst7vrqSloy5lDPnjiFx7ViVH8Ehk4TZLPXVVEuNdXoB6LHTAhxr/cefy0wHfC
iAdOOfZmvAXvpl+cOnP+uyPcDxok3QG8VE7j9b27GjGeLHEqY0HS44N4enO9lmbVtgYh1Att2/D+
yLZfujV4mQNqFtA5Ak8W+1T4yZ87hDTwSWrYHcOUx3LUh2DdhfCPmMvwMya6Pbs/cV0ty+aGHXpn
KdiIGCX9i5dgkhw5GvE01wK7XOKUXUuCx2o9qXG0cPlZrMKK6z0iSynFh5Dcue++i2hS3emtMl8/
IzTfT4kCQHoqPP0kY8uTymiH+qNoIqV4nLz7DhRdE+XysCz0rigK3mjlCkzLPFE3VWCeJ48ksnzc
JEWa29J0L+lzAwC65egCzUPSMkGI7PHsP2YSI3M3SqvqyHnPGXOnI/U3UAtRjVQEJzvswhq2UN02
ID4m/BZbQDS0uiS2+vw1hufIibN8+8VjV0yPLlmXdCmO/55fAO0zM81XqDSnOqFctqn/BVctru2y
e5p18aZ1XiENmRKVnltDI/2Q4mSE1DV6yrdhpk+P6D/C9+Jm9KGkBoljhArMaE7FSpPCp4byzTbv
hnFx/jvxY43yCOJUH9qEVVk46wqUTJfsdzoPBgYqGz/bT6NGhnbz2Ie9nOB9mmtM2lDongJsxY72
gzqcyu2PMRDjwLfxmlnpphinpYl/f3A/+IgnJXGmnPd85nURxzsB+krjkk/F6XmXizwDWPySbnqd
3AQkojDELTHN6sD5+W2lqla1k467RChBP1PhcKqnNn9Y95DGaw4dLh/d+9arjsDiMswbbyIK8A4S
KY7Yc6Cz8PI26aPYazHmvQTPfQlTMlRVLEectXSBSrO/jvWzWpoDvdE1rIYhemmRNZ0zqPryaz5C
jh/RxOz4mmHghBhV/jVISVxkx+obvVzjVYxrkS4qWdlQapSlKHH7G/H7vJo3b7bcvMlmqaisIGlJ
lw5kjR4ESKHGtO4bZTi+bvNrN7iMJ4Ucp+WFK7Y2crEdzgXb1c3YWubUKeEDGiy1esWVWRKsmn/k
AS/YoKfh69yKY4JTgvn8LgeXrBp6Vbb5C4qUQ3nknenUTEozyThED1/tAnNttafu2GY4tVzm2S00
jObwAh3OBYo3Y0851qGcz5dXdGxjJljv/OG/Hlz+6fNzXopibeD3q54iuBHKhn7J0TvOCMteMR9p
zAJ5n43z5BfsI8vpPBVwRwmafT/5mI4y0lwbelCS5Y5y6ilJoUyDJb4NjGJ3OiHovbu03CrFp2WS
T+rPu3dd4UFTrASlKq9N9TQ3Wc/URnXOfbxJLFLSHQD8hIjUIJDJ4HQ/bNENoKJ92XbcuCIrlUr1
AAhq4DYcbh0+LEXjdcejeqdmiVXJtXew6v1wRBZBf6hQ/eVc+eMtCm6yOrAy8BL3Jynh/6tAihtz
0e25P/vbVMAjODtLgd0WrHiOBXQQJucaCS0h3Q/Udem30JF30pmVFa7uNq7x38yMmAcroNCOjvxp
Y/vDGXISM9iph2RSiB75buZAEoQ4U8WKwjf1tvfjBCfPlRmN2ebvstq2gZE4d5TsdFtKqUd72eak
UEOmQ7A+gsfT/cVDNy07rIUIfEVI/MYZltfSPHnmEQ9E/uZreGZKvcl15+fWIW0jmXJMxn5voC8X
OInv25letzG3vvtMl9j3Mow4w1l55DxEUTI+ap/TBoBpZO7sTHLUxUPRy8gGIptDyinW0hIBjZm1
ey7OybfNvdv/YFSLf2MyK8zvDJ7mUEsSy0t+5ewVUx7VdE1mCJKX4cIYPF3yzhZBmZvyvs9Pdp13
zkLZ5M3rTeRa4o2KUKkjIg/83skUafXNWw8+AuckW/oaK7ObBAU/Vct9YHZqaY6xFOXnECUUQPGW
jXCw5mjSgHSHsu7AKihtVKGHixa+AblPNBOMMMJGULeluez98Q192FBYaPXfZe9B2nDL64XioAsd
xjI8ziCAxXuVEKsM5scOYj5mGMXHvwQC8oHTWB/FVlMVK31OalO6GC0lCXsf/o9z+UwI/a2DfUSx
CBLkjAwhjEXBWVcUzw8bLoHqsOtbXfGLCV+tRg+75aFYeAtQB7SL43PdgRvOciWdjw4xr/FY6sEQ
Orq95A4pGwq2rmBqQ1g+IGVMsuRTxn0pLLiFY8KvWCLybHayK5+nT1vNt+srIAFsHf3hWZ0GYqCN
WbaIM5cRhQ5+pPIosdacdAMlRA0lCPEHUcy3VpphE6WWDJW4Npq6NmKZstwTzvr/Cy3D37kphI6X
cJdEoSYGyM7JZn2EcddWuDcdpEly4QYeIdPjpDeakgfbkCqjlZ9SAbsWi0259TjblexS8HBBKSAb
KovssYCVl7BSUnHuZ8hiFFWMvE4atTobh085FBm7emj2LgtQhUhEEcVCfbcNN+zQX9XfG5Wx8E4S
oWFesV+HYchAkqNX6y7avB/y5BLhCe54p78Do6UTpq7E/L4F30jnlmkCf0DPk0s41GljBXz5z7xh
PuZtEWqxybeflzgIKEFWCYj9HS62P560WSc0JBhAdS+dv+9dSVfCi84VE0EYZ0M+ZVlDIyLIjMN5
LgjmcjgU4qaaGoOWXQX2Tdp30Uogu4zOyIk0WKQqZD14CRG0v5HMSCL9YlhFgNjZ1D+dySnJy8TO
ZLngVW57AZBMO/U0aMcBMVuXs5aDjHvxH6H78b9qzR6wOJ7kDvof7KYN188LwWA6y30fyuu8YXnu
qnnIlF/rUu9jCKfHHgQIAhrFclZ8nVv4lvmWwgfDXnnZ4QP7XPv8Un0NvLgJy0jtw81xZ6P6PeSF
WyeJy2bRa7wPA9JcP/sOwI0wekEWHBdgdgW/9uAISE35hLLnPatRb35etwKmPfBEwElIkmDXm27i
kpBhyDDqJR1+ZvYbZa9R6AuzDtCWLgppEW+FngcjQg187SnZzWaGZk4flHFn66dDyhj0UzwC3VtF
xiSej2kB0sMKZ5MKOgh9VhmzeW9VaZop3bmKPehKpXB9xxScC3+NP9SyUCTBgOFmHz4cSMo4n6Ja
0P80+j/uJU4VhZMs+j5toXpNJnlKNf9ritI3UQ4b+iKjU8lslmt6UZTOdgJUSglIGG5vGq9AZKuE
CeaOj5rbJgmHuLcdcW5qg8rdjtZUIzVEWAl8LFThKzzydsPJ8TB3n43pSXP5R6tS34xPPQzkXLzd
gZilqeUeiNtbqgRxZfK4gCf07ioZbuFgc6DkRCORqNlHx03frhmHDprVsHMZnqJ21YJIChRZ/VWr
NE7KAtQTRW12yGCLiKP/Pvb/YiR4vVpBE8LBsuZNsFmTsy2kt/hQjAvmlv4Fto0ds0lGYf+BJYu1
se0FDGYd7ZKJpNBVrecH5JSJQnC4nL//HG/e8GhZvDdmwXg8fVBnyoz2X4RkpNjoha6HeySxarLd
a0C+eVHLHvp4FyxbBny/Eo6berbt/5EaLC0apVpZ2Sk9/2XycGA0lEW0lu9BVFmdL168hoGF0bs0
jPt7Rrb0gTzcWRUmCWmsoPCgLETiFqXJlIGP69qlCD70kSk98PVjQGcoJ2lR9ZH+ye3R9JTfGlrE
/LXM5aJ6MAO9I6a+GDY28ojaI7eZeCqbDRXFH7gPY906MUDbmCcplXFyhCV4D2NMz9KqYKea9TKu
cv4ZiuRJb3MHNpreOAf5LCENSr98xnhKrbCACVq8+0OTJmWMs63LsmHgw0k2IKgm1TavWzTm29kt
y5FyhcuiKEF2gKi6Ewzdp/uX1CwVo6oqlMasiuwG0EwV2MAifH5RDh5/C3h9JklBdVjST5+Rjgac
GmkMmq+kS3+zs/zHLgUgI93CxVoL34tW/dVW4C6c5Uf9IIVRetD8y5IraHaJkV4qM9/LliOXKDoX
UtsfOE7461+Z1lk4GXg+sa062eub14GwZm1X9xFP5tDUlxbEdl+nj21hLjyhonwNE/4tJd8PW9CF
RzG59z6k46FTdjxqCVPrOLI/X7MNEXUI6lFOszTE+3hlyOvCzQ4jPe5xkUwa4DcUHnspeBBrn8dr
YN/Tpjf5RdXWed3ePkuaMfN3Iqi1b6NQHGGdx7y2jwdK6WLdf2TrJtfHpNfABimnrm5oCfnXYBMQ
mWKvWBHNbisNOqd9G/EjnaEK2ULFHbv9I1CtnzB3fsKrWeFA7nraJRdT9KlE2dcAjqiz6RKNu1WA
DakwmdVbOllDJ8hvZgPJb35nIdyhEVXsqtC1P5rhIaTzajiMWG1BV2Vo9Zi9RtLymUyqKSznGGVv
bdI56+SCKpbPBlEosMM6gx9RULp5vo8XDxDWr+fkgxbqyUbpvYuu7PSibpgSc+xEaIC3K2eODULq
uUWtYOhYyyVibPXq1jMLrXOY0+WiAq931wC71B+90No4gOyQdHcVVyu3KQktBlQ1WN6FjAiPaDK2
Zh0VKcQAEdY5FbtyVzbhOq44P08aMmC2EF39eodOFu21vxftrF3zL7mzq1kcq+KyOeZsE+YUWHol
6jF2TNvEJ5IsHl+1U6PRvOHmwJhsVD0/t2rNZtJmMBZbWH7ee4gDLEZyD+HwDqJhYl0IpVUqaAGD
wDBeUtDqRSgbQryZCPLjPYLS1zp/ea4QZhMgrf0wC+aQGzGlb1cU6DDb3QufzY/5KXeyREFl8Y5B
cipyKaYuimoA0fMgIlvs/sM/2yKOwHN6DMFhH+zM1gbnmL6Bp8Cgyandg2QZWUkCPL35v/wIgkg5
p8HhFVZ4SQKaZp3NXDGJtFfs64mRAUt0EP3qKuzqsAt8J9sIyqwEC1PNvceBMzrhcug3IMWi6Fvc
adeReTXsPCj/KVH4KLjuDNC5eeTRKaKS+oaw5W1XS4tBtveUfzpds2ic3TyIP3hnyFKDhZVE1XzP
OQ0cDg3l1zpwxXV8drJxSmVNKUd+U4/b9P6xiFZ9aG/LGx9yYOhFZotqWuq3CQcb/nVEbwflxmH0
HxV+bOCjyiMaJp13Uh2KJ6AkHFFLAdE5qtBThanC94yteAzP7oHuzpvTYs4uTwcGDoKspuX4BMdz
QDLjGR/5hwn0DOh5xlAASXG2rLHreu8NDUojCKNblOCNNc3ahLh9tr+etMAtUP8mi3LZP7KBHPo1
cUGJuI74ElO0U4RaoOlhlPmyLlDy75YCnoVwnaesLbn8Y5Bmg1nvgVB0EeX5TW8p4tSDsaMoPpZg
jiT5ItjOm7P4/Y7xV1b3h30xRF4ut0QzBwN5y3tkxsSrNS5/Y/lUVfeFYOmUfOJVUJHloVIZu+E5
FdiIsgCoLA7eNpFKrplZlDWbU/FsSrSNyURzOzpbFvOAD8TCHw5j7ZxTJcPYe0rWtAT9W2QVIhTF
9SReoM4P897JdyPDGSccp03zrlgbEFNVQp43UNEtWLD8G521w5KTQnIAjbx3Y7rxagjYFEOR9RQL
7U9TJCXLPXEgl40r6enDq7JxZlZIntpkV0mMWAVOTXczCakbZvLN6hYQXmVdGy+JpGjFnlWsBIc/
q8p0xk9gT8xlY6sPrWpOnMzDT1BxCBzEFDU3aud3ePE5kFgcB1hdL9mCOwTTKJ3sAA4x1bcr+9sM
j/Cm5xmhgLrVL3k0ngjj6i1L9KparLgqSsbqcWONFxRw3lmCC/UHGqaWYtaNoyJYXcMzQQ+j8Yz3
bnUHlYV7UraIjSCXwFgoA96AHY3NExCqCkUlAAfpwP/U2WB5rULH3JvF+JmrqFItr1zcWLKGBnTu
zTDMUHgHf36Qw1T/QYXI4aqf9Cv4ydaTtzqr9TuoZ4KMzVhvVejDqAyZ3BT0zqnvOivD40ae1JO4
R6/OqASrm3vmtIU3AyYskS3QA3Zg7AXZ59O85ZcqgahB0MXzd6CoeW4wqI0ow4nNVZg+uf1f8eCG
/HKfugHbVdoj4yU3B9NIpHTDK25907/zGwsUC4qJhtLRpEGPAFgbrnGZU9xVml0I3ogMcGV57FZ6
a9hoxEr/Yuv2Ro+q1F4xWYDq9m7CugmZo6epAvCEw5xjSKBC92FffkckCtK5awUJDoZYfAsmTjsL
f00Vkh8iwDoaF79My/DZMwBvbuhkmoqqRw5zKv9gOLV8HhAUfH0TM9BorHc9TSvGe90CPQcl460M
bK12z2Z0y9b32AS4F8JqiEAIQpCvRcPiEr6sZAaGG0bnkctPgygM5YCJJXuAQWOM2QAfjgJ1vDAe
HlUxyfpv/qTb7RlqRoibH4l4Po5SPia+jrjipH9+xFRvab+7ErvxuhHEZqtPPEsSrryNbY09U8M0
KJJUbh/iiNfyqlMZOpgqkclcQiUUcqwn8Pkx/htk7G9fIvcvm+kgoh1KuXqOmyslg7QxO/h9jREh
1ktJiZbDHpoQljaGgAMRsRdoul7NZpayn5lmXKF4pWuvF4BDXSEmvYzRXRCo4FGWW6yH/bhPDfxV
DeRv6r8gK0l9L/0/2M+29DBFOoERq+NVsoIX6QylRIQ7nY2pAw1WLLXA7tSD31Wxs0E5Bl3nKAXv
5Fvn9tgAFqbtaSqAIfC7GHQINpvE9eqe362dIpmWJJd/fhoX1khu8a2O6O19q2iOvIaSYQLvamYI
SCX+hsOgYrNr2mi3k2IR7ljjXaxXhHxZTxaaC2CCw1ne32MhbA0wNtreqpNOx5tmxGBoGG2KWPAZ
ZSbhw+EDFiG6YOFNgE9yXjHl257gdECS1Ro2wTNH25YB5pT7yapZ6kbr2sEXn10mFmYKtioMhiFC
TNU2DCQGxR/5GW7sqC70XnMtpXykXAUmuQBig4OvjJsudyx0K1UY66vn7r03KbZtefGq+Vtxt5Be
4hxr8ipFljy1fErImaDpjctsqKLpFGKhOqgMu+ewNXk9DETGubpjyOQKGCrkFo5KSHe6y7fir2If
88DofhGx9yDES/iWBD2Mdy1KcXj3VYFhXmQcJvmoFQm6lQYEuZ7QNj1xL1q/lhlcorsp4+dOaeAh
E1BQUX8co68eW+2sIGmR3ooTjWjI/y0NRkBZV8qaEdxIfsB3BEIiDe26qTgbFmso6nB8cXdKbDyw
9btmG3mMCNB3MFfGOpL1UeV2I4JzIGnEWD7glB90aPo3pMKwCdE0a+1TKPMvYAvJ3PIcqVuERPEf
E5+muyAS2KbcOQmO7eymlaaMmq+5YDvU9hs97ykO4W93pbMU3YbZPCL3tnPccpDyIt+JoNzE+MOe
Jpk4+69x+rs6KqCkfIAIo1KTRIpSPf37EPL472IzhmdxUSPWs4qwCes0Qi3gJR+mMH73ks4KbGwv
NYeQeJ8lnnpbRy350ihc8b0XyXLyhHPOwGuKj6VaDyPuhiY5L6tYFouM7HYIc4YVaqCLAmHyx/zT
4SD/SGis4sBvXitU9f4CnXbNXB9oZOjYaLgj35SohRqmhNR8yr7+65eDcM2xxeL19kAH09oofJbX
VA4zO0ljFK/psBfErhkdnz9o6FMvRa1r6wA0Rag0m0YjqIS8IWLoofUwKbKQgJYlZuQAwM+geH+J
DZwqnVBcH9CvelITRsycnwNDc3T7zY9kwe4EuXjtUxpqIrUSBs+yV1cwZuQolZbwHInEV0poxmkM
qWWb0UfNJ9QSZAWkTm4GWBaUMPnQ8ECwXXrt0ogIqutb7WWOJKErV2uflnAf6C6jCfDscsLa2kGz
YGqjIPSIJllFs1e0axgkYGPG9x4lDwyiWMNqg30YmByJxSdmlrvaCOfB6fPba8IJSqVBAmwqZLcv
5Oh/SP4kccPcXZdkGVCxLO3QUzOo/OS/3Q8KoOglXJ/pcRO93cv/pg9mM7/t1PaDWmJlzwxhNF9l
5mh5Lk0JbwV/4w3mxh7FKEpH7VwPWjUAph+Sks7z+uY4MN6YeKewG7ugIuFFRp26yNJTC0xgHWUj
/TtfgCStzOSQYscXkmj1K6ESqeJvgzyeyAbt1N6AukVNGLxQm96ZfRUS6K/0QWY74UTgme9NSKnO
lHwJD6UGZiOzFNZMtiLiBwf9Aq44c03aTaZ0NSyyU0sk0G+bkMqXmb/082A4mSm02kMhe/CBbdGb
mjnS7T995xCDn5vgKQ1NcX/7WrOtWyU+O4rI0b0ISyDWsdYZzXtFYUkjc1NdamYwERRnnE+VBBcY
ma7vPmpYGkByWoUvYgyvkNrvanMbEgwTD/gMD86BUOpW8ywgW00NQy/ky/S0e8yOZyedVO+r0xOb
UP2PmjXKdW7WYKKLmwSbtV6o6jP+yfPdcusiwMEetzkk5O6qNe19WvsaCaSHoWkiV/Cn2EtdNYXd
51UxUmDyxgfJ8aJxNTxbCC4prwbRpm/D8nE3OvjL1fiQrc7E3JduInIEgTwj/cOMA/8DePTEkOje
fYH3G9KsCzh1fC3JyO4ac+4hNc1RhZuzF9E8wjMorpfRnGW3hId5aBdkMcxeh7I4BLYV5nvlJcLe
s1fJyrYZzhgkzlMJJz9GnfZgiYWOH9sN0fTfjA+HL6+DoE/nPZnPhmr98RtgvUV5UVJ4JdpeEXbD
cEuLcZ4PuocAiSj1WQEGu9hBAHUmr4gP8kKHl/xO100EEtQ84HdZoeOo2Z6a4S0mESjAVkpOSZIv
LAOBu9z+lC/ggWnQKvPCLZdBy/AxkHCDp1vWzee0czLONrc2vXw9JMYNGsXF1Svc8EoVIayxwWWP
xbaI8eJhyq1DWzrYg9S/0YlBI5CWfQ6fdX66Bp6CRjs+c5O1nAuAQs6LiuScHgL8b+GCTPfYvPng
3F6p8MAoB243HMbLKLsyETJF40MRvIvlbuqx6vdZ2PTQn4VjzPU27pTG+dH55cBsS2INXi2c567d
mR/uRG5kLZQZiIWsvbKacFbMIBOBm0q3znwLFBntqH3Gii9/ssR1p63cmK6cOXDM2ojJh//N0HWn
X3LReCGr7eM/f1U2wZsJUNNDbFYb9rFq0rTmpn25apwSwVMeoEYqDyFts1yoYtkCgEFwPslfnuYB
PMymPEqHyPMOmrR9lER9feQ7i8z+Dr2NmrDP5S1iBNaSYOID0+yOcCj5A+b8j4+lH8N9fhDyj1Nj
0EwqjRTFy17zweYVF7DBS2be/JCknEc8q27HWBFNSW8RGCavpWIBECCwbhPk0xZLP2xn6QbfS1/a
WSPc9nP5oteJxFm59Y6PtKVk3SfQVn2Ry5whhlMGCL6e21jDGTfVfvnwFtzO7RsdcV+qqOP/k6tF
h4pB6G55VdAwDGFyg6fn/dqE4Aewu84T7GtHY5UZZkmu3+OCa+qwmhlRCsbx9qJkioW9u16aggwF
FMi0+bSYThy2sbq23sD+5CmSV04VFqzC6fcpKbwOKH2IE2g0L0Dg/j17zxnG5slsrkyRvnnpjD1F
W+b1F/usgO3s5+H53KtcinJoMcS7fbPR82i9os1Ss/TV0HbIg7nC/1PHlyfk+dmHxgYvBls0TvRl
At+xgtCyEV/vR5NbS5assnNOW8vMu+sPoOP1DL5RM0Hb8n3a3wlxPKSafr4xT/nMiMecFj/Baz+l
f3FFRinZW8wfbbfJjMbEGwiUJqmS7z3gVlNRfXM+FpICCnM22gAC5G6IuAQj2Jbviv8s0Xn1yej4
A9xqgEPb3KPBo1zWK16wRRGvC6YVKtJt5CO7EFBiO1B6zA71HSg8kXohRAvdE01+g9OQfeFSvN2q
wd1odxqmzbF1h9R3vXj1JRoPFD8pDA4fX56V6Ytyd9wKF9ASMJIG5RvSr3alaUqSV+d8tsWCg47m
96NbbF0d5gCrIMZ4DiVSE2+d4cXRvOmhJME618Im4AcdXud6vTUnwT0/NChTaUzqyyBFh7v3k4G7
kUjDvVMeho9LYJQpOLQhJwlN08eTpYuiwivbqNs75iv654bN3LURqxSBVT0QgInCoP4biz/mLWE3
YqRHPVWvEn0qHAFtDMEJ4MyMfn4QofWZkCU6ggKcwNO0cVeXlJnHSqhFztCjmmHibOw95wIfVqBA
ptmFBb4hZF6Uk8fY0Nshth7UZV4cDnEQb3Wsmq+idLcAIZuS2N/O6j0lLlyjEG5iKw+XOHkCFyMO
dQFoekBRM42VP2DRLFoUIGUADkb+dvO0ehuEis5whzIdWxC/rNG7vCYZarWIbGLOxDeV4bN8AWcf
3KxpX4qrcXx3tBDRVZIScr7D+v8jMZaaUEwUY/xW+3yIQronhlTUH0JQ4hI6cDRm25IshbMIJSBc
vZB29g8YZRb+lUUm7uBCbS2w9LlBGlBo4n8CUMEVEYYanbRdhaToFCxLc41ANirJ0X5Vocz36XZc
AhZHcOFAdA6cOFBXY2zsfsgQJGw/CDNFuGGG88Q7w0zCVZcnbrBfb5mYBMIcOBL0NmNcfH1s4iAA
dC1ElhysGIPRztjlZvh/MRoBiW4J48X45/54VGRbeVAm+En+1Jl5zdaoFEEKtizl+KRqaQ2orIir
jsBgK+cBQco8SYXyEckVXWiiviGh6/DoIQT121t9N0i1MS4jJLEQ9tCT+0OuegI6erIWhKMUPVs+
6m4vuZ5gLzq8JAZedLUDiaFNiddQ4wl6nhENeHf0zUHyM8eWOvifhalfqFD+tS93QSu+rIojcsAU
ScbZ5bCvcj/GkzgE2zctF+gOeFPxS6s+YebjlGM5M//hNr1B/R0OAC2I4lHcyeeTPMy3E70O7NeF
dKw/Qjd1F19pr4h2V6J6D3UMwAsaVHtJMAyNO2OYReblgASaJBpdAUUJB8YSnojNYVKTd2svHbj0
ocuFgbIyIFI7/U3AU4qisNTmQPM2IaTOZn9TjE8YRYrviB/1wMVLjg4YQ5/NLN0Id8dfAM60I9et
HEmQLHyqY/VvtNqQYMNQyUNDIhmK7wOzePiOYdm7JDCzkfV+M7mp/ugm66MipiR3/0L+qyoV6ora
la9Q9ncRObBWtTtTfLVn3XFhmHkJUydxJ3Dpd84xq/HQQ7/NYEO9seqVvtpSEkoHeGwHnMU2LTPG
e8+Z5sdOCC41X1hfzDIAfpD0QCOJucBHF/6UmfhyCbzGziX7G3dFrHDBy1jST6PI+iE8fM/cypUf
0UMe+vkaIKxQFHIvIwKc6eWvwgxDhtXmkAIHoS7WuFBdXQE9qFB9ybnRj6nBTV3sOLz8CIdF8YS7
5NfMXW6uBLWkyP0oSDG/cI2P2sa5DHR88R7hTbWK+8k6AmVdbRa5DWqAMc1ZrEIVrwnNDkTJ87F7
EG26Q1bitlfpE8XnZ7euSZ7tr2hiNnMJv3CDJ+dmqRCXJvi8hGYgLwBe7fc4/RcXQ/0HwXGBcexQ
qDxeMAG7LaC76Wy9sfiufF8M7rz9Vc6/+4gKbOaW5eMrDPpGIqTL5iz2bXOVYsT2/91zPmDMIWPj
jPgqGPKSkCgytEj0Oaa3nzPJqf5LbPLWFCD5ooWDgFbVc19mHCwSlWI+0jvALVIK8l77TBd4d43B
mZdeE5ASFtYyOkutIWtluRFXvx5bqvUUwaUSi3CMqfHUmYQZsFBGavtsf4nfak8NNNADzmFQZLwN
D33FfoLwRl4DEFUCbgN0EUEmX3wrFa7wurRqM3H9fZ2HnQp44k+lkv0tJ6O6uxgeAZ3nIblz+DG7
IdgDcVVVBVDxW1yjhrcnbMxLUTHI/xqQBXoTYlsbtuRsy1IzsfHLocMoBTXorODJDeSZOZX5Tg3g
jb1ZBctk9LiJGi7Jdei6LZXgjShqaKGI19Rgu0+18Nw5qd6aA+PodQo6jjTA7RzogoZijCYazaHN
VngQrc61AM/lQIT50pdmcK0OFWwtPO3bia7wgaWs5kivgF/xAuuRBRqzRTfSerCWhaCzAUIakCWy
qLpsQP2qqYq49yRZX4cw+p2XvWozPZhj8Sgb4gQCwEE+2H8GRuiRjSxb+VRKYqbrPyp/ligNSQHM
eVxmoTfLYQbPnjdJMkC0LOaAQUZUKKIUn8KCDILP1j4X7w9Jhl3LMAFedm1o81S21is9vGUJb10Q
ld4QNdzsHwVYH7LvtlSueI4K7GEBTaU0Fwdl25bliUF3oxIB54VVhvPo8T6aPZuRWlMj6Awco5s9
g0sy54k6TS2btUdOaev06UnxHMgeCNWNFCm/IEkJjcDrn2OYwd6LaCCcoK0yZpZJ4d+lIhOKh1FE
U/dIwSRmuDFyJgPlw9YdNtYegP7e8FyPpmPE78eLbJVqVeqs1QsvHV5aWS7JcD7Fv9jmU6B01Jqn
NHHkZ18eEPnti2ICIyEDKemDLh/J4pSCBSaOdXmY6KkNdcVwdpW7w1W8zaSbepcUp/Lqs4uk+xt9
E8gvy++6CJeYtnlP8XbAOr4C1ZDPghfmK46imK3NlUqi41EVNSVPci6+5J9s3InAgVXKtlD8+ana
PHvyiHSVJ+M0h4wDv3aA2uSt0YqKZLAZrZo7ZWFeuuXvCmpa527sMHkKc8IbgmNjF/zjUpgMlYeZ
S2/z53pkzxTvsGQI3lRdOkVeuUrou6E8duTO6ZAmwPfGjpLufSODTCUpUlWznkRTl88g5EOM6RJX
W0EHth7HcMjP1U9B8P2qFaNspmZItqFY7x78+Wu3ayVAsI6/lEED0i5Dwgvkh3SLTpJvzuUFuKKQ
A86ZywmHpiQUJJCsWUcs2izWLE2ojL+lBW/S9gpS2nop1zYMEwjfLSxVus9K96IQO8cCnvBOCwhd
9t0QcIsaB7imyKLnwkZriAPbmoQu+0GAxWsudeb4jH7y+jHK2MjRHljfWTae8KRX+oD7nT4n+7Wj
XV7fNiJZ5tOkB7n0rx5GSv5PMR8bqDjo4zwvP6hbPLyqoroPIl6txxse3g4cf0PuQje4YDk9KA3g
zDZ1tHfm19fipSwKR+YAm8sJQKhf9tMWFJkjImmaCn4h3LDwGpBNzTxabmX0MBjmrU2V/YemK9f/
8Nw6gc+Fx7qQEZuwsLw2UigQ9ykTM5vumGmQ94wK5dEbeyeo/Hd5bfXi6p+qMJkC54dpOrZSVDYU
QWStf0/QM2eCl0mzAbDogfP3EKlW16hX/0OhRkUJ9PAy9kjN4zdL7+Ru0TrjnWSnWC7zS0reF8Td
8y3OlYAb6ynxNCK0mmZFlu4j4MprVYyGQEX8SQjde66D0JzUj1t9bQdAvM16o7IVWwTx3XGUSodE
lHsi0jPDCBxND9PBMb3BZkqrHl7QCZaa3faiCFW5eu6LkJR3jaIRIoff+pwe5HfSLgPrCGWt9vo3
k04pVTPh/fpSQnAWgo1+6MHn28vW53rs6z9JP4cBSLT29kBVGZBHf+yWIzVUE+dTY+vRFFM83CLG
MWh++zEdUvs3l378FpQj08Iq+I7I9MbKsT3xBhuSXEdlMyM//2c9wLdDB82pdv+gXVFMJ3vzlGCb
V1cCEtrqtokzt51wowxZLqsaz03rXj1CqlMqd6hzO+LoiE5NSzg2dJ07TXh2fsOy7/sJegyo0xTW
cbJfLFeSTYWiqa2+zC388o2D4T/obD32AilzBjZkDqZMU8KPmhAIncNtHt1SG5qESr1CUW8jViEl
+6sonHJQ3YXX7QmhDoT7tIyslX425Sto9C3QXsDON6lwXeE8qzcnNndRbjYQZhzgEjvi21JXck3R
xUDwzlG1gmiRTZx0e8Bs7X5JxPlcYYswAq0CxJk440NpevWx0i8gkcs2hjT+bRCA+ksIrm83zWUp
zCXYNJ/j0F142Ob71TE8kuD2RJS/gziU2wXXJTxtKjzQOZY6wSiulSA8BadBCIUUtOXHWFR4PZzW
UlDuutA/KQxJf0dxdvHBBEPMURSMbbs943DJv3q9ovVVzJdu4JPJjL/YwzlrdinVyFJmHpX+cl50
ZeKMSJz6s/A/UyUe+Ujo1rrDYOkk6Gm3ufpOIYYr8N3FIMbIwtgIpbBn1qSfTFCjVNu604MVODWv
v1p9HBlXtkiieeGXe4uvw9ALm+kfKxZlma7K2IfR1wHbRUWsEa8O5WWmTKBIwvbLVK3VG+Y5zQS1
XmqUgqCKqEEqv3iYZg48qSbEAvhc974oS+FL1rwHc0c8gLDrIXelrX9heNtyDd4NVPenVbSmNbGZ
JDoqz9T7TjO6xx4mhghiVvMmCLGZEQA/CVqlZLt66X8vaQDhNLFxaxz448gkV3oifmDhHMuhCkB9
eSRy7cC8AZp7pTvbNnWG0G+NT6vD6Jz58JA1b3fORr9u6D24UWmSn22ShRNSNWNd2k/aBj3xBSQD
inPfwpICMax5AnElecxiPVy2JFG693PFostC9nLfJYQaWf8ZQ5R1HJEy67EfD3tVmdrxoRTgXcW5
YlkFooqoZQ1D9hSqQEtPAjLzpA8MejpfyENarqGU4zE7osrJLRD021B+N3/ys8eYwXBJCsvHzz9n
Zu21EMsB9Nv8oF+6e9JaaWfNs9qQLGECE6UlCvOzTOJ5fj2ANDxgAvawBtsK1G7CHqSUpn8SrIWm
ubloKy04FeMLH8aoETTl6X89kJiOeV1YQ/pe8v2G3GlxGudXrCsAMhFUcv5ATl4rRfl+iSJgCoSf
tWp/J2Lh0DNuwVgCNcWwtfe/st8G2oXa3tFDcDvtuu/gVqR3DEWHFHVyl1YUdgi7D4xg8ePaJpZh
wAkZy21Ty1IOV8FTVWrYmZwlZU2gD/RpXEJFreuVrPTQIWUOSZb+r6vWyy6mNnab0CbLdNtPDi9W
BijF3j2BB/GVbKdhL/wIWQc+SalsZ3Bn959B+kefwUv5Xi9r5dqTpz6ES3noWmbtT58iHtk2K++b
QSTLhP2MFPX7Zq45wDOw0Rpj+HBEStoW4TfWD2982DLn6L49qRbbvLqO+WYEeOqgLMkAPrK9E70x
X4kR5FCCIxfK/833qH+Jt0L42neVdKQXvCy1kUA0ur7QKW2OCBb2gubhKXBbMYCZjcN0s4rQo6vx
SrOlKmnAjBls6thOcvCspk63/xLy1cY/PcOctLbQyDbXHMhvy8XhwjGogxZT58rQWoQejoBwDtej
9g6/ky39mp9QGQ9E2AQPf0S0kd8cNx6B99YfOxvPHpRvkdakmr+FhlixGdXt+5+Zcz3Par6LHzyt
/QSXL7pRnV025bt7Fy12vMKbXE8bIEBm4/rfCc3EsuSDFr6HgxZSJ84sgj3yroENhJQDN6wMA8Nx
5NBLip2sFH5eEJheL/E6kmcfXBjsluf3O2O0kysKT5HqlxTwSPJsEzJGn689zAW0PiV95l0Wvgw8
YdSrXlSzHYLzkNlUXtZuwKdZSuHPP7pEpDTvC0JwS7y/lUtKK38q2ukozh1iiGjKy17gkkBSRQWc
5+egPd6JaCnw4zCGCS/phUMel8Jh6KFcTONMnNkJU+xlocAc3TNafXx6TMy3/nNsqFX1ZoDWeYOr
yUH7loi48bG5WDuGukK39bMU7lAZ6Qn04l72Z1DGwYvZhJyUq+dRTWtjuBSrr33rebFQ2JtIvOLm
2mdNpLSq8UtfFnMLQdEC7jWQEXV8h0R0HoZeTG6UMhhQh6s64W0RUa4lbb/YC+Slc8DAJVo7sqRk
Qn9QiNmHeRh09/E+414R2Q2S1teCcbs8LC8eBxEd8AuANVkb0SoaVhnAjahYQH07QGiroIGYR+g0
bym/bjWYR5rFTlCJoL5O5N+75jFadu+tRQzkUGbJ5AnAwtyRmShHQknCV15r8O04V/H37gqLPWaq
IW1UKCo1WupV75cHjWn+3LfRB887BHd+E3D9HmhtvhWMSm1N+I8Sy17EQdUJ8y5adHm9N/RpumLA
i6DrW4ticLHh/zr+fPwDycDkrNbcgzw/U2pM3bSgJjGbxIH1cXIOHer92XULLoMK1ccjyDNacPeU
pn+wcNu4OKBt5Fb0iOxsU8QJOK7w3QALo0Y5CSnn7mfyNymsizIyG3iDGbnH4jJsbQBTxmqca7sn
0zmurH7q1tlXE5XVdUibmDJPy6y/pOVQxiQk72jAhnIjXVPListJWtE7XAxrMpZXJFcRUAvkum76
vsxeA+oFdHTJBRCkJ2clXJoJyGh1K8HdYCTJQkLVmRSkgIAWvwf845SjhLDiU79fBGzuNS77Sog/
xlQ9n78uS+Upo6s97py6IsCGNyJplkVQ42lraND0Rjy5wzbu/+7X3oxnvOOu3ZJPURWsTFdeNXj9
R5vTaj9unwpEF8Mfb1271GyVb8DF8kWZXOhNUpOfL8fNSeJSTmf+i8iUwl7PiaFTkemv9VpYyNxd
045w0R39cl8CW/5z7IYrfFuGI/uw+PlfeTJnnxCDrQod1iZM6N3NeduKYmLvEItAhgdlRp6p3e/6
zA13LTJolMFuCgd9loHgU12Ls62aZ7CsQfoj7EsUxnJx/lBWopU0V+Qhv1rh+Ifn/cBsUgcl5GZP
DR+juqvx/5XGpR7s1qEKFrUB2IcWcTSiPLy8bqqR5NNTPTW1ScB1rDwTuGXbXp1Hi2+k5lCIT/Ab
s5lL2H9b+pXxKWZh4+f25RIlTPfsBGHiwK26Hup+JIWneA/UMIXMhFCPUXTGUjTA+tPBMYS9+dCk
ShZM0Co6PVxBI0Z9OcFwWn5Jf7IZi5a5dOkzui2aEWlb3U0D0F8FRJ/IRv2PLqnlXZIh0VjDHqij
er68JhvSrkz4pFn34nppSewhkuwnVMP5RF+LEYoD3lzTwHYvz7KNgkJkDKcKXt0ZfLYa15WqUfUF
VNC5PQLPOKvvHS4ToZb46qnLy/azYGyZ6P6FzIbTW+GlVJIifCjw7SqoEgt6PJTQhzmpp9aXLIK3
aMAW9CSvVpw1m3k059rAJgzzfz8tdcGFVYEkdyXSBOvGGZLKLtT9XGEGuCDfsERqSxGzOT2IRC6D
TKq7mhXlYGn2XZew8f9DIZBan706F24l132B2dPKh6E7oDq3yK6mSpUDHEfD4TxQ+MXeGKh4ECn8
5r1BJbLlkTclevNq0VSk+KblscZ0V2lzk6wJpocyQH0a5cEHE8rZ1nIX+9P/aqSTLV2X5T9Irw6V
wfC16A6rjw4n1F0jgHDu1COqJqsnCfs28E5NFYgixtpjPVhQ8h962LIRRA5SLgSnNOoWMnhZXR8q
ErJ51vv2Jp7eOMtCgvKE/AG6xRRHSRaDF5S1JAEyFsIGS7ScHpoj/fa9Ko77eU7SdtEQcOl01Lbz
10l61NLO2veCwR/cebOfwiaDaC8GgSfF/4oAYoBeUeZKDxZ2C15lryd9BbBnbmyPBBEyvgC05xBm
7iK7SN6seH+gt58ECS5kLyVoRQWQHUWh7EpPu01qQxIBwJCNPnlQDfG8Jw+o5W+ebFqjgdhSR3pQ
rS9wTparjIAxF6xRSJrlJ/RVIhiJyBleVD6AH3AGovqK7GJ+o/H21wmcQl/ECrQ+7Vj1AMMOVAh6
MzGP6m2PxGgVOgbvdElzSFn6b8FqtLaYFFD9KKqdJQKKKYO2Jcbh+kpCqO78f5FKMJ/RImMQMn8o
IHIy/pIDBy5P4pi29+cXhLUnkZ4hw3lgggyVN10BBshH78fZmAC7hAFsPHYXsgbWuefsS7cyujLE
6Z5LGvNe/LD0csNxTTOvYm0F9yxNTDF50xvr2swMTV+b74QDHJtlwaZCMbF7VpoT7+DgFiQmyKKX
4wd0+kqBAD2AXuc5jv+/yv8xmbPUVM9yTLOQJaYc0/7Ev02G1PjUzNMXV9Llhfiyv6eOmaCI8mv9
vGU1HlBNoN5ul5Gro0zhxdm/mwKvl4jhNcKyPU6HPG3d6mN7DPuWcw8uSM0AXOyfOgUnay39VS5a
c91P2lEIEXyLmhFSMUJn78MK6hjqatfDTCLRCz9A/pHpzY2SKQ7qfYd3R7JPI5SDKBdRhYz0lvMi
zSRGXyM0oYsLjB+cvljcHfJJ/r5MDTju5BRjsagiqepi5a1yjeGR+Wf7cQmppMbj081gh+Fu80QO
ptvUo7k7/opoNjGA/nOzfnFSL4Xl38PG9k/CGtgZx3Fdstr1zk4LJittUmNRbiI8E7iUycviDpL1
/SvtA9gLTYSAs7gu4b1WZgDbd5wpBHqUaF1joOY0WXgrKglVJV0HjFRkdzvvXRmM40NtjgTgPSWS
Pk/tvO3X+Y74RaqL1bx5QCRCLLjR7ima1hgEuHOYvIDgRxY66Jwn+tlFIt6FhVuC3kAAvWY+7LbZ
hzjVcPO7F6x5YTrqGTwYNGmRZTNKvOSGKob3HwA5wjrQpXdky4KdrDJ9IvLlYeLaG85TiQn/nv2J
44iBS1w5ToZnfJhKrHX4Hs6vfeETXwW/ja+62iZbPB0XyHkU1ifQgE+SZa2MfY8yxDHg4xX7yyrc
o4s5xurQqQ4RzX5SKr7dSCwfGhX0Ni02Y954kaJQY99YTieLambZ/bSlBs2vyLCyA1NRIKbd49fQ
ZXiVZgQpCBrmY9KQdJ/MJblxnxECzfmDbfzeXuLEzd5rlFrKKGV8qr+FlohTwBxIqbpI2aZQT0sp
AWyu7AwYGFB1fueNGRElU6tW7jPYtRGHlrzAJFp54UmowC+ykVwexerC1LtJ7CnL6Ur3pM4sms2z
1k9InsLBkxuTpw5Egw84jt+aUhsDemDGjALghI0lb2LLsog/JSXu5vZRH+2CuX4yQgdarqPl4acr
J2utN/0uPG2HYa8hMy5g6Xd+qshfKK9KjI8C56TfHnSla97/WTTRPRY30s9KAaE9vaYj0A5anzJW
Y24lMt5WWZ25FuXqWvr8lRY7A/+y1ZmzGXeyL2eBmfz4llKKXm9vq6G0I7XvLkOQQFf+uji9X4Kp
gaVXyZTbk2xBuR4WYctJm/BDW/RRrJuEsCQjCbGxxMl8MXUvcE8tU9gYnuivPLkv8e7eYTsEr20M
H/lHNij06D7GXLWdrHFRkVA5pCK+JUJqZVLn89y8kY5p0GMV491tuqVdZnCVdt32yWiMxt66Beup
FIgQW3WbIr3H7M53u3cOgTTdk20SjLrL4Un6y0JPh6d82SGfpTmInBPEITNPvJgZcZYsVcC4ilnV
GkBBCisZjbnv3fU8VmUrxQS/3VMHSqddNImAkV/KElUeNSr5Zz2eWamL8zlQ0axkcV6e84IZNt0H
k6RZfAdq9RzhwRkVZE0yibHn5QXwjyIZR5DIogVG6B+5aVUcnsuy1xkrCjw1yn/NJjZGjvC5FW0S
KPBEagTeT1ECBLp1tYyU3ZNRtNfYzX0wolX+YSiC5TI8TUzEKHxw7Xj+XXx2KkdA9Kogylzlb7qu
/Qj0sV7NPfrSfS7l58PkhK9gu2tgvgWTiIpDkxkNL9eS2CfYKutsRRitXo6YJzQOZ93qA1sy7iPG
rW7ux5BoKROLoRzhAIZFTv2DCfkq7YAOCkeFCDN3kyC468x/7mvQRvWRrWK0zTMW5hXy+ZVnWL/P
n0VyGp66ZvoMI/n/tDp8dAjsvCSeSSFY6zAvH/Dn3jM81vU/Uktw8NJRfJ88a7aEyYY8V+iFpDQo
ULSNCyeKvjltqwifuQa0fuHmFlHuVdKA1GMTpsD8CiuE4hVPUULBHaY+LqSTSVxJ+2sEDGbDpUrH
acEJD4zIM/I20S7URegOm3HmQcJozVPi/3uUH+b/3v8f28JeIFjliLrR/Z4e/FbjeeO+zs0NdN51
z0+vQSnkfnG1A58czzsS0F82Xj0WgYKsfyDBmUecUIv6DSEHD0b6uQcibP/YS36iDgln2uWn1NXf
VosMIQ/Axm0WH7S6dOs/HuU0bm1RgPSMCgAmLp8qrtk9ubw5THra7nWCbMUXqephy0K2bLvu6O7D
oTNcfPvR2QbzaIRMoaIwtNzmjgbtIQUaYW69QM2fQO1cEkKFEZTX4DyKEeO6+s9ImLGsT75Srxuc
oIX0vi3ELNOtOYv3HlhUu1L+Vk5oZuTO0xqeC8GFZNlu2CW8HdgTgVghcxPZTmIZ0u5wezfJYShQ
Z7Q7QvkQK7YGqun3LLG16XRvWmj2BNegtAhHO4a+rjyIlMrXDAhSmQeO2bykQ2ayyEDZ5ELWvvtD
sTshrLrIYm82Cd/dxmbNQkTIVpE5CctDctLz+4s8dSqcaBV6zFM6roZdJdesEnJRlefBDAbzsu/x
uztKbaDSyfaC0Nbh/Q96WdkUpoCOIfX8oPaWqCRbUPY3rA9/jjUQt49DOHl8is8raEex48xgDg3q
CEM2JVnGtqE1FliI6SDrL/dpMfwPHgl7YjeNY+wb/CDXiyXPFUN0+VmhE3gd2nQflk3hlHZBejl2
/J2XE4LBiQjgbZq5TBizpXSgj7nACKBpWze+BHW7tC+In1jvwwnRtZGwNlDDtYOsDidYvokj2mf/
KhyDSDJWPiWgfwJIl4hZm0IirUMgguot6CAkJ5gnRFFn0vC6Kmb/DNGgc55Wmw+CDV71lQoyA5RB
4AdnzYuMmlxTQTDMvgC0M2p9t7Rm+KQN5S4ym2p2oUbUqUcgwJkHAEgdIYg31MaEiXRi19dqBHTi
AsfJLj6TD3DHeXmmsUdCuQz8Nq1n9MLu4soWDNhU1qE6bw9BbmX/5rfOlFuwY4QBs1TA56CAFaJq
IwCpctxZ+Wc3FuNJ/oQppD6rSx0xdwWiLngjq/V7mxAbluVSIClQAhRpcnEJ15uAKdBrv80lB5lw
cVg3s6e2r9kbsUUkGmEKWsvVYkd75vGRT3hsR6j5BwBy7aJ3PC8DIRkIfri49HIIvM764+tNiJpH
dY8spSJ+fXT4jP+cxAwAUvzim5Jw8/t7MyDP1UwxmNKojNHQOscHG7Nm6Od+59AHNEtfRtIEzbGQ
a3PcWp+JY7q2aZ1Oojluq0cmC3pzCvsLHR1Jltar2tSlI/GcYxZkcCLZYO3I8/a0+qazb4Sxvo1Y
fzhGLTzz8WSs5z6vmiPuv1LPACSy7mmBiKOGrfQnJHXc4qmZktlIN7ufVhIK8ByQ5ECHX4Om8kwN
b9krfIbgXJzB4Pq+LC9Ac5YORk1T6Rj6Omvmuc3PN4s6KKW4Rp585pJr+XHoZxnnITo4B27vRW1S
s8El+P/iM0qynf93ulGr0ekrgavyDD+gVnAkb3g7Xwq0xgr6Xp3qD0uYUfWBoV1Iw+4foTgwk51e
o8cYLQMA6hk9RE+/79TZY3BBwvJs7vzfs0I2zQuDQTVq47WtGjzTt2W3wMTJ4HQb44wBy1mz+8vh
2WYbeyTvbyJ6iBHX8iU0iy+8LU/wtOMQ+FFCWY5tqS3O28iP3wvxeeDphwlRPbvDNGfke+LkY3W6
EwL4oAGo65HkZ6KkMJE/VVb7fglvp6c3kdWy20eXGIEzYHJ+E8QIKkKNVy1MMNkotkcSr9/xPtfh
s0SFKUJAaFVEYdPODKaSkocCjMsE9jvJ+q7SjW9OpOJwmTArjddatWNrpb4Mcw6MAsBQW+moZnl8
BqTEmnk36vFnq5YkWbqXVLtJC8vswpPuVcDxEAxFOGWEgeYr2BqN1D1kBKLwDpWpiiHLKk6OI4lC
6mLJ6OwXsqPnIbpSWpyQMXUl8c24mGPBEVJwRZhrNHF8mx7oFk9K3Kb4HvWez2Ohe/p/5m5ZNIAE
BV8aUE2bfvDmisD8M7W1DGhzofDQvxCP1Ukq17dxWgqhf0gPgGuVMwwVeTJBobnxfwLTouL1UGaK
t6ALZ4FzliEAwQq9pcxqUABL8NovO/36DMSfMALu6LgAR7D0Mh1Xk4DihIWIrMSDTMLOocWzSKUV
oEQ4xKsgD4wJ1NsrECE6OnSlOCMXkcrdnCxk9yyfs5Se2VcMJEdHMzXNRENXPjKlHD7GyXwEu/lJ
/18BHCQSiAcwBaCx9RYz7aCKolWLRm68lB3dco1+PP7z1umxQhN6zECWJzajwtLenvgs4rCkhOQI
69h66c3YFp2z8D9F/J5emZHbIcluh/ke5SQAzw/MpExZOLyui45hwr8U8D9fFQsyf41G8jS22/2m
mFpfXFbr7tbnb0ocSjMYSRvS0psyHDydu7zAWUxfOh334bk7/SaU0gOvEeGq8WpzgNq2IuPVieY1
lBvniNAvKonEhbDJnTcpDGTFspyDbFUABUZmB6/bYCu+3wwcAZXrgZ8Z1RClQTK2QxYq81b9n5np
xU72OaFycjZuZGjSCE3+KNZaec+CTFzgXYGsNzklbcrIFbkuNVl8pYJS2FKZ3Y1/imJxnNN15Ft6
FKKBchlXsxRAe+reZCxEws7CsI/dnHhhFvCyMelh4zg+I6weRS3YmDonqvQXOr1QGJE3sMAVS8od
z6TcHxy3P9uOxdxy8URn5+TfMWIwKW+OM87j8rgKH9IM90RLh5nfHbdml868wTQ9q5s+mGq4/l1K
/6pKf8KmFXqzc1hay5yn34d415xkME7RE/Q40/VLz3hK5JnnZsxPgyp+g9FsNW+IZUVmd+SZGTdU
OyRKDkM6+gLB0UjKLG+OfU8SpIRNqOsWuKxJlOe4COXZuf3DkFxfyvCzahq8LiOyv5jDCp7IuLYc
cU5F5skMlYBEEDDDf8Q3q9+UMnnNymL/Qq/4ghuN/wOWfMnVH655Q6i5ubLaxEw6vzAmi07mWHTF
GFiugJdzeaO8ivTlfUnoj5x3FWQR3pOM8MDJJwcHzZ0O0sEbyjC0+rt4vHK25zrzkYDS7wzQy4nA
Nul4t6fWjxPpOcuRCRyLX3lpuO6uJ1J+i1XkV0R699HMkX8yJtCNLwM1applE51An7SQfDXDKYtS
CX3D9xE01nSNEkXgeUD2fQRCn+m6GwJlU1A8cWSjR0v2VUoMb0esez2rx6C3e9N0Jw9lKCeufWqF
43PJx277laFvN9avrj3WG9ZBpp43xyIhNEIW9iaNX+yEyTO0E+p2n2bHArJhR3ArLea0GpjH8c+l
b9GpBWCJK6EnowxUgSlSFOr1XFlMsYq0hKuiNVrupHIGQvWgFiMIbG0LtX20x8SALY0cOyIiJPrb
HpiH54v9IpnGJ0o2JVEkqc2gzFanrnXtjxKRSAg/Mw4qBpY359o0jkic/wxSVsyvjLRL83B/qwUY
WNsbMBnf94on+zy5YAopGjQCc79RNlXwrJaQ3cJ0vzzskSkzjrJbvMj9xqBRIVkzj2UScZnYpvj+
2rLptHkmRx/Mh/jgVdji9I70lUfaey4sSqy17aXohZhVFjBML+O6YhfjS0z12pp8EBt+MB1PYgv0
MHAtQ2hqCac+xtvat3obNKaTXNG78hrucCy8ERCUl8x9UgPHyiNeU5G9gyelfrnnORJ1PC5Sl6pK
KMhkY0D7YvbwH5CNOkmTO9erYFBep6EWEIX73+hJ50QtgMEaJuTlsLDSiQx7DidsfU6jee2TKuUt
sAViC3G078AsKOhoaRnmoeeULyydfjOP3bY2/6cdvIqquHDgnq6JqGgbwdZR8U/0v10Hx7ls0M99
lFnmDZDOsR4VvmNQ/RyKQ3Av4Wqi2qKVtCwkWI4kXOrdR556zQHbBFYExunjKggLOyevMctOcV8V
OJBAlV2JCsdujDyCHy5kHO4FEl3U3lepC4rJV0hg/aIOHKEBKaC5nPEieQE3WEPuPEgUUUEDapu2
hq69zzqpXnTPCFjTtxAVow+s60h45A1/QUwZTpaGmDVcgRVx2AIiiUwtUC8hG9GFmFLUz0gIjcxN
h1u0TXlEUbVi0qDiJHlcyQ13H39BGlB2V4AMhoX4qGAn9tNL3zOz9y4PpFMolMtlqcJ5BkUfNU0D
hCBA/8b2xCjlwQI3vFRASd26c8B4iCa5R8ePKDNS8xSnHorgPfVNcIyGqNEiFBSSfqPhCHtKznv7
73XpXHH6ByqkpFzMfYmBJbIAGUP1pFrCSC2kkZc//fQOCXkaJRxuRZxB6nbV7sTV4OfRaJnL/VT1
AP5CgvJMXHUvszm+agQ5YHs6v7H4i7MFTfb8UjCuuShL8IxOwbhCa2KRdPfVZOcjQs+d2BxHgrjJ
2NvG0NA/s5SDBAwPFAlRIzXYqY1947iNK0mS+gMxmV+NfLIwlqdfHCoXCAz43HBPciA/BPZ08Hvt
y1RIQFnxioY6Ca+Sm7h5jg1/qpqXesl9C2zUXkqoquuMh9jq1pb5A9E7y7xQLSkRNepJz5bQVOB6
yHxF1i64eoUJQSobZ8hS4nHph9zNM6iP8o0gPJRMUlHkokV3AMyNjr+yY/NI1Vqg9DXT7rgHkSW/
TRSRexvhnROaDdGMZf8kq8uvyh69fU7kO9d7WK2ueR3GigcQbId/xA340H0JNfndd0+tU92eSZ9d
Mg+w4P0PMKgoUyr6LcEgwca2BJE7CPNXWjDP+ObRUwTvFBnYw7WoDK6itVkPxrlMP/50HUva9C5Y
dvMPaUD1Go5558tNN8TDJImml+gXveq+NOqjBTBvcOkuOsj1T05rtKMfcJ2V4CQq6XJG/gWj7pa2
jeK5HnVSPa3FVcyS7dQpsN9Hzg85XzzIyWnbRe14rQ3PdKASi5PNFxRrVgCFfatp/uvkKdFwuhoL
GfO6yw/oLnYOJEJuLqxGUsGNf5Z29lSScST8pk1eLjgCcv4hmVTWR9NaeogO/qGOtD1MWQvfWg3z
c06iUPDt00BSqqWRahn3tS0YRLkdtxSihdrAKfgKCZv0eAHVoRxLvcIML/vcsaX+oh1QTG7UD3ww
RpOld3OodP6E+v8rWlTktbHmmMxaKV484j9K1GU730KQbTXCnfFu3qw5y728ajTWt0v5TS6uFrkj
pB+3MzrK+14TlZ7O2MhPXaY8Umsv4ly+Q3jb1+jndbl2Bu81ERokMlveObG4S5KXwZSa8NG5DmjY
5GUelDpChYnNo7qlFrKZ7KA3optAFwlyb+r3yr8bP4jYCqawaqoS/fc3hVPIElnv8PQIwvsJKcWG
dpFTP7ANGENLYgKwoAtiqeUd8Wn7pZNSBqTcXoLzTpw7UPRI4MemX0K3PPE+KZV79MMPUp5mHAcY
hc676U2Yhq7uUwauOUm88N1BO2Sufps6wTuvF/XxRzDPv25QLPbOduOO5LZ2UcPmOETJ3xM9OBIc
6brjJ2MncX/d5Z0P1zKsk+s28rWi54JmWVYsFS3StibJd1yPNc4YjJhk/HAf/IXO4FDB8wQzHnHQ
OWl4QYN8F5jw3Ph7qIIAhYpgP1DaQpa0rwBfljw+eeYRaOL/w4CmS3ALyqBdCtcrv1EAVv3QKyaN
dCI7G2DRbnxMTXK851tlt33g7mVQhdGijL/whsLGQv9c3o76mBlLTC4q02bj+P7tDzJ+Hte/gVid
VfgPdgZrkQh1UXtCA33sROO+Sv7BFgxs8J/h4eumqltGjX6r1ndidhjK/c/7zMc7d1guZ1T9G7Ez
1uU/E7vQ8OI8+UAacnJArTixkkN+bjBKDhHSLL9SIwLMRo7qQImturQqrr1Jh96NYNUM61dAp9eh
RkS+OEVr0Lv8/0n4qw+pGIfxJaE4mZ4wembOE39YV8/vkLpwObyedjzt9hhAdLiMfxmb4DvIX3C7
7rFgaPKD47Hmync+CRQSHE/4WpvVDchhQaQwSGJO0fxXFqckhY0kWqRAKtnwFgk75u6SwHFAfrph
ditcbVPJkqR4cyfpo1FY5u6Y6Moxwk6DYBkJXuGS1um960Hh9TwBqLLqfa1MUWjKDR0SMLBXHuwU
Ut2hKiGKROSkhVeaUvc/JvSEiI5FyquCVLmXh1DBbrBEbmHoqbE1nhxJqeC15rBK/Pvy3YeeVwl8
OPVT/sx4Lj0j0GbPn7XL/6LZBS5fPP/zBY193DTUMy7w1hsPsAOWWflS0nVYiKeDDQSTtRcxsgdw
XvH0XPAU0P1Kf2GWCTGvfSyyQ4VfpjdozaEtcmDJbR6+coagD8C4DYH4vqIpo4WSaO78dvU1iwfb
mBmkP/8ASfoL9oovHPxOgMmRxNqMU6MiqzrVBdiQpYGW90z5aX0x7cDLWtQfc6gF+ECPbBlwMyIm
KRnngkJ/C4UAMIVZf0zpwwF3SHWLLVLbtXjYH6yn+0U88vSi0sj0yteyOyORuAU8W/4vNnTr6PQg
Z+B18o0nJ0KVSRZu8Xp+bm0JEG/iebyDHFQScB/aT++soQAD/ZTzYfccME6PadZCUuFhhrS3WT1U
pjm1RKbWgnT7uKqVBTDyg0YyIWH1+h0W73Z5FL69rFOaBoUJ/R/U6K2iyn/xC8zx3qylZJYWXJQn
ICwnAi3Xw4fD7l3GdNEp0ytXm9S4zgjgda8CFNDyIsE/+wIWCxNuvTHrMhg4rlOEkpMybF0L1KWV
sdiO8Cdp25qGWXaElUyLvuHbNTLdh9U+dX3Js7SgafIyuAOtN8yhY2WgXIJOU5dkE3Ianta6eaNf
renGRXPm3V84zQxMwehnXrt3PbXqexoYjiCLQ0eCAwJ1F21BEdHmVNoYKXdhfB0Rcq8DCsReGYf4
7E2MjrP3jXLmSro3TSzst8mxyBe24iS+yS6uDJx8tkEfXWI3YJSPkedESkON8Mn8uhPzhnBrG3Ay
vOgUXvcqflTrduqWv8kEVnaqqFEewVjR2KZcJjg32ez2ewrlZM/e9KmhASQJ/ozD7I3xiBR4hEw7
HKKM5vXWB2fLYWpdn1chWY0BWvfYlTRzCOag+UhxzUFxXjXCYRAdDa6fS7NQ52dAIlG7tsSqdIjS
ezhxyQk/RnuGUWr4qsS465wuRW8Sc1eQ7675dffORYlyt6nA1YDOOzB60pTC6LxED4Ikt8d+1ndN
Ldjak+4OKY4vWEUfthaNdn8Wck3nd+gi10IlzryRloLf216limkZR/pb7Rjblwpl85PJs3vRxXvl
+r31FJBRUgWWnh9yAOztie7abTkuKrDIYKrYb9jPdUbs+JxuzqrJE+QL2WsgcLbDsIUiyOfgJlt9
jr0kJ1RsVg5DHBpqaDWf09DXlpGmG0lZzNFyexLO+oHvP7x4DCr9tCeoxIQpYejxQoBWP6djhNFy
CQOfQbogCtvyQHP35gMU/UisjFeGEc3Wdi0M7ikQbnll65yKHzjHfKFolzJ3iZh9JwWI7DMTdrgc
Ii2WHQbqa3jSoHt0ToyrXWuv6De+AzeE3Wc5xMK5gRmXUnUCQQx3FlbdY7/u6lLt7wybG7uH4BqD
zJmME18MxoM5CCh+9bVBi1ieCmMgPUSlZ0z4VxAzvUlbjt4oGu0cwWyBYZ+HmMDOvlX/s8UfP64r
0++kCWEr1Oe5WLlj+FbWuZZWNZOXHwmph0KdcyB5F34WvAjm4718Ks6R0EucJcm+zMPlUkugCYya
7HwQ5Yi/07PEkj2y/t/abZ4/d5wkXeY3PoyZR/3wfXA3tGgSAj4jPbkAo1MAK2T/SoY8Gtxjeo0o
ck1i5MnguYN4CIPDOrifuUC0ZOOqSvwtpFVxMwEww+b7JuEvMYID1PsU8+4ct77w1bMZAd2t10rR
1TUzDy/N/KJHkKbfyJQd242MpWNnMAbRdxQu082eFILrxpSEEVnksunfSHiGqAnWIdhBDGwHDqGm
SZhLq015v1dBbdF/PJOcynv/Jrv5xoKdXFUD+JoOB2hrXlBN9jcXLmRNMcbMtPquTNta+sXMZgXP
+LAAJQ5HJzGQS1PG8I/zPgru7UBb41mH7BNLIZ781mcJm9wqfZUWEgH0YxM6cp5mJI2YecKXLlxl
GmjgGW6Vh1bg5mWL/6VL2+822k1xNuiX23P+SQTxArGjjlbn1whb5zGES8pnCISd5tcgK7i1NOQs
eOWqgQG9H2V34kSC3WvFTuCzzuHghFo1v5tnbhMeDLz8OvzcuCs6pFlsa1hPWMv101jOZhkAx0yK
+QHoGIA3XJsdzJX9qGElyNWXfRHim/fiXGHVKGk/1pxDYmkU3PBETpdwbAVn+A5u8jga/mIE3f94
bjXNLBvrpjPT8fmOd3SkFasaHc4lIFAcGq+8oquAQubN5o4PgwstrJbZwXaZ3hLo27OSXYY4iGzt
M8B5Z+MxqkRa3FprQqf2jL/P1/OfWrvCh2I4ufY7Ps2uM+EFp0HT+BjNpsl+D5NXLoK4QnDLnzgC
u8UMLa5lmYSw4s8LZW/ehn98U3EGIb2w/DvkY1hpg4zJybXwQRu+b7XhwFe1WgDyRXFyZTz0561h
d+FN3t1ur2RuKpsQ9H7rT2F1Qdszof423QOLnj8N+oTbemkhtUYw9xBSWkEEg6CCl4+hNBZZ4dsl
QHply6lTTeDonR6TydGQWlkSXhvUwpNEcREqS3mYbwJrhjooCl0dAJFgb7Mce90ov7BC8PzFxY1U
jmiNZCalJOGC4ybHsQR9QtXQZPF9OEbqdeLE1QWMfRbYJlU6abUY6rFiRVrnAOxIWWrDM9Wbl3XV
py7enRmo16khysIR7htES3iCcusztMPlOVS6jA/aqPksWJa/JysK/cGHI7ruV/YOPjC7X8WD3I5d
HMIU03Bg4gxpV6y7ZU/1sl5AJ+wPJ3N2zCPKPZZKDzTGc2mMJhBkfGp6jg1RcATZr0Qvho3Z87hl
rDsyGENasYIHLsm7j9gfZCD2sIgYs77QMWB7ADbuEme87uLRVo8DkPSDnN9CHActnDAqcbGWFjk+
pMDpmL+u23J+gysGpvtFH5y62NRbYUV9kG/50pw/P2pDRyHeoNdEPtK7ldCNtxrxnNNSXuExAk8/
MVFqyikAKZId1iCmT0/imeXCEeTlylCU3iLd+BEEIw7cCFAVJFNiOKKO9/bn5NHxKsKsziYhpKSa
Vgh6Pnk+TvNRnfG7KaRFXpj3kx5WCujX2jBaDWwu3vt5/vojGJrHbFpT59bpnRGy9G/0uMFrwr4H
oa3gliNIQSgav+a+FtdL9l9YRPIoQHs9bSuqhhc8l0327Nc/oUDo4EKr58hNfpUaMFi1dHMzy6Vn
EYKlN/42YZ7WYMv4YcQHH2b3rCUgypU5fGq8ueg2NMEk8d6m5pOc3C3WO0KVrh3hQE0LKi/Dn7Az
MbQZHy87hPyU4wEnY3rAXP4fQm4KK3fHkvmF5+RWSWRoDgnuW3IhgPNVW6FNt5J5uUvjlY+Rx5I9
h1pNdfenqPtX4e294uTRKCukt8xyxH9ecNLyazsVEx06poIg2d0XkPQtE314MJFmK6uNF4Q5y8in
IZd1fk05mNEmezkYCJXTYbJl41CbOXr/M93Fmp6DeK83w6R+a7GpUX/p8jr3DzxPyy3vjxdTrnCi
XDi48eXqrDEhq3b4hcTIS93/Ls8HzQfDXRL9vw40wPK5AeLro9ivR/2fXBPqPw1C4qZMK+EOznN8
ZCJtnkEHGId0QD6bxzX1JXMkcQOLL/Jt7doSXJfLXtXjHeIZF1E47iQ/AK4qz0y2qnJH8T6zjemg
IAagg8ISHZUJn8ORetMSjwqg2ihB9z9J1bLg+DkLJ91xJnQAo66wNkWmIj6vumRxMeR5sVfPw+JG
Sk9opJDBOXr7Wb2dynZ0lI5OAyxv8l8k6KpBL/v8aVc3tdHKPWaHnI2QbHI/uK3DjqsgGcv2Kn2f
9hgk42mPkgv1y4b9FaK9KoWtrS3C7DQNAUD6VkJetZFIUo+wWCtbtayHGpUNW6euY8d5NvJga+Jl
PWdDuOw/KAVtrnTKq0YHzn7WUcPtmWY7C3mjsZOa2Zbb+6IGImyzoW4BfALnKbttLbFoN4C+oxup
rQaF1rXD9nM/umJoLQUgud4pZLo3tyH6s4A5xFQqGsDlBgBpbEZxFwjhOgC8FS0K8zQ6RYX4aqOC
8KgZnQwbT0MXfFy46hh+ahM73evIN/UwqjedulBdfzUVB+oZdClGaBxvqOLlZ15BDT67vLUUHmXA
ETQHvTFpFfxoy2PIGUL9nMN2snuc38d4ZTj3ai7oW9mGJLy36Uwdo2pauhUYQV6SwwKNgdf0YyI9
dNeyHq2M9qrDiZV2hFfRW09x4wrpxpIgtBZx/IJWQ4MVVQ8pNgPc+P7H/btVsGFmYVBOdrMjpAAd
UDtB2EAEmMWnTP8QepLCFRDgXemg2H+8EoPoIylYXtbDu6Sp63k6vatUdUPXd+iOKF4O6SwdMFSv
xlnGxhPu1wp87AV6cXTpv5keVxVuuKfq0AwrlIMaX8P2zm0PCJTtO9TfU4aS4x6d8L9rXlamoSVt
qyT2tXp11qf6FM/m43Rx8567OnodAFqrjbTWYPiDaUZdDjEdn+y2rKOjbA3o7DgSxyRw7knjIwix
ZI8ZMEkfkmbqCFj+txPST4dFHv49I3lVDp6chR6x2+x+2GXWXoBTvNewJwSnD6/Yt5vVHIftUsiE
IHQOlluq397CqlxVbBhCtnv8Qnp/J6yXVvKJVIfs5dc8U+rX7GfN7eemXqectSr7RZqL+rOVJBFX
AY5JklZurhToYG8URoElEnomSucOVO9+a/osVYs8OHUh2ent+O1c6aPaL3Uy1N4KuQhlUHYRxYW9
T+zoSdBO5EFotWphTU13QRQBHJ0Iv5JWNHimf6X6frAiU1Y5E5DLt1U9syyLUBF+bksEwdo4hayB
ibnYHbBvX6GyyRS6v5xNDJXAg8vU1PMJUKXuEK79x1zOsHB5WTQwpkXWo4/FNe+QyRrQwLs2KmWa
cKTYe8O7r1n7+vPU8POId+pBsPdrhawfBnTXvg+gjxc4r7c+g+afeYnzLMhZMDdtPen6AUHRCJUh
yUD04US4dLwoiZ13OEiNUKIFhynIC/Rr+qJcan2vJ2j6AfqwIcQJN6vcXqkitKjfcy6Wn4e2f4We
aTEwCaOPHI+H3RiFExVCdp2sSoTzryPIB91kl1k5rg+PsXkJPNqBsiZQF5ZMIAttwTkrQDaGqYeT
UM6yhqRRsjMvnZkVr1zTTCtFw7j9P6sZHMBocACB8Q/i+KcrnwUndx4FmT+o3Mpkn7s1oKoyyfhh
waHSHS299k+Y4OkiZ40TzzsRlu7YzuwtnTjuDh5FIRCF8J+U73n4fzUADBUZFWy8Ae8mMfJ2WJ0M
8z7g9u04CU8Ete5bswaTgP0ZDYFXVwsBX1fdiBXr7HXRTxWYvZtXx+AHnB+58l+3Bjs9kTdSj5RG
IHwxXQfQt66PYL+jIgVSDJB5LU/X6ksWYYsoLA2rpvfGmxtZfGOB9L31TpdXj/mvx9ZANQo3BCaE
Ithio/7xsui1p4hIKep/gnKpsYdsvkkwzFE8nlE4Wq2M53rvin9ZCF3Wb4k3pyi6IuSiFMURKtBb
xh36ZkehFV4tOvXjJc/w7toIrXDri8b0tgsjy0HFblhFpNqdz5jY4FaY+YTiKVCUrfF24i47FF/n
pce3/oHlqaJqUBa8SNY+2DdHa8P4WnKOaIfsZ6j/8cyiFbTE6ZhVXEOiy4MNdwdSbgjzlukoDOdq
sT5xw5FlyieiyxfV1rte6ypScWyAw0nPefmjdcZNw7F+0wBL7h8cyD/+l03Vbahg6oM50sdreKWo
4vYFPcTLMmpat7AXQ54LwjS8qOhIB75C5VV5rRD9/HyIapd4fvxuhBPV7BHRk7CcuqRKz/+eGUiq
7SwP/vKk/2bLIAIWqgBjUyBgZb/YkrYo0YtMLXgpVKIaiuBZq6sqAtZIMqnJO+am90AIBTGZ46cF
XOejagyVXAxSui4WxDuEHosHdwTirw7eAIbzU4V57SsyaFBsZ4nFv8wI7U278Y1IfZiAaWxJsVgk
vtDcIq50Uy5HPuO3ZjhasijGocxInTMRbORV3SpuYeuZYNFM6ybQq018Pr0LnVdRsoF/NoSQpxU0
1J2xI3gZWvHRu4EJtuWuBw4XvBrsdOUORP7a0ypTZAHduYoVpz7defTfsbVbTr1dmvIF07i4NYWA
LfgCw8XCTektyoz9uEvkfXbN2tqw4eRqdJX7tYJIt/1WL0g4KOp8b16h+Zmt0kzpmRwgKPGLo41M
jvG9ZeI/F5X/BDkkWB6q4dg/hJg+v6y+9qEqrMpXOh/Uo0WNEitb97s1iISe8/Dm7mDKtY4l4Xa0
QtUoXCpvVl43GxkMG6Ebusnn1OfUNZhDed5yOFGQqoSY26vix+pYVw6IxI1zl4qJ1lEQsK6hpo6Y
6OI/gTVhoXsAl+1kdD9GLhSCPs6nMLHlml8iCNby83mEi1IoC9+FOfbygwlpOqHWYjpeLbaG4PLC
w/DONLumHtL6B8gZpZ+ppYIU9Jtn0i/HkQ4qcJCKaLs82z74I4uuWaaTRPVvCvhRqAgWLt7I4qwR
EZEf8t5xsqtDxo6s7EXPLFOxf1QV+C6xcx4aoumcu2op+NhWBLp7Qf50Y9ZyJF1h/ZM3sx/XBjNV
2XRDHJPOwAQ/YAG5bf9G93q8rzwmhy7Mc+kX7jRrhV5e+7tIUPsLJtTaFriBBab+s+LS82EVk0y1
qlGuXXh7zTDgzgnEMw1V69xSV6H1lGqUsTXhHPcAsMNgLIrpXe/pZcs0aSxDoGQX2bPGAqoXdAFZ
bB8o3cMN0LDzdeG+PlHQkguhwkXQ5M8s1DH+wtJd7ojKIdKhFBuiR04Kn+1+gOcaw+496+izbC5y
hLjIF/fKv1MFAlb5QrgJd/1O+IYshMNsGph94z3zf6ZqHZ4CimwCMdjuFteIaVnM6HVYJ/jjC10u
7rDucDiqMastBn5ddq4PlVRX7BahzFFf9XlR2qJKvX7BaxRZUOxjn6URWN33KJhog0gs4+RUsZG1
hf+/h8RjYF5qUO9fZcLHCRiJAn/MYDP3WHjBoDew7Qo0xEeofzON9G7wgUaU9G5HHH7MlVcyg4hL
iAOgTPr64VqB9khVx8EmOk8qYX+59NpuD8+Ud2tfdqja4Qw8zotE1XICKHS/8mk5lKgUucKFFTYA
0JC198uJUJMgmkW8oH1L9vBBR6ZLh4u9Tg5ODZieDEx0b+dAu9eb7zttERCF3F0lm7AuZsdnxohC
qaUgfMJacdoSPz+TOpNjNSHspYRp5SumGpLSQcHbHblX/y3OsYt+Dt9fnsgIXgwf/mVBQ870J+6B
5b5JtHzDuDz0Ank9EzY5GZ+eIhKCjhwG9GyarEBnyuZKDUul+ocnV1auFP/qVSVF+rUQ2wpbbPNN
UlzF2nOkoHJRcpBwrAyIr6B4kZnvD1wZNDYaxWF/z8bgpIEZaqnudRgjYTziCo52dM/HXQjmHQC0
62X45SnImOiuHFHjaO23NbGZLQfMnwikX56OPzodFBzGndtRjHraOBp8Gt2cDFl1FEHOZNBGKohJ
7625Ni2gzqT9RwKpTTduWhOme4ZPlmI7tMbDS7K59eVElStI87N5VUcFW3ALZJaTiIhSf7wU3FG6
jZaWfvcP5ckmJihrLPhPfTNuZDNDqZ4iT+CBNMVziKGZEA2K11tl33WJ2z0aeXJgzRwkzNBC38JS
djzA9Bw8PuB34DmSWjtjLWTo/+aX9apbCOSXzazwlF+wpmWyqXdw8w+F8QJCEGKfJd3IunoZwcb4
ZIkHbQM9J1A1jbyf30NoRGOoJdTT6bEMwlVOW+brUYXfkll/SYUuUyhRwUAtg82cG+zAdjp9shtA
vPNR96i4OQvUVlPFNOEO9HmIc10PfUWKY64n69t5EZXr68Y1i5pSE/IZBhNVYVCLA8eJj0ozCu3l
AZUjkTB914qTGtkT3pM49WjQg0PkCaosskvXOOcY3SDO+PsDk+ztZnVqhA0591Z5+uk+n3rqgNCr
BR9PXQvQO8SwnrHpPrZa+AT+KrU40xeVk21ajfh/GvPL0nL1mZ1jqPKdg61P9b/LKPiMMaVP2AqJ
TKr3heCnsMQ3Y30jMgtU/Jy6elN1ZhQoY4EQgZWRedY0T5Y6E4NkVuWHB+x0sSCBIfrlKdBWeS6j
x6/4ugHrnTT3ULhhx234DEr/swyEOYPrf4LVwiTdXoK8ThQu2Fbwd6T6ijQxSnfULoTHrkeX+eoZ
bMpujmIzdrys8+GXYZWe0/zJa6cjsbz8MFLPgtwJUyuqARqf2n4T9CazEtRsRrwLKcoJCp+vTvQ5
xr0i65mAgQ/tufJz0NdtUmoMJOamRXP7X1wFLRfuTk7txrVlYFGnB+3NjW3oGz3NqywS5SPb+yJj
69Fov9RtvNWjoAX3t0HxTXPbi+EKPJqu+IRnVMzA+LxlGdjvTvcxiwWLSuddVSDWlWBbL5QKSUUA
XBZQit+KMBK0jalGVPCXhGCzrSIzZTzOCl7p6YBnUpqXXGJdYPPgYr0n4bLWRqaTmVHVssUrD1Vd
BWo3Jx6fHvSOO5+DwfufEy3rVFcXNpYg3Q51ZodNjc4k/oDt89krjorqYGAktx4PaCPb/4mSc6Yw
kbpgwHS5vWP0toUEoTIqndio4mcHIVtWKGz++gBcZSu6hDvzleSqb7kSn/BKQNLOUtWeywBtbgir
jC1N/sjBtI4TSK14ly45lhdokhAUQSJUPwqUAa1WM7+fbREHbEH2jcl27KZSUC8suaxjqpuDmkGU
id5sdh2sVB1YUrbAE0ZMpMfVqSfQuu64KCf/e4ANcP21OBoPzD9L9UBI/HgARp+GoX+RhWMdM0t6
R2Np6yIaIJJnjLpTuS4huj4DE9p3+KDQJoUY7DSaCgGQVJtpocBNrCimQhjQkdnXmRct3Q+KZ5+W
odfYsKNkh7zLCDgOz223Xzq9Ln+MHtq8pZ2ze4R0tuB/+isf59d/WYzILdZvegt4hQEr3Z90oR/8
1LqyQSwvGyYmiOUvPvAP9GKupV5uUg4tyh3g/ZKSsEHW6y3nHKWC95stMMB5SAjCHDwD1FrZuu61
vN9Vw6VZ0FyygohX7n7GB/q9yfItTPp6UTMHAO2WRWTyzG5MEZ7nxebbkQ4TkpCPpDEwlA8euRm+
w7PpnXYbn22zC7n/nsyNmbrmgynJ6wmHoT+FPKfot+GKt1gPRr4e49Yzay6w2SAVU/SQPNsZiZBr
+OW6lYYy4bfQpZr/CpZLzZwbSH7aSypiN/+kevwvZnjJq0eJw9eSsGZV6O814SSJHIjp+JO+tfjc
pcpYPkLubYhwVIf4gxJMKzPM/J0aIexaKQR5jtrnAUOCVwr/AHAO2pHNMvqPpaDBgGNQ/P1SU58S
4maJUi/srM2kGfH/dSH/kAyEVe5eLRpi1CrQwMYoL1EPpRHQOnA5f0fB3h6ynG2w/MbmGaiYM3Pv
u9FXaMAE01Xd2EkwFmsj8Ufq/AGiGsaLs0dXwckH/vsXnOZe9zU4oR5OCirXS/vub3TmdCJPNLC9
B0Qpeb/cgAz9zVdenHV1HS1aGnM8hcyC0ajOyVylaNKcgK4IUrxS69VQ7GfzqgPEuksO+W49X+dB
LsMllN8j0XUopUEopCE6Sq0WsTCXYULT6MeDNAHVEoMH517bjM/kJlZ1eCcUma0h6QZxlIk8DV6m
1LNSuWsU4DMHXDBO/1dkhHYDkf8vXCzrGfA3+bglFKP/Ll6RFpmtlJcG1x7rgIsSDBndVBcQQdhu
a+j6jPIHoab9O7nN+di2bfnpPFE9QLRC9g7kpYWfL3K2t5AOqDtIzYVQ/Y3Zih4mS9rjMbLaqZk0
x/MPyRYMD33+mQmcfmx0MnVPNnLwezgiRu5lUp+PAixf8LXcdaZyPHHZMnXu2kO8jPBJ3efdDTzr
L04sV9PQSird4cVMd7HOJ/+Y5VM7+o1dyU8nKGkZYRTV1QdiO7jdrDuLUSpUjkDN93ZrA9wuyV6r
zGAIfCkHbL+1tDTAMWFm86yifDWKz91aUlolpMnd1w0wHeYZWbBqcb/G7Z2ZuhbUQaOnkLJnf1Oz
dUQW2aIo5SvBHhMNeum5V+R5UKxTpPy0AA45krdNcFwdI7QtuVcpPioSJNGV4Viv4JS67HTDZB6U
pwGhSi0SqGh0yJfCAXzfrZxngtSyoezb67oLaYkI0LyLmP4N0cWK08FfVdZ8Ucb/JRuvgnoZuG53
DQjtkqHsuEFV9zhA50jJkz+ebXfpuPDthVkHmNsoJAus/BDaks3E9zTYjdVkmJRVM2QUn/cyvkdw
5WolRW2K7YDdlz86LJLlk8XKhG3MbdqHunJfwfgUIKGflU8lox6KnUar6iuCudmrKI1N/utn9zDA
vW3XVNzCvDaTCZg2f/uV8/zl7OKT9Ao15PJ5VECJ5q0wbxn5qc4yoaqNlwpC7n+HOpB7P620flrb
grT2fDQKYPVjaShZp3wGKzMB4oZa4+9AXZtNbE0xTYwLeEeFn9sMBXPYlZR3VKopMN7CnIDfm+XM
TqKVUpfXrg8Gt+KhzzlGa4Q2zF+z1TqxCRQSj+2sSwKm8MN9J2Ld6po9sHsgo1aN33UM9sirKWin
iCFjAcPs7yvQ+0LwYKOfrELTxx7SxhzyRg7KmB4pgIIQCew9QXp4JLf+blmVD9hIOLHYNSfoTUlj
Y78o5SetyLObg1qevUUiHTBnKWxdVsI/vEvisEPE6ITJdTbclu+9q+5yEkuiAwuqc4Qko8oP39gO
r8yQLbMFR3hpb5rGwxYKW2H9FZKFqh3d7uyPg4m70tVcPMEkcgZ6hGKFPsUW5AfnS7+Y/ffgE+7B
oEF58U8nTy1c/AEgOGZFRPBtbDycMA3Aphvn+bjMKNDRtLObzc3MUytq/QOgoBPPcWMIOURs3uB1
sK8Rxim/zCylFHCJOM1TE8x/MUEEb9JXdjIzR62ZhKUWGTjpVLHkEc4L1vQZd1btTxSzA5ua6LFo
ZbJf27qFGTZ8sv7mFdMLNK6TzWttytF8yoFF1IBSQCweH/ri1179X0bYoQXuwUJuQiLz6tWXDojL
cqnniyGPZxD2y/UUztVrwKuh061+kZQ3IMTFYrBMhl8tNd52ZWj4ZKOOsRLkcyTZuOJGv0SkvUio
Blwdxo8hpSHJ4V432aNRfvOtml7bSs+x0nLCsFFnBcG50Y7ERKYaqF/VGY0/sIyhHn54u8Y2Zy3r
RZzDI0QZUFuvwP8/mmlTD1FUiLDNVLiDZI1bn/1B76WiJoRwtL2K+m5ZzOT6Lb6fKY/J9ZVxG22e
JezVwNPYiyVL1s/oZYpzVdyjHAEG2RbD2xONHte1V7IOXklVgPhE/lBzFmtekwAifahl+XQa0irB
VAbRSW91JNx2myNgwnn6i9VG0Z4Vxzu9j5bISLEEeOrm87EyZn2Y71RA+cPJ/LJUqe7pIVU7Yy+0
O9lmxwqOSxnb7ME8IQfIT60UGa0NCASevEXOio7TC+t4ZZTotMZ2E8Ped6PUo//v7EV/d7xU+o7I
wlJOkjSV2pFbuM9q3PhH5vGhl4abxL82kI1eqzQWcFXJikAlX5xanj5A9Yyj3UOZElRjNMR0kDjd
DUFZuqng2F4C4gH+Dwe7ZlN9jW7tg/YTZQV7tBjogq3bN3+dZaSlt4oB1hVmzZ+fZDAl+8nmeFNS
o0HWGTsVbqOecchqJ4m6VYPkTklO3xLg+PB+Ke9o1nzvEf/WG01UGMfv4i+Ef5LeejSBkBOZsBHK
siLTyfpLxOQcyLqQXirNOHP5fpxAMvedWiumK9+Xtaw3RrTkhjC8nYyscY/+U2EhiGlP4zjmxo/s
/N8zDaKt6QCj2idPNozj+8Idiyw9IQOOzsxI/VJ5svMv0XakirkbL2m0J0yIyp3mBWYtbzG8pZxp
nNry/RhcaXnbqYkM9mXI46Tryad4jnCRuZa5Pu+46QcRzVdNPEYDN8O+X1CUWzg5DyDLiXixViJu
8R5oaECnOQaw7IcnGAhRtNih0Cyaiu0uJG4uDFFxlaJ3+cKLSf+pT2gLhePe+B6STxAh3wdJZqjo
ZikSQity3JiTDW+TfHbLJo7GSY5GqKK5urLL3l6LUaOwLVxU96TAgJrhQD/XZBLqIwFYh2VHKYFr
yx5S1PV+h4YYkE5wRC3J+lHeGtKB/4RTq5OVY9ZTItenSvRXCjkyfFhzF9yoJvTwEgQ24OhFtuc7
qPo6QARwZ5nP4nJeX6BPEx7uOT/rLa6CGTBl45zbgstQiTjwoVbKmIGKmPU3+RxxI2RuhAnZQD9H
/O/zICwD3DVa9poEWDlQTd8OTqKOaxwf/xgHT2yzcC5OxG1Uxevr22Q8Po92xKg8RI+LvZnTtq/i
S/o40f1qTyj/ACDYILQl8NRHXLH8JCXWHdiCgOt60aKYoXzUzd3qeoPTA/rjVe61wARWORWfGEgJ
sPrUOOpg0+PtkS68phx6kHyZkL3BfvOF6uApkB2Edga/D9vh8qfbk28Ih3znTRf8aROaPZf08+tH
9wB4m8wK8Ism8JbwIF9wRZMOkD2l0k4XeVxqgPPef7emqEjdx5/Jrqja3/fC2Qj6PFKBjrTmV4VA
lSAvmc2g2jB8zWgh/YmPftd5HYdq1Bqy0xvddVbDGYAhas86lQWOm6iBZSMg2rndZ9xGuna2H+GT
0Z9LhnbHKCCMU40j7qTQ0iAM07b01jMOgTqwN+Z326poNjfPXnLBJiEmS+kkbbpMyT8m8XA7kHvZ
gBPHKf4S9iaikxhuQ0Z1SL/uywcjwOaPQMDF4qhi3f36i12ZANd04dL6Ws3y2Ge8hDB9CeYcRinG
0BKMG8srfrMPt5Kthc3ez3GUqzYV9Mg6b0UXjzBJItMKNLCQzlMYc1QrqpnzNFqPbCy6erxY8zov
yXXEiyiRy2qjvUSVHYkR3JxHaTYZdejse1t8FX3yOfqKu7RFCQB0zFxqvDOn34ThpDf3w1/Qb2K4
NE5BGt51ujnPaBjnasWP05a2H+Eu+MbYkmkraWb9Sns0oGzhw4yt4yxpRrqgh5/qax2ikSbSGBG0
LZPHVKDKXW3LMq1vI4I1C4DgLQh0yfpjAViwhlwkvEx/QZlKnm367JpkcOGYYkfmqaH2+Y2F3ktZ
N0ztGaY+0WMisSrbq6cfQisFj3PeKUC+BHg7sJ8WbFtNW5FLvNZF689rUrdsS7CLBaaIu61vllde
Aaf5wh2sC6YoCDAbRHGEZaeAxpcqcuUf3dwjh5q8IvUgicN71qbigeNu4FA3ahOo0bo2Sy+MMKfs
suIZZOc+REGo/GqFtLKmbyFlIRS19qyvIQ9pWkt4zSastNBuARdMYvZgIbAdd8BKjWfqreX2QMf1
FyH9VQCmyIf68t/yB3QNBqeNPLW1lCxzC//pl0pS9kurr8OvTK0VLbz0eC9oZJIWeEPDtVXFmgJ/
Ms1ViuKV/MNxtZxPepUmFxj1sU7NcmU72daR4H/JgJv+rHIYwrOHw9sPaVo1NscH+h18AqAaJKh/
OEqHG9VDsgktKUrnEpZZ9WXXH5gh0FX+x0u7eAfSMnaIIDptNUP5KP1K5dWFLNW/FFt7fJ7BxsDp
wueiYAGd00j7Jtu3Zj2TQLp1gD/DWUHQJwW2cbdBzxiC1uY5BNEBiv+jNrhH1RAw6nCSfLBafQTY
8gUkOxRlCCzYH/ByKBleTvEaVN3CDHNQUmACPSgWaLu8gQxSogoKDiLRvzwN/YZN8+uCap0Hl/7r
nQJZMrLBvTIew0Kgu/EgDDe0FqSaA7uYB4ZSg680ylrH4tNb5iBMMXRYcO6zOFhthAwWFWG/jGna
MTh0W52Kr/yYsVLv0s8Lr3bNVUC2+L5LYWZ3Q04tSj3fRwUCfPHANWJkg/bjmBj+SeCKPhJ2do6d
USwnrEf6Bd40Y2LRLBigGwAlw8OIUwKfeOY0R32mcqaui4i2uZBmKr4Tamgt4GCiyRcB0ZAYE8Sh
0JSwym4oRIFhcuSstJoYxfnQhuhmHOFX8bkbaKuRJh4hJhPhedY3Yxu3l3/QiyJaUGF6jaQvERS1
Ct3RYjpgC2hzd9liWxO8XsUOZK+sMqNOwE46Oohf4jPD9hS3/zr/qyXVaNqrAg0/4aTAfgQvVMfW
jwLrm/WzYcJmT6YAjXUxZnBo3JXcP6P0gylvEsNtuA4WJMRYY0Ts59SNXqXhLjzABCOtByaC27Z4
atLV1qmOV2jt8He9Ggaz6+XivyVkl7KuIDOmaG/lz3uLXsd9JMw+xmCzIigzO8YAF/46wdTqilJs
c3zMeXgT1kGoHZKO1fakOz17qiXokulslxbYIWotIpO8Wad19zv36QMZu/C4T9F/mOTWNR6fuGK6
QCTpdPFHiOGgyaGkmKpCPNMiG2BNpqSZfjmpR9QMAfLgBES25KyyiLIeUvKe3F4huW6+qyGeHTE+
5l0PnaoSqZhDQpXlXqHEh0Y56HWbIEkbtVfEdfe456vGGKpxgvPWA/xdU/67GrHodG29U4EB8TlF
LG1LB9b/9gJcwZOKN+XdlKMID7hUa2QScgfTv7Kve/qFVvsHROnaGJZmtU5rjqXgg0Ae8vjhp0QB
9IyJAsQuBmYWneNNVyvfi6hzXTiY1e255z0Ioim4cUBqDjNqJeIztKfQeBDwrhzO7nI9HOMGTRRm
putRH1i2D93GYyi4zVJeTTyujN083V447QL6ELBybA84XTiCsOprABoaInelsLz/i2c8wHVQgutH
1rPFDAJ6dPzfqHGoPdu7mU82kBjV7ud9mIqgyTd5tz4NxrQrfX6rLn40yEpQQmdi+ERMTwsMiMvQ
DWhDnvLcbQK/7aoaPP5oe9MZR1kthCtThSmJyKLJfEtRFAShGQ7uKn80MjfbbcQYmNsUwMOaoQOy
fhHsfXRe6RHRx7YK21RQTS4+W8qzOcUmmEBPRadlcVZgiKkD9LSwsJggaNaapppbYn30exFBS9Xc
Xk8dLVbVkW39nN6Rs9x8lnjXJ21TtrwtE1EOwzkG1ZM4QKVX5oRjeKFQKY5WAPVpBcqGIC1LCgw+
xv8aiOhzbTh5xt0gCOvK0lSGc9mQf8slKcpS5c9pe12rgnClxGSjF9IQx51bLHeuKky7b/oIWBdC
Rw8/tEi2t9p0ZFFu9GAozVcInTKWd/UdpnuGSRBlor5vYO+WBQgDcyLZZWZBa2FGpSXQltteaGWF
yxuryZ6N+tgvKut4FPi5Dwr3MP4raHekBuhcJIXdDQK8wUa+fp4crGFcrRDktilu9VcVfbyVYPH/
6M5FyqZfky+Hy4IcSiKgtHojqp+wSG22qBDKQOpjok1LNXrLL7Ppd4bT+tuVi6WBM6iGiFromZHi
O67Bgi/rHsbOw9wcqvkhfdCHQudBcEdl1Ehcm78rAO21U8OzMq71Z7UDJ8HDEM+3gjwTekTIMhe4
jIN0VvaXz+Q6/IXjLktcjFLa5w3I999EOQ5cwwmeaAFS1C686fnswBQKaoz+zAKaC6yPYn1jOPIm
D/FYuvaheEh/l+Jc8VdjdJQgp99JSReXFefU3A/seU6vQjr12kNvxNapmLRotcYQv1eLuFN5P4Jc
YIITNmfylzaX6OvhajU0G2NeIOSHiwbcvJVvj9C5BiiXc7Cxq36JDMeat0xcgmvUA5DZwE1ms4TU
QL6gnAhl6Uf+Z47p2P1FpWx2F+XJjKYjNmeg4EBU2hEB+PtYpLKxi8vyzSJoQNPWmVvq+g2EP+b+
Bx0taaTuebl9PkE9bqs5zZ8iI4SnVxy6acg3pV/hDOMKB2cheLAEGN80Q3s4oTRYkF9ScPslecmO
Z89b4Osm65w2/lPncid+ChfuLkVODhxmgo9qP+Fu/AUfKRX9B2KpGIwR5lF3HDP5U7A9DrX8BjEZ
P5qjfOvwMcjBWGAz/6AKHR6lojaEwMx6p/mgQHnzSr6sOsgsZ+cOgDtpgxYqMl1wVcPYTpd+wEgI
W0YtJAtJ4owmVJJ3kz2VZHbE/4UQwwilln70xwlMhDd6bq019URPU54AZxjggWkPM3Y+YQoDNQ+y
WmjZTg4WLimyjUqsvGQl4KXo5u+Ge1PVzDQiEX/4b5NKSNLVKZxKqC8z+NxHI+DaLwkjXuzs4Xyb
xQMATfS8zN8Wh3Q+WgaS6R0l5GIIgifDobbHR15iMkP1Sfn3vxYrkwm2iCh0N/TCMjzqYitqx8gl
gHGj+rtJXmqdPWa3JqYPdtE2bywS5o0PekmGkdO1z7w3ut06RS9+pTI1cN+0j4nMNJTI6a6njz3a
XxyhsM4DKe+b67xf9hu4pH3+AbH8rCXP2mJt5ekqiVczYp5BCGMj9/w6u/jQNZE7eBtYstvofvPt
h5v4efROpy2D2+WNgBRu7gqvRSQPL0l3k+o4+PMiDCptSwM5yfVPhvijuEseQpfrUMMBTYhJTtoW
LSMOdeIE26VLx+p5M2W3iD1TjIQ3CQaNHqC2NJPVrVLUJ3+NNQaZfKCM6/0Q1wOWonsIYA2k0InM
jwKVUiQiAUodnNH3qp5rq4eJTY9ESnAaVOe6Q/m9LibXHfo5TGlOWgwONcXNq5DJrVC2uMdrdcxH
XiS5EXu1ZZPeO17s7Ns32Vh6n24yjKHXya1HDc5RHn7xg0j+ne8//RKtPP3qmNAyRzqrt7cDZPxY
hkNeFNBN0jihzbiqqwFNMRD/MoFuUnM+RkbCg70eRKJQ20ufobKpbg/2iRiDbIwUBR8Tsq2llIY7
Yc82VvZmev2WxXQR6IIsoYD5J6pqXXCsWTFGww2f+4aQS74U/GrVtMzjId1GW14nfIDy9fR51aSA
iAzjvGEAFvaEPdwcuDyO36G2k7zN8fvbtC+wOOeGinf5C34Mw5nhfqerl1OOi26P3X9E6lb9Nk2i
Kx12K16ghOKAIA2vQBbzX5dvK8Pf7QVknlcAQsgLAPb0x7tLVzjERY+/36yhrerq2azRZIQDgixe
mbdZ2uQxyWyWTSV7MOFZjWan8G39qF3FcVZQU7ACL3oEVFmkRyxtyfwOgetJI4YfmbEtO109FOwg
Y7iUc/RosfV0nlsbfgqvngNJhTYxfiXnsLLb1aC9Jre0U/ornyx7QI2epmyzxHrkaSfIJbkX+3iJ
c1pQEQnc53Rq6cX5HIh4Hzj+i7c4liSMFPPRXdRTyo9LWDapNQDXR+uHO0tvGUy2TvpVvDTEkBqY
6Tm4OoZ7Us9lfaYo5kmlYmciQu4FdXD2MIjQdbYB7FQOLGZOWuB55svLXtiV1F89Th/DK32hzAOA
5rqRD578M7N6/fss3whNVuMQOEWOB+md+WV9fGFRSWG0ug0YSpFbB9xwzybpdxlKYb8yvRxWb/0O
tMO8j8VtjccRaVtJ8SP0bLlnPa75K6LDmdaGtWH9syDeTE0ebBjAXy8JDy4WuRWYSrpkCof00/zV
OJZUbhMWTaeVkfuGw1eXRYap4HAAnaWIdTX30h2V9KQlffqXdZ0YmCTlYEUzh+WCJhB3IfEmwUYO
vRKCVaompr2583cPqD2oi1LHI9H16nsLKzkowj3WDtb3jflkn/16VOCOrDOH7dAUYNQmTSKGFLra
GWukojHOXRn8s9y6ItO3RQO52R2xnhcspDH4RS2Y/esZu+x8K8h1OgsTFOxDQQZiXr0jMBgkoyFX
OkRdMVYW9gSn5Er+56kQezKvxYUbQSxl6Hf9osZ2qgEAEca2rTqKNK7TzZQCacNcFFiQWqKUiZtI
kfl78y0QSjfbWczqwMs3JjppsDxvOL2+OS2jjPA5DNxDPl8EANbXR46ATCWSBZn2Ja8iTfGETSgc
/MezVfLnOcvv8NfTBE6XY5HCjA1369dblAVS7OxPypa1VNnr5Pt4yWnHEs+sXXUpjKCA8rOzTJ/l
bZF9maFQMkFEz1nkAUKFWo1rHwDEQn7vdlAhxQaUG7NeUh+uFWoIoPC0gophBYmVKpzd/o7wGpZW
qJtGXo+boR48/wiPN32tOMDAKFRHoIMvXEopA5GXXJamdLI6q3DrzAyw9riPYOCJsaNb5yhVoPJj
j4Slai//db6H6LDS1dorLceZvMOIFTO3tsiI85JutSOvJcRLW2OV3wzyVw39XHd7m9YLkgDYATRX
2qvtEE5NIDzxfriDJ/i6uJCqsZXMkWJ2A6dyTMhquR1Dzmwf8vCpmxyfBJUY8W0Mfgny890V6ylY
USByws0vfgPShrEqFsG7s3yEwgicTZXaTyNUCj6szAWOrUmLiYTZTEd2hhePOLea0t83DKmFiPih
AnM4n/VTSbXt6uAPdYNECdAxHjEZHu/h2GC3O/0w2JV0ofvccaa+uYkar5sv45SrDMOs2RMwsQLg
EiJgnGiczGHAxSG7jVj0gLa1A7okRjfQVy5wdF8THOvNJd2MXJwVs32KaL7TXEGGcMrQI1RoAYp9
NECTWVAIAG39oEFzG+tE2enUGNNzpTSVEFpZnxGA392Yhdo9RyIMnp8Q5veAkRUPOLirC0yZspe9
m4KRPkR/rfueTZ4XRVNWmRoprYOelkYsYoYtP9klyRQrui2Z/X1HPnuxF2KEdxEI3wbK/Ojx7XAG
9kdN5tKKzibSR3JPEpivnzUv6mKEkAd/MhyBgoRcJStM5eaAj+bQF446PH6wKeQd9uKBnRUSNCIf
RXxCJwmqE8VZ0BqWxKq/7HKfTHkAkesOr1Goyxf8RNoBaV6fhEZPGHqrH5M0s/nHZxK5oMMV0KwC
vSXr9Hej6TuQF7t3RGTL6GWjgeYq60fMfdoPYle3NMybgWl3LV402KyZDW2lXEcBnvGEGk+R9oQ0
/w3YlQsFUTW2yKuGzF1hSdA6hh0QWkdfj/DA/WQCrhS7Q0zXvsVY17mxktuT9CCdebauNLl/5/0u
NZCVN8vYjoEZCPhljp/XRHOflVsydctwW5dNH4ZYdTisBqW1FUjZXzRAM428cEH6+wM2SfeYUZZn
0sHgd+ujVKkXfSPAXInnEPSZo91+lLzo5H9Z1OvIuecPjIwx0Eod7WuZAk2cgEDZMBmX2PeFtNki
pB67hpHX+F26dJaGNpcatvMAbL9te35oYAPsElyVJdwqty+ZDDyVVNI3DjINfbFmQjuQUdpf/ab4
Ee/sqsvi2/fDzF+DfB91FOkc5/IRqzW8xSiPMluUPQ4vg6Xt9IdHOmIAqbZ+2fkYz9Hjar8QLKUR
OH+0OphwCp9fAPt79CqeG5naPKo0kdqnSDecOdpv/D/LaPmaj2w+01P7bZp6EngmD/wo5t8lPjid
dTMbRa652ddy3gsFhIxd/3pPS8PvUC3rzIcbRWS7zyqIKPeTxMqIamMpe1PYBRLQU6fHcXok8K+o
wLKJRFWVlqUJDGX0IKUkyHLAN5aXcFHAcp2Aehp7Gs4TB2u+GCLX7KQIZiYnx8QXoUVitI5cqEeT
Iqg8z7i/bXeSK59I+atA2yx2jnO97yXQixpcNoqloZjF8w7dqNnPxwpWYhFEASpviHHSnhUhKn4H
fvEWbIF/8T8V1y/HAzPAm4mu5i6NHqX9g+DSX9uR1KaIA4TnnGU+Ys5jBvFGuafBH4MPEH64xc/L
034sHDwy8ADeQCj8Ze08XJ+ygjxNGHguahdB0DUM/0Ns0/HZMbtOXENJI9SQHTqSbW0Yp2rLVEPw
XgvZguDpV72xiLLxFbrCKEcaWju3JN7JlW0fAe1m/1VfPD/TPP86XWg+hoKUYD/D4o4+A+VQaHNb
vzYH/u27wZoUbE52Av1KeQ+C8rluO3DLK9Fw8MrsH4bGV/5tER3nf+9m2N2Ob8QCWUCE4O8B0nbf
vPhCd5dveCfpnpcoH+0XvOF+lDLjTknU58K0RjEJD7L2XdrQ6dZ5VEMKgLsDazRESDf7h7PE6iMD
pohoMh2kymwTBlm/jeF5LL/cKI+oOBEpIrmqrdP+Lg4f10N10T80KNDg4vdeVtskjSsbmR2jGdQP
Na9uj+JdUglJyKjBzl4Z5ofAU7/iCgWGAwKsvuFk9tkLeXGHyrE1TTPYWHQGFuWDKFzkEK6MHd/j
BZLSTyrVa2WF1bcU+no++5rVy8V/dOxkZ/9xIfju2MjZVaDCI15R4eOgzKO74a5d9HpE5cn5OzWD
9C2nOFRApMSqOvmmHPA7jDCsssWraJEWhsYhGxGuYr8kS3tYwgGazc4b5VZrHQix3n1OH5G5wuid
Kp1PoW5y1aA+mKotbn+1Sl1aGzQlhO97zdx92Yiel1MFYfDOxrr0U5zQDa8S/tPQWEZkopeO4IhV
JKgfOE0S/YSkTT12dm4o14RPNq4xqL+YRjg1IoZeX94syNSjsdbovZj9g/iNMTBO6J6bkO8SSFF/
HvDABgrbkW2MoVfAv4VkavZQ9B7Fu8VHVBb/KLuF61X2Xtr7/2w3Z3vU8cvZhOvW9pPCBSlK1kMQ
PhfFYZo1fe+EXJvZm6ql/2bSg0qTk+bmlI6kXRxESNXEdIXr0k+ekEH+lbIAxHtS5FajwjsdWmB5
CFBN22dfjkxzQnNoV1fmu68jXHs110NGR4v0xey84xDS/tdBgKL1tg0NBZ/LW8bcycXNwumuScA1
8aM9YWzFS4wgysakc+JkEvvgV2DScN1ycHS9g3EKMlDJcDjDLT/DT2y30w8wuWTYipDxKyaYwklb
igMIMbmAL+VrZGbzJKLeFvOTGZ4Qzsbeycawr7lI3ZQYqHstUQFBvqfwZc2NEHzHw8X6+1wFAegN
Nj1iDwrAmtTWKvSbxk/V8VJ6aEHTHZlx7TW38r11JQ37EE0lVNIbaXy+DO8ohELq2Cno0afKsEUu
sWZC0AwKM57n5tnqUs+txZU1zGRfpl15ECgK9VzaMqcDCWNm/uynDIFwyGXQTEZKFM3c7NEMh+BW
Ylhn+RHI9qG6fwDKY7Dx+7asLiBiT6a0Y95L1sLb/ZDDpjFfHCpL/f57Q2J9DrsX2fEKt2P9r2Wt
dRC4u83IlIS4efa5yAUs0viY7QttAMgG8HK+GOgFY2DioZK4YOz6VxLh/iIE3FppAansppL1osZO
K6l1M03C4HOpbXhLXgepgT3UO8lSODBVMWPNWVDVYlUkN9Y/Ok53oqgLSsRS6yHTXVOE8rTctP//
W3K8Mc9TBF7z6rA1BCpOJeBEzF8z9n1J6NVQK/LdXEHYVcPCOXTYitkxnghyY8v1EUbOxnixlolW
Dq3TpDCg087MDcssZobQnFgIolG8OAbyzGKCm3TXNk8ma8srybdKf1bRKE+QPrzurIy7Gj0riwvx
FH/B/FEhRgnRO/NR9FTXplobodYxH038l+0l29uvGn+cb1uqar9dDc7WGffOWOBjYiaszogJS90E
98f4TgsDZL675hLW0MSNj/y2qieOXS8BCj6uZx9xrhYe/GonVwt2OCQeCb0xadWoqmtD/EowxRwE
M9ODHqU8WKHZ4LsIZcjo0PmAMtsz1dwIDxfwMrAMBUyWRTDTQZAjdN/F8uKU5HPqWQd/rKSGyE5q
SjbHDLrY8gnbmKmjK4OCRPieR2Jiqo17l1Vje1KgO7mXw+nqoSeCG7MSAxy+U3DOGHu/Bifx1r7X
BdSX5UEVo9quVa+ZITgqqxwUyZkLwLwaBldipWQSUl/xNhLxc/tv9rPhf1DZwq5eePtXZyu8i1Cf
KJ8N5bi9QdEspyKmL/iJ8kZIGIGUrzHBwq5svUJ1adh1gKE/aqK/KcVGCIdO3ShO418kH2L583ii
YQStu+2GZMJCJhhW22KIjwI9FD5jstOerO/BR2mkvFTWeYNcLyoYtqajuRn2pcgggJ9RTZlrGS6P
VI7GplFXeTmVruw23EVoSbf3bUxTEFhFpwBrBdQooS2nDzpq0lI9KJaPzXnf682ZWWIJuU1CRac9
eD4q7hmaZrUWjDeLD/ZXFTw5WJ7OLtYcv79sqDaykUQAerBo2jNEM8uPiOGucd02yrJb5XDFfsas
0r88+a12Jg9XEUO+GGmSs0+PM4RZ64eUM+NwgNqvr5sLR5dbSiNIuimT54OkwAiiShggvxifEyvt
zhNIAIrjGeFfMs1sKlhe6EgjB1G5jon06dKF2onSUg/3AXD0ZIJldkX+fje/qmGoH1qeNvtM9qUp
8ejMO44icIHXNGSn1XfleCEd7rjUytRcqYJCbhn/XR3UsAwQMsLBD9Vkk9U5Cz2naRnEzTWyjDTi
R31xG6HF2EbLm8tbtriAEnKzSTvApg52qsH4RTL6u9NU+TIsF8O04nUnHzC/URHtD9nSx7BG5l2f
U2NZVfhMFkDASXMxZdALfxUcG3mBWnPQfjWHeEg7gtmx8MUYYw5Ei7X0/9+PESoN2J4bZVWA8+yp
+fHgCg0lze4X7CKW25zNuBJfZ8Sxch7y+RZwaoXENFD+XINAvelqdOUlpnZMW7s81eYamCc1nDNQ
USzi1ooONg2P9s2zd/ttfryt+d1GcOHoBH7S5v8wsXBimd+ZKFrsiItTMKYRFKJUE6J9RVvs2zSo
3Rs8ADTzjCMUFtSEnLztfkUAHd6FLqVoKo5dTOfEgqaZUGGnbs62oVoS7+hMe3mLuil7F4DmGvEu
jSuQ5d0ONUq2Yi+BOVD5STZwRDVeUyaojVAP75f2RsptjMpcIex1tzE+0sYcgXMOeE5vUFx8zMU5
nvebPADp8BrHJqJHxgK2k21gLulG21v/lMSOxFu2BGwYxyMD+1FqTZRrQRPnOh62mOdn/+IZtoaT
rc7dksvNxZ/SEsGxIFGQwwACYtP5Dnf+YH3QMiXrNLKnYGL/e3sBLJMSliu7wOLLtLoTFZeZph1w
MsZPkjHbR5k7e/pzxFb7PSlOiuZCTvB9i87Wo/tZUJuvqFc5jYUl81dBazWypzhFti18YNke5kmy
HC2H7lJ8boszk6VHhq0b/RfW9PUH0xASPdEuCK6ahE3FbVASCHsKxWxTfvIHNR2oGTGa7R7nMTGz
8+JpkeO51u5NpogxIK5tCN+/ZOdQaFxFTgoyT93miim/4aG5MSpB9Lmh74ONiSM8iyiMffHsEgwY
8A6lRF1SJzQZ6kpKySsuGLNMpdPii00/SWsqSnWCk1XLYmPyuUHKZmjUhOfc9K0LVALo/cG9Vz87
V8SBXnpmGPZBnjrIG8k8XhifLle/gpJLPmRXfFaK4JaNOwvlfSivFVlO3ggZ+bJG96QwuwvM10wu
QWrr+q1EoumJcB+jhGDGiMRV8hbKJlMk0avRFJNTJmsI8oqpjJzHRk8fvUScpx3mqz5mQ4IH/j34
H8Xf4wGeZDJIl5R9MjPWTHZLF/06qFTvjflVyxy3yzANNZOZTJbu36o+M8ltZMaS3bYNXTGpov/Q
jJTRJec3Yjv4xDkaj+aqx63i4opT6Z5skGFZvsRG+FjoTPNnNCPVBDLQzVf1AG6jNPpIbBGeX0Ta
jbtWiDjD9VfoK8SaNCz7lNtXTU+v5afft5jYeGqSc7wg09dFC18i1VovveG7vd9AmFO6p2eoyrLb
W9WaUSG2WV4wWSLwFuOz2I9gm+ddWZ1SoG9s+udqEwMDizVbNDAqUNn69JFtnZTFl/w8P6eAhK+A
H38HFtY7CfByMwff4gTBZASxgdAcT96gXvFdNNhfGc//a695EeVgbolrCgFT/R0WhGX8EMUfbhSU
rXZQZJuogK+TGEMSYtPmRwyXqmPQbilI59AoExbE3YejZkZW+V4MucHyGwSV1s6I00E5tmbaxhL4
Sots4zXP7c6vEv04E/83VpodzIwio65MB/Mp8CQMfb/NyVaBgI4q2YDywGGOs0sCJa9NkIKXd497
HqeYfgEq9dcorsjuX5q8OuAZcdLTGr284Y0Nhl3FkEGeOOthtiXpkCSjPoxzgm12JpDS0SnAUU7g
59BJsm9AlkZhWMK3a54n6M4pkziXzaX4k0Kxuy8RGtBC19VNqb0JOfjqK71MLPQ3SktrDr3qP6FP
ypg0TSZKmjuLt3U3+Q2aCZ02LVsgrroeOeWIZlHGtxwc+1WYnME9wcrETryJ708HYDvF4vvNb7Rg
vaUEdrCergped4K+vuHxjG7E7x6WT6eqpp1ck99jeX4v6lfGQ849e+U6HR7fRBXpNel7VdcHbmZb
rjZs+EUY5t3oTA+V2q1a2L0JaD2kX6B6sgTCS1kiSWCBvaCtIkK6LBTC+eXzBN/KUjwBJ2L1msRh
1rhhkW6pQI2jP5rwxvO/rahXcECpsCbq/M3qmJM5rpqKt/GKPMF3zR8JfMHbqZlcYryKLpRe9QP9
b+PUKEnvSD2+qFznSMNG6+dgah1I2fdAfgqTpXX7b9bf46LZavzu+Lfdh1z291GVP2lGv1XO+jDW
D8kK7wcN+E+H5uNUsOf7ZEgoxIXKcHjz0c2WV/BugoqBmtoGn3+hkNPJ73LfCfKVhWufm7aaBroh
1LaNMgb7QD94cllNj7EOVLRiD3WtJOT7uCtrs+6B466B2hdze7M0w80h9zmXjbTxCBt8wR1NLWI0
IuUPekl8BaH9RE9xdXsUthPwNcJ87YgWBpzaoBz+gmeAoMHr9TeXw9qaG3sJZIvShMLqji1xPL2y
mg6ItI7zfo4gHpJNx4hN2iQoUOL7gNkZTv4lHRsAVKNzJmttl1sKv2hjbUWihgEeBtMcUEjxnFzW
vH0Hbyg9XITqC5JLSN1HkFIumTCxxgtSxflgF165kQ4PacqIWHARC+S4Yx1OpLvj1i/VupcTNjS2
ATfhx5AeZgmkCi4w06iHQC7c9EZvsk3d0lt5DcUMSii4X2YvJj6YkPYYrn8cI+Hzv6yvGAtID3Qz
07Ii4pOmbVNjeSD51EnuoiEQsYnLZsGgG0hjdCj1tSdyFgoLUfDPHi+31+GPFjmZKMzUItJ1WVTO
+eWpZWvYO4BnpzfyWUNDYf8oZDhCWIp/pPWxB0Eb/TeFMiJDAveqWOzzzJ7x0Z4RXrlwOTBmaTud
Mpg2RrH9ah+PAFZU1+sjpN58xgx6Oq2YST5a5fBFD/VfKFuQAp2xxJ4T4hQ1FgXtEr/Uz6XFsgjp
ZPnySzGe/+wwKMznzyl/sTkBMRcxFFXatqzfIOIFbpg3Gifqv91uFM0/KP4ziAvWrUyFM8UugzDE
4yJYjIog9TsdtuWfMshTB6csT+1qdtRrgXJE9Pt60OeB1kFCcTZANenKcfKRiY+kopohNaNk3aVp
d0M+qAeXPuB1maSfBhBUpHq1h/1fgiBvVdz29FprxmPHEtzdcO2/cuT15qzYlRdCZI4YWfYr+DMF
nUaQQkvtOCk/wQItYoifgoVhH0eEyk9EkkqmzwAsV8fz/kuvjPcpfQDAZY7KA2O3x0KZNSCKO7SP
7mMxLrUUZgOP/0NBlittJveZb1132F5MgQpg0okM2AOcMwev4NW6SESo30sS38gKvx9MafBJmiBU
tK6JN+loOVmGWUJJsexmZU4JvUHGwzKmJxEG60ywkFjFkE+uSzAAf+GBu5scf66DPMUyUDlhwSA5
5GjPtTSlDIzhNin+xBbSnXSojSBao2EoGCth6/m0vgsQvpx28+su0k3xv90A71v89miK5CrPXLwU
MnLw/TAs9LIVmHfFsOXW8ZR/3vZKKL9nulBWv4MaJ7PdCvZ1H//wg82mbApB52hI0nK5UlGK4ERT
eOwwByDk8KZjL8DEF214R4S/OMNAoCw39rSTYOIyigAdTwDmTiKDW3cmcJ3vq0YM1jhGUBQn7fT+
2yzpKyWMejcOJRlF/x9QPtFYKx1zPUms83EG/T/QmaMQph4r6NZGH7Wjx1VJ8g9it6AVueXf/3U6
FpQpSbg8uWgUC3XB3zqBQzT3/hECUXyljIS1nx85AhTGjb5jSk+R9EaUZhjuvzc7cLwu76+M44Wc
GAJaWgu5TaHDT52VRFZjlJIV/BfFunyTEb/S2ixlOu8Aq9W66m0NonDX/SxRrolaQKEJE2mK+Wk/
Y8FA9ITJwENfmiA/ZUJUTURHoK0JUNBX5Clr/RSO4Towjoh2WjlVHo8tS1kRLs23IUb7pt7bqwUK
mGlQPVculVh1HCi/1HK0Ec+tXgEyo5YMjDh5z28VaIpsXMoaH5BLbkfVNUqrJJJ+5BFYelnc6uSt
TpE4aITlG6qdXa71PSXtX1tfGT0bGNQMeC7O+p6hVa+PqXCQXUSC5TUlOuRNeWf82TG9iHRojqJo
C91jW6pwRU56nB4w+Q8gVzpVjlETC3JJR3vy5ZFpIWtXuUbi95sCFRDIfyNxXTarY63HZyZVD57x
iMf6XSNgK144pjHQWIidHkUOZEtW6ejYjtndxVqlKyAL5qPNRaeHcUkDDk+S2hCDKSmi1EeJMDRy
O++0MRjjNU4Nfy8MhSIPZGOdDY1wq27wkzXJ9znZabBpVNAEa678c69PS/06MWbqLaHSfMj+UeT4
eG0FW3JTwluD8RgAMzj1Mtir7eCKirk9+tMX5IiAE34hfws6FZTovv+xgVDOIO7aPc6qlRCF7pP/
60sAlrILhjGJMm21hbvzQesBfu2b1btckvuovt9mnB2YxvavBN2gZ8Skt4l0cJ+QYCJuHZunWdl7
R5NrpS0PDxluvWw149jxsXOFNRNRI2wDQklYC7Qz94WZPU73FpKiVA41xufF6vlya2csUCFVeU25
CKZgwZ5KD0af8Gt32/B1NunLHJFe2NNyDfcsgrfL0rAMYM2TMuYyJbAsoCOeN6e/QxAR2t81D+mu
+/gqhmZG+E4MR2ytcQxxFgKz1H2LdGsiKb8L1ULlJMbXxsJEGypy8iztyeT0FjCggAsExdaMWhP2
qa3riqzothfUOytoWe0LwvTOpI6ctnnyYa1ne7ZFhkYrVnYqkE7nUDI9NXJULj9raKBpIRFIFO4u
V8BTxNRHyM+borGXVKEM+/otd7KDelJ05iXHSNOR8ySJL/PWHtvu4cTeB8MXBIpeNIZQdjU1/eN/
pp3GA0vh8tnZt7hVyaQhamQbFVQpbW+lYFE1RoyLDYqKoJjF2il05TxiXuMGR5mDtN9qkrxVAIdS
xWjT3PZx3PCXRXcS+uSLhg08BGiexx66FpEOpqD/16QY1NkI57ECgWVZOUFe5r8V751C5/BIPrTo
q3HAv/3afiR9vJMhzr6myayBTVfT8/9YpBr1G2IN7ANONIG5CURo2oqGqt09ahlw0IWDTRjALBMK
JO2nYmSyO4LRBzj+6t7b177FAr3f1um1qVNyMBRij94LNinf724Fa6hYnVj/FSFJnDuXdbQaSvG0
EutjHHUwbOIbkWCgk7HlNn1TH7Lk3scTGTcdXdLd7nzJrQ3fqIlbplJyNi3P8BvXFWqg5vUKoG4r
hh0++g5cGwzGxbyg+KuFyrLcsKsX7taPn3xaxnYd8Uzp8aYxHce2L25qUfQGVY74MLF9W/rgcL1o
R0fC+0ZAt5Mtvt/y7m1X29+zZBOeRFfvTTw5Dd+JFAooxVx03q1p2ubmOddIoRoTnQIqpvpPCLti
PD8aV/EOTtifihr55jRPjzZabmoFIIjtusDqhnYF4bv9uIz2hMwDfw5Nkkmb9mIVeAZmKkMWtjZ5
2ldcWSOfJ0C0cbbPMH9UnnrKK4iWdPSU0Y7z3ceQ4ACSmb8CvTFLg6OAjCru5IYMJ+Xd/zuBbYXz
mAWCVPr1hCAtcwCgAPQPP2P5fiB2aQTo7k4Pp/nCqPPDtgrggTCOVu/069ew1E+rsnqDcqiehFgg
2x+B2PFNTbJHj/05y9OnaOYF4cYv6MAl8QO37m4FUAGQEqHv4Rs+Sj29Gyz4HpD8XrbKpWb02APh
UthS1Ily/SBY0rDbRENyriFOifuvqqaONiGG6/+AWlTRYhWyiTD2KOLU5DwCkqZ9joxje8bdulpE
InmQ8+e/bhxKTKK4gkXl9o1HJboDG54cB8UvSp9FL0Ai6QIw2CYBJDKpPHlskVP9pU60suvl/AaQ
tZ95tGFsbjuIP9N4JXpjsfwfLRY6H0WmLmqMvxIfYMt7G1ALjT1OEPppcHfUvr2xRt1hjO0KgXlw
m1C1vhZKF1XqaHYSuy6VRvOekoS9jOBENAIkYc47tnomdXVBKdL6fa6KEtwkN2KXYRDc2wIUX+Vk
gxuU0RWz7zxH7vyDLjKnfPP0ska5tsTkM+ssgPojRh0yjy8ntEGtYsWYgGDjoOENRf7JmPjvnsL3
eWBcZgRI2PFlzQ1qTf9wCfPtHv6a6b9ymlYtt1rnNaoXq/Bihes+6bab7hV+xONDRlpD8qM0LMpD
nds1YjlrnRJvEXT/y22gP7ocX3fKxJEtkdFuXFT5UEppLqeUm+oqOrDBcD2TbXakZAaM+cOFQKY0
ywQah7uYBUDmnMeiPPpX+NeKraukCxjmBvDvRlxcM1RqgtvBsmD4wmLonzKTzknY9tuZNU43VY9C
WePjrCaQPB8t72yUDCGc1tKyZQBtZLeICfcnrYAlhdYjx0OR8YrJzPFadGGE+uDEtHXF5PaPqIMV
FtJeZ6J2uo0DNcrEyIaJ6/q2ZDoY5f7zZtSexmGE99n/vQZIjbw1gZY2EIRVllMizTGDbxsMUyov
hE2zWlwRtn0yVJ4ZPeTk0gIKlM8axLQfgpYwvHraIocmyn8XdsT49ia86skKGdVBraPHSu0Glpfa
HPX7/arh7dTffEnCX6bLdJ/Swg4oHjWKTCqjpgl6XbduRqH/b7zelnjGfW35MTIbFK62gBFP+K4x
zLHqcYRKl2KIp+J3O4p7dnOFaUjMOUl2qHdxr43liUmcU/Noc9f3ed5BS1epFxlWAzy+3CDL4BRm
/KnUW3MilPa8O2ZU6lqETH40kyIXrDWQO7a1W6fN7h2Ddl8O7A33NwdGLB8juNlidNAqTa6akf7B
zs55ysEIA+zF2h2jzvn2+RFmyIzfVZo9dX5OeOp3dj5IAbHAqM8wtn2Ry7LiXtmdEzFAcCRVWSiR
eJqwwCv/d3qut5zR/0E5VBQUECwa66FodOSJ6wR5GsgWgoy7NkB2c3yUU9XQ4q2HhZViU7PnOGZu
TZDN/LGJBn/MmzfW2q4QysCEMmi6oVZ1Iz7OoXXLdfYH5fi69sbG3URjhgOQucr2oY2Znp9Aoe19
7buU5wASdhffd6DfJwO1exZZ29f9lhZjfGHJ44tZfM/lGAmZdukkuSEX+WN09Jp9rhJXgEsME3CB
IlqKkq2wBx023SLxykaB/2Ns3EY2aSb5/IOLlqzNUzQfaYFQBrF/X9yldasOszlJe60Vh+BrnXZo
d66a1lf96rXkJzOLWnLnrK/zqaSjZqusHi98/184HRHH+u67RkseTYqI0kSw1NXx5qJfWBoG+k8I
mgthkvwvjFks6VbKedSNMLBUKEW7OqiN9rf3eOpff7zXYmkgtGV5TNINoIcCZNu6sqsYl76epRTK
Kb+vQ6H6VxcxB1izujYALiVHley98N3mHd7/UT8qG5askgsZWre530ZlCeUebLlU9SrpFhR2pETi
euW2a7FVED0/AzWBQgwKy0G5/tFABDh+bKSAeWGx3pOxIWpBX/vjcrxCdSRgZ7aHcrObwaPMDhu3
wpxQVhW80xQX7tGSW70hnUtTsUKrNtN9gDVdtgfsPa0fqPACgcAzxZQfFJvw3KGQzJJbSCThnxcg
Ad4fvt+stSh3yMwNIPdnJwyUjbKDQ68k7bBkoA7+SNKioaT/Oqc6GSjptMA3SfAuEADQjZ3xKrrY
wSj8BYUWfVc27LEGHY2vUfuFmKZBmvJ6bdvdhZVeqeBNVJLXbx5hGBVIQ+snaguKk7I/9/oMcxyz
WnaplAbMtckhGTgyjfNlreTrB7Cxa1bVUlaxn5XTnZwjR7Fip/+128DRZjnfeG5kx3bKccr0kjH0
s4DaCRReuyc6kLUaZu1zWbXuYwzfu3H9ZsT2ikMY/dubP6HNqwcIDdy9WswaxQS8hYEp1/AbLXYH
BeMq0erJGYBZHjG6i05JgZUsKxNrDJ9uuMDxD59WuMkAfTvFJv4qKP3VWZ6u/v/HUUbDVdG1sQP6
zxU3U7z3UREqJ/NM7pjgYnqMKdZXFX1YQYOH1MVYPpczghP03fgNyC2PILQJsI/XHonVT0zfoeA7
+qOyuo9DuE6yenCljxOvWpxwwnpLEap6P0fvOH84uUioqQnD55+zGX67gKoN3uc4wJMwDzOyKlB7
WMY+/U1nwD/9jP3kgFOiMoceZEsRUPEHEk4Ff61mdQinKNmLXyVmrnvGx69/4YSB2IdKKdBCqZFD
Im/nYgP+54fUQ1Bzo2BomW16uSDGRxhQw12Lk5M2EvVdMQLFJg/Hui/TjoM9rRKmALnKOO3kRyQt
SdJTCyMygTFXjSn6dR+T9ezwEOO/J5byssWZjUDFD8GJV5RnTAPy6cyBYGzTLw7emIdRUUXGUQbN
3LK6ivyRRkamZm65oiIUfqA3r0lNIzb4mIA1jXs/FTTaSjDjrqz59vzbkYB2ln7wdMGmLXb+JtdD
zgAQuFGNT72lEnILJhH4n211Ot7jUHstiA0Sc+0F5xwHiUdKJYuwnxh9UtrPeDpQntpkXeqkvqYE
nXpNtD87F28uY/oSlBi4UdgOOtZNc+IBFlnztQsSHEvIoRE7NT6HmYp/nTI74oZOC+u87VagVTkR
/kgd3x+E5+58VpKLCxW8wqV0FFqmHsCneoQ2HMRiLfbV0RfclXAW+5syWNFftQchazx9tWlpBpNW
mrvQS7aXqWRUQr+iH8PpWTSkNg6hCYsdWdM8QBGuO3YKn8gSR3W9kAuV2ACu3qyJ6FbAUFOWXztq
onX+VXgh9wig0J6JcQba0fpIR81Jxo8ePWp3CwfQi7F2G5UFN9l63AhahA8U+Hc6FPs6xqlNlguX
/UEeU4kDOE97oF1ZVIzFgVupEBo7WCq8HGkslfoPfDxuO0i+SDTbbINz7wXXRLMhRVfC0oI6I5Je
1Necm/RvxibFu3t99kSBFbPdUBmVl77NVBaq7VfdZKknZ4xa7VSKDYz2kgqHfVexcRM6lnyu1tbT
EZm+nQEPs0rO5irfX21qZeq1kNf4lT0VH6lj40LHgaXLsQEVOP9P5BkbqdGcsJ6mgQkgecX8T1VJ
r9cW4QMIX5vHTNVbfAckg8i57H4HBlt+iqKLkCUJx4s4wG9qo77FyxKb5iO+xbDOmRfO8tSatvX6
Z9i9+KTqLhmgNyBUnAnlTNM2zM4+7QczYw32d8cgmJH/F2meXYZ/UtzTFgqcKLsJgdB8K+XWA0bO
fukTF3njgtWq38TX0bhKPhP/71ErPF9o0zp/vSeUwFPbl4VWaJbWSvZ3NErKuF13mFw0k+/KkXks
Vz1EcV3R0IJ4rOg5KZRH25ec7mqrsbcOzctSElOixfQbatHRWKsC6DaTvkvWFXqD7titGPMlPwz1
4yRkORZkrTi850COT+zeBDxSRtoUYIQtCfdf8drHXVmvS1oHi2AaHb7mn8hDuQldxo/Zqsp+cviU
1IHAX/vma3nYB6D/LpgJDqRfQr5cNHiaFu6Vil0wMX1kpz7+W35MmTAPfmuKG3ihdz1vN5iOrkFy
IC9OaCFFRWHn9ibA4vYykDivI9yi5Rtqh4T5gHI1+ykZhdhALPKJ1GvWJaT/QneMOeJg6PLawJ1g
0CegPIIzFt54S4cZ78Uz5xyaXRUwWCifMsU/5fqGcHDs36RNrDj1K12Bb8LBdFpwqI3nLqW6wNsy
GccpzatdqsXbV0+F+qyGilUJJ480dxCIExQh0KKy4EddC0++LmzzODmvETlPsxup+fFBMCcxdJ+p
YsqSQu4Ms8cave/UgxoTa6na65JadlUA8pAvSO88KkGosC9YVsLZJ3ogWac5R16yq3KjdEC5jthb
p/neGD9eYmMk/37in7IjWqEzytkBoxxvqOUV0ZIdtX8L2jLfS+PWE4MmGFSa305zzejv+Pox2GJN
kS2jpixWbLDSFphqw9Bpa8XxSZ7c2oxLeN7K+gzxFTyOYXwuydU2vyTxU3eCLQ6OWmyjr8DRhJmz
icRzwZd5JpRArtgxZQVC6iY0Aw4maNoQ/8SNWZu37KhC75SYeWRMbYjGtLgBMQbN/RmYn/3ZPHhD
tB3K3x8ZEAbG3BCNSqnYi3YM6zMWmIPQvRYzWgRpyJ+LX8SIafNKq1XJBicyBCuGfOGrBcUX60Px
BcNGpq9WvOWqf6o5AxIVZnVqd3nIgd+rd2/5HGE8Xm8yBw+sknnvpcElye53/eMAIs3pN/Qc6uG7
Io+Ott7863j4FGFgI41ANkNgllzsvlrao1BgsDW1G5KZYkTA0zof5LXLl4V19+4deo9+lFEv9+1q
W54OuChX5LlOmpqLGxpm7xRn9UNmerT4EBsV4ajtpEfw6uXqz+kvhhOo/9EHzkZsuJ6IHpGwrDM4
2kOt354W9p52PMzZghXqCInakduAM4f2tPviJRW0LjhWu2U7e5ckHtDvJy6YyrxpmN6nG0OXNzoS
XJH6bjsmKJwutNmfndWyrXmK3iQl1FG/DrfVfnxidwohkGDYfhEFy3wawy2npNmIc2L+csZbui6W
QfT7bpYsGpJ7sxWXbf2We+EYHTowOovJtJBHpEWhxX3XE9ApAdV1IrtA6jC2AEr5zfEyxFnWmxbm
puv4OhTyt1o2rcW0riq/fiSLMLRqf9w4+XZj9z5SeLu9X5r0kLzuaVyZuL0OJSCyytP1Vlq6vUd0
EQPy7Cq+YLv6AJzHmtsvbPRmHqgDlpJx8oMQ8RiFc0nutZFj4sapvF8h5to93U9Q9lH5RrkfetMf
5iKUDw0BkNGWarapUGPcDu9non0lIHYwcPM66BoswQ34d4L3aQEaFah7VuacOeum6wAxdeXcC45j
4Z3ekCIg6/bct834pVCshMGu62ubaLdN2abuwIG9azFZKayaXqB91Wv4z5zzOoWlmhZohS7NTmUP
7yfOTAU6GglvfD6gCGTd03aX2MqWrjunfNjyaFI8ghMEjEJyLVqhhmG/+HBmsw/qGio2cSys0TDW
RjNGEZ5t+EhA//4RRFGfxbEAeNJ5RdZj2rSEYZcb6yWHSkjalPXYew2raTWkvEQeJI3z9m8qzh6T
PK2llDKa5ZU+3GcNWtCfdONqcsgxKtykiAIhtRP4rNqkKMDNns6lBhwbUKaR39QmuQgXBtrbs/NL
G5x9Te2XjoD+dIVRrzKtmGMaKCmDRjp/BfHUX7RB134aX2KRe9F19uaMlXXkEjEXT/rLend4MyUE
0YLAah3L1eUolrfLp4CQAfApPlqW++Pt4aWEwoe7a31y4YuZZIN4ylQ+688tBoZZyyh76XGX9san
TK49vrUT6tCkG5n/SPA6WOoR2MCWNIBV9c3CsLM8KzJdqsq8tyostj9KndbNA6pofNpdBIApSxk1
z50OPpO1wMf1dHx4j4csfvl3vNwvM+PHjsazlKfxLf9zkzZiGnoaho6Em0n4YaRB/BNXlBjaBIXa
OUSoXXpGl6vZNimvVQNkz4ij3+Fpirw4dycRlWP0MpO5K2qzvykGj/2JRkDy8wFiooC77JA/Wqp2
UCn2VTqVQrIHxTqWR+Xrvh/bEtKcXCMRQHITnwAz33jdL/P81t3eWKadjwzlrt0wINIUrxhguxjY
iwyL2tDUhh0sk3I05UIFq0JGh1DCPZn55Zwkn7aF87+b3iPntBkDis2HGqDbZSkA89BQ/IwE6f+p
G6N8d5IzTObgNA7CS17FLpopEk55V7nNBV4ZNiegoNpegdhRxEASH+fK44XqUr1wvzfHmHyrd3d8
43ulLGPQXY+sX75wAQyqa/8WkXynNMj35AWT6oiEyG9inOhfc99YuEVxIceE1h7gOdAlbv2jqzt1
JBZehun6qquxGCAWA83hxxQ4IHA1VE3Wq7iUtLJD50fdl28vYnMT07wb7WAEVFDgtGBs1EpCds4s
OU2YB5o1VGU7Rh5WgsQ1hFbdvo3hqZVG0FQx2tZNje9LDFHDqHJJiejksQjPUSdGstDv09oc0Y7z
MO7GQamdam7dNyjp+FbkVaV3Rwyr1M/7Udw6dyJRz3/0dykdYETDp4urBZkAmpL6CVIqq+VVn+I9
gpMfx4QPIKi6qyFZCgcNEfXPSLSYIjn13P2JZHixT6xUUWXuYcoB5yChE3GeFxveKMaLESj94v+W
FASCk2pC1yDPY6/pM0ZaxStYVxxfMGRSpZvV58J/+m1hN4xT8LbiVMJNQxUjRioCwhHr78PfUwhv
UFjLq9dgv3ezuTfsAaJhrcGpNv70XIGQKwiSIxU8cLmZGMEOZez4UIaL0NbJJmFsih9085GSiYPZ
PkbjJF2DPThRZfifse8Xn0XOVrysVKbicGI8+EH+fAAappLm55Xcud8Op1WUqKRA27KmakWOqGtC
MaWWaPwzBO8IhjSCuP0jFtxsYG6ujo8Dp/xGZdXPdjIvkIkT6YdkZkW/D2mDaUGWVr5g/CYis1pD
3IFi9Ac5hqedaaj6lIq4kQBk3ECEjvIfyOq0DmhgIMC00578SJ/kfLdYlTWooDTuWaPH18qcW5CA
BWR+IMJAG+BZiV/Vw1dXcRmjuhIDkD2B0j6++kgmIOrVSVzSfroVGT37Wa9pmU8ecqO4Hy1rJnYj
18ESmIiA6HnStjVcMeBt8gpVzC9idm1yWsMw6V78aZy+ItJHD/26hOmyOUjxPwkHjkXGUdGvWcTw
/Ehz3qHiBw+0wV4+gCfe2raxG6HNzW/BNQ3zlYU18NIDgTavCoOvmsxRcS8Pd6A3hLBcK7s0jKPw
LyBjTVhu1tqDgdMBCoeoj6B3UZnTX7RnKwj7NEnSOSzPxOxoKMDO2PreCwyxd7VPAkeWnhsl2QyO
lnJPGPXg9Cic7oje+khSKGlWnenFCWb5H0xyJMevzgp5Zv3MdH/bpLBopyjlO1/f4LPgM6Ni3vY5
UvKMPP8SSQCsv2ikrV6IlLLley4C1bw6yf+qX65qdYuyIusDyWdX5ernkfVPUZUEq8KibivFNjMR
27IGLsAbw7J+zuL8ooC2yxeAx2+TbcVvibNtAjAxib9gaJCjtYDFId3oJLYwk/rex3eer/BdCEK3
xLs7BwfRQ9ml2nroDt9b64crhpGipMcJNGKavGZCd6Stdrsur++bFdBxblrX+CfQzFCtDCNY/rcO
2GL+OIQfMdIU6ThVjUPTIv/uZ5MR5DXVriRlESlsfEeJN8m4Vo/pPGMMTVAv0xMle4JeKoOrZ+RF
NYZc2GRpoKPdqm0Z/dzxb4M9Rbrb0d7naVhImEOB5bqZ+8QNMH50NGT9nyEyuHp4klrRohKMm9fD
ZcpjYqnQ0IlflYwj8CDYGulbNOQ+omkINJpGoHsbLIrbSZOlcw3RLyCi96OIFZIho73Lm1X1ZjTH
8tVyoPcONUlmZElZfXSKTSYbeiyOeU7C7xLVtaI1amtTIwTgmmz42nRSISPT8DxjR5FU5qH1KkEM
vSSwsKcMZhRXTY+Cm57NyHbTIG4QK/qgWRPJQz7ltkWxsyj1Cii54GgO7/uxUqK9GhJYESFY9N8e
lmVkXRNc7Yg/0vIP2qtjGklkOGBhixIaYAiVcj2L1qb4aWuTqPEovajON6e4ueHw4Q4iPobrVwPU
AGvP4uZkANv3usK0Q1fYpRK6gSTXad/HSTmGoJx1PBeGaAmkUGYbR165b27KTT+9xptykB+ZM0bd
+hK3ruuaIYx8dmaVl93kgjdiEn3ndNuGEXGUiDsdoUUk0HshUmrW9nuAW5nZDf9lKTdoNpsUF+E3
lF7PWHQQKxpRO3Rv2+Mm3It07y30IVZzU02Uhsl7Squ2a0ZD3SQFy3k2VFQjoAf2CalO5qJ7gP9E
g2ItrtkqZ+ZoGSLrgYPbvsxJXqwWiVlS5TZQwhYSNIKhZ1x6AzGzuOIDKyQGPhgqnmCYRxcleVFZ
lKVh1fuzZwO2kDWCjjPj2Jc6m45lKpBqGToepFbHHoKsK9A4Cd7s0I5mX397nJF8rF8MyzBqvCI1
2Lp3Pl4cYZjqnSsPZGJ/UrFSV7BKSLLx19rd1QpxLxjiHHGYb49DpVqEKHAkIZFwquQx3fjvLPqf
YUbb/AYqIkalzr8tWjbwdTU8zx3K5KnGC1WcdGTyMtB5+aJDNwOpgt3HD9JsgBSBP7bl1UZElMF5
W704y2wr8y4gQ8dYQZCIohsV7lTRSLDWM3zWD5Wja+vVf/AO+gjcYFJsUBuGWwdGM4ZF3zQN4P3v
6XhHAaaQ5NuSylytkMouQMKki06fEKY+23xx56PhaR3SSZcshmiC2sh6wO5ItMds+oNQAPfeOXR7
j2vBeDGQq10rk55qKjqDs5xMZf1QP+WKhV3ycoXERkzj++yS/IYCEmu5ygX3N+19rOs007GvCUFz
JyKhzlaOhEd1hz2l8QPCgGP3J1UquWxnrIwnJxVOMoQB/KzYqHpuDHlkfZdl6gAMbmgGyjIpK++N
k8bxZf4KYXi+nE/zVDnkTveu1FLXgGu92keqblNjZ5dPtz9ymKzvdnoa1U7A5x7lX07vP2svmp34
u2BLU29J3CqbgDzM5dK4hFgGN8fcgL1A9w+luSobyFbnP3W4E6s+d4xNO3sxt/1rRN6G3kakAPcV
T6fnmy92BmiIsoQisKhE6mc2P1s+NBEaKG7Ne9Ay+nFkLxbCbpyK3x7/bfxmKzbCjVT0u/uYZldK
ZRkbCQSL5OJpAZ521ZxQfyOYJOKtKcHeH2PErgj5ye3N3RM4IU5rwbVYCSsDhEoYOXS8dRP7DjAr
ubeO2hBkZY6Xr0ebeRoy75+rHqoxuVXI2XWg6QwJ9gylkLKHH6YSzY90UnzUujgRgFFUFk/34433
UxjMEtw0L19YrY8YWFbqbybQiKk9mnG8HZyqf5hbJad/yO8EqVm/stJDaksKOysTtKkZSbbJV03d
x2icBdSUv7H/Rzef3vDVrxeJT9qYH/XQlRpHFoRnZUczc+n6morka9MI+gGPV3hSn8yAsDe9UH7z
LDN7wFfnHmAxaIVzD63VEileCO56uaOrra7FRCWavvwm5q9jX2UWHL0V9Tfv5Yo3X4yt3ocloJfS
ygaOboqpiCTbocU2yTmLkUvkkZm+6A3LBJquQxzYYi5AbrT9dY6gTNvisi/6QN913KUNwOMpESxJ
TC4+xcG3HDEecrsEPdAOp9OeewJBKMuk5E/SyEbxIJ65/5lXo2yVuWZpDMblgYI0kLUsfnime7J7
t+GFkL05VZCWWjOsNc49j3pcPvqcyiyiKs8x8UThJexHJVz4by3Ea539o66kWK4mU0ZJp3dKB7bX
h6PM/+Qr683Nhzn3I44qyARt1KZuilz6WsnnDgYZ6RgCk0rSqFVfbj9CEMntu74wTmuj73tr9xcv
b5EZC9riU0PeZo4hN7e40juuuC2Bc5Br+tI52gVQW/UqEcoc728Nx0rP3L+qYFeQHjvnuatvLRX3
FNVMacGsVfnrKszlgG3SZCugL655C4fodS7D4S5J5i/qY+M5Aqvic/DoEDeKTucXYltGMuwkWP1D
a3lf6N1HwUBIukiBxfWxa1ECp7pC6grRgPVlJRVSvBav4rqIP90iyLjd9Ee+5s0Le+8r4SByI4vw
hvYB919zX2wg8ONZH5bkMQ/0JWymCxQz7hAFT+2Snk75JLoajuB/Z+lLny9zhf+lJeOqjYoDzrIC
WolFCaqdsv4MZSjrGAsocJQlkw3aFgRDSTd4l5gAI2+VtB/kEAdtKWytAsQYWDM/AxYwwdLB3NEA
7vRn4L9YxXiBRfXKAvAH5ht7xgVI3UtBlboLU3jd9pWH/1eHkJn2FYWeJeUyjjCRezGSqrUrD8Qo
iSZzoEHU4M0Y33cfc9n6E1zsglArUJaTeYspene+jf28Y3kJ5kwr01FzwP8z8nBLIebi13LaXJho
3RCQ70EtjAjV0L/QCWVnDunHOAIPW2NaENbxRbui5GvUaV5jXAI4lhGWtysY451L/++BkSyRLKxZ
Lq10svubssGRru/Z2JJZfvJXzLMnosK6gLApXNcxkrrYUloDnPVdBgpmw86znsvuCZQPJU7Ancm4
/LS5RpDT629GWzIEZViEb6J15Qj7olZCItlZ1b+HydgH7wPOgqobUK3iW07s2n8oBpApSP7Xba7N
JeU7ozrf2n7ji+3d46/hEPf0irrRy9H9ljZ835iwC8sSCWUwSwzISihu6M1xj9y5RMnyo8dENJpY
RBEncAVPMjtNW8DTyTMjtRF38jgqmDQLpbbYSNJlE1krnqM2P5MA4b6yccu8AP2M9vELJcI6HN93
kUVBvQZntlJ+XhYqxfgxsAKcWWQpAvYn1TIfsKj0//iPUI//aZybOD8ltLwpB58ZZe1DR7T1DbuG
l2XYCS9kHZHI9S6Y/pR7ruF9vaztA7WX8FqUZ08OXeRX1rgOoSrsr7+eISR/YLF8fOEcpFICMTuJ
Fvq08fl+/QG+8TBCUAzF96BEhjiS2gKbEowAxA5kdDy/kH8f7fCJyFy3vRq9BjrFfZJ+mggQBA3W
4k4E4I1qgYcjmeFfpDlksjsuwJnFdBc/IRMMkPgLQiflk7jSl5XRcpHyDMLFmheRKcspqxjRGhI4
waClRhuPa7B2wnOiFwiNd7kCx2mBbdDLitua1h74VBJmt6MDxtchRBUr0z2LkJMZThdgifjLgeAo
Mske2F3Pien+qvG7vQszQnaSL8pI9CllmZ3R6MNnHtNg49TILn12XQt0ALNdJyYV951f0SaSijuF
FK2g23OdcsV665lMcaYGZQP58KOg+A9TJPcY1wmsBoC6jhaVCbAsRQtHcQOgkOYqlmQWUz019+i6
DnnmNqUeVtT1wqWOc0xtX8TYxWDf2CCl9ffqxY36l+YhcxadYnlpNwK2c9wWNWdrr+WciAu11kla
e15+7W4VT+7bGzFkT2NtGx26sHqQSeE0pdhnv9AmOz0Qv26EFxM4N11wlMGFNlFDlYGj2XvG8oyR
UO5iYljyENSeM9vDpO8JMWAsbCALIa/8mzQDCjW0X5/+s6qQ+jERY/0iZZiy/8YPfY6Ctw9LQYns
FtAXxgiC1LjucgX+GDaUfEDqeHJfJM/HGG+YOz4uxH9p0XDa3F0Ye7+5IgomXVCAUqx6fdFTiMZS
fTbnUoN+86hG/yFg/yPAY30eDDqQE7l7olaUQ2Y+EitIiCPLDgY19Y4GiCPwTCDZc6GTGJPRhMKS
3afKW52BddZNlLX/Il6eg+wHbu1xN5EQVe9v4LjpFpwRfQo9B2jylYhta5tjzJbOz4O2JtwcoQGD
ovjBOLLLuVYyi7YJJXbu0aTyZ1Q56lQEcXfxSuRCo16sbxOz3XQXa64pixIn4WYK+4Xr1mwfDY63
Pn3LvcbquIeobV7Mh/J/dUzff6JSfQYzwaL2iBNw+InpgVTqtUjJOg2MBHUOyC/5WOK5Um95a6It
B1gvoTXStzEDhyq9aUg/9uAabmNBqlpubcnMQqVqkF158ow9oQKXloT0N6xs+j+ZsffFRLCgz5gm
keOuJwPhAinJJNWF2ark3TF3S3K3OmExex4ltBq+m9E9Kg1y+XaHp0bIBpk8tAKTCmlaEonZg90L
o04EJTSS+pP/dGOw/UG6Kwr5FaJDhimO7Ya03YeTN1yZjlljj0jHRVMz4LWITAkc9+26J+ygwmZW
g3IDSHNnc2yTFQus7rGwLxAn2jDOjf4MwCk5dIEBBvEvpvxHdnD9vlNptiX3Z2pPF9U5K1O8tfxZ
1EWU7rXxXPulWy8Ml3ZV9VbwjjOKu9Z9GCXf/x8vjE68paWLbKFq20eZJ8XyH4m1IYp+EzuVqv2k
osUHioD/pgnH+UTX4pF71YDvcgERzHMP7xG7d4mDSy7XSCZnuhQQHqisxufFBoJcDoNtDOrxlW7j
dFhW6G6s3FlZwD4QqGPs4dXeEwxpLJBrjGf5CpxJ4QhywvUZPSc55/YF5wEwA+shElxVro4ZveJc
NPOKzTfO1qZCla9PACwndUESN3kYtdduv5T0JaGBOE0fmQLLQy8zno6PIGUWCCYkb+Sy+BJdMGwb
2QZQ9bj01fz8+zIaymn6RkXy95lH1JYoNwEBO/7C0V/0wbJbyl9H7YK4j4Y+J2nP76ICeFFSL4pW
CxnYLs79dRjXEpL0m7svtai1L+uL1BjT68cnAPZ2d8g0aa5Edbg7AEnr8pbv129iFajWCsWZampw
UKuYOpoCATuHxKwgBQG1/GjrompgFWx0dPkj6ZxcKfu0uPAuPdqxsVAsuAHvZS/KJ/YAwpdcW4/t
zYOlQzum2i5kpf3JvNwF+pVVVJVGx4c0pJB/jul0OvNNBSYYcu3sIy+spS5KSKEhoK67h6rwND33
uaFn6squ14iY/TYeyqc9L7qQRIZyrszvpyZRDTwcq6Z+ZAR+Bg6kFHDSCS9/ekYDh/EH6J/S57My
v2/PL/WIaaK5QwTn9TxeRru+xX4gJm7B3ehV7z/0A0SLAslRnQCa7b6ReANxQzBOdsbBjTHNhaf+
PxbRfR3QkPsMRqsPE7fmJFaLWzMAzi7C9HWLG/Wpr8do7/6D8ZzJwH3J/ff0/RtWVkxXlT4BJWxg
+UKNoZJJeSNLysfQlchWly4hKJ63YhPdTaJbAefVtgYoIOmQuWDGn/7wJXYQNktpIKREb6akCr/1
RETnCQhD17qTNJWap6OlWrZzE6+NAJIBFIP2Rvixusl2h2gxYQnIU3b6LWTsK6TdNOwm0gLFhmJF
iFALkM3vhTG0SCfCrFhPY163OueNsR9FP2nY/snTsLP6xuwgQvkWfZgToG1vYekWBdBaX6IvkaN8
tvHEoTarfQV1Hjq1zaPrjiCRmX6k7wATrLxJ030AG4ygn4+vcN6DIb1JFM/uKQItDMZxnt4QS4my
BVYhTPqbd0klzqmec7Ez3sVPHe+QKwJBsn8dFrYvi3uLEyUtTVm8jheKbUPBYwW+zLEadxz2Wmqd
4ZHjjcW6radz9sbFAPiZJ+kctBD6BGjDFb2lag99re7XZ30cZI4onLIHf5vuxcTt7Rij5NUqY4bB
oHwyH0HtVDRgot9iQK+appjsZ4esIQ7eCw5bpokKATtlIdD/s8Lirl3KAGhD/XDRTrr/MdpJclBB
LP8sHVKBmOTcze/S8ObCTZ30CuFtS9IYlDQ2uyHNP4ZvFRLF2lks/VKjk31i8lyC5RVr+/ezMYP1
DIBabIks1nU5CI87E2t3HgfXjQbuKnV1G9ikyc+6m3xH6PmIexCDx6i8Yg3K47Bp5KH9LNsNfRNH
LgG/j9yx81OG//lTf2npBGxwN9TrzZnVkzxk5iEZVxVSpptNPW5XNjCesHj+73T7C8F4mM6D/NON
7McsCp6z5wK1tkvp1iz2tbKrvuroMK2SWUjcMUKtUSAXMt6Nke3UlAMvqvWaVALsmU/vvrQLBEX0
K4fy4XepOgItRRk4up26Y6bxS2pz19CgazyKZThQNR0O34jjPEeILs2yKWet3BWrDr/pzqeoP9G/
Xu4VruPSL0/ksWDhsqKlurpwQTTKTs8YJosi35ZTuGt77jyXsGxvADr/GrIv+/qMmdx7U8G1k0Ya
Wun5XGow+unPR56JWqq0XtiMlnT4Zb+U3p9jPHlwA+uorSGwZRV6gp1GY8IKUjs6Ogt93JJNkx18
QIvayZ70B/rHlLrQAdpnynsJUv5vMLW2co5ySYkEbeulcEMCCgiANNILyfx8CcZignQ+HBXpdsYc
j6fa/aD9igOZrtQrsoT5qynnU3O8lPsH/QL2BZCnME31V+Q9qSE3zIHodEM6mD2zDO6tG/P1IQKR
9V63p22fFSCMOL/CyJ1s3A00MN3lqs9+GaZbmAE2DKKmQhGL4yNfX6AEhx2678Nk1T8dNawtfkGt
AhBPwFePjuj27rf0ewhZRgZMJYVYwVOh3Oo60i32dUl1kK8anIQrCZf8lcU/byINnqB+T5qfrE0j
5WZm/dXzQ8MAu5Vw/5AusoXjJpiU4aPtN3twydK3+6tv6YjJvg2d4Xm0HdWIpvOuves9vvvfcvp2
M9VRcgbYBPDw0dVoY3fsPbN/BFRgGpp5PoGLexBAl42EjP1+aGwJlHafzbDZlRiMsclQypwgfmER
GzLw5xNFpqHGYOtzER4A0IeMq/4e+SdPSu12k3x7exXHgH2+dbEWfFpObMnw+B8SyybQt7GWtggK
fouq6+F+NEMdg46agyoOwxOe4w7F7Q2woxFg4t1eEWbAmLjNUEFKUDN9bv557sviC0kHTxB3FqkD
sh9NKSqHYc4GTunvFxI3aoL4FqGeLTmnUxR67/2uXOa5B5PbxCKv6alcrRSvTIEmcL1Z9iLwbM2A
/e7cySe9QOPCKszBOVD+lpIyh+Pm1SyEPR5fjr/JujYRlNMXeSbwdfIlYqF0PMvSxlsZaCHCysh+
x0RBWAESSDa15Nb+bsLI0cyLSBcK66a6Y+VtHGwd9RatYSjBbx/PDkugUNRKt+Uo1tarr1qzWqwt
SZlNdSijBXmxj9MNeEbi1TEFvBN7SGy88bY8YbYgsFLtUW1nsH2PuCFfcXnlqsnLwfbKSWNmdvHQ
vCmWsFlWuIIhPOSMYR0i03gIhhHzAGvobDIrcyKqHB6xV89iH/pZk4lksCl7qvU+wsIQ9LWORvfp
S6Gthh/w6xWwcWiT2FLQgp1h5Pj3dI8XR4361Fl2nNDVdgZ5GaoiPTHai9NNM/gvzl57PG5A/+9g
fi1781xEsrqGvw0l5m8RdPKamzUjCEZdJiHCmNQfA9ExsxpkTN/PymnOCG0UmtAr+7WSyWyH3Y8d
zQ/WM5UGCFVVc3EEiFDr7lwuu9r8U9cd1vWWpJHzN+PjroJLObrNJ1+gRHrSH5grNGveiYB7DCGL
+XHMD+voGJhFrIfAH52jAlHQOBVhN3UJ9WjMghhliqtxIyynkxr2B11/B0CDJzkesoApqqAEJTMC
ZkgwVc2m5VDcoG6Gtg5ocdpMqUOR02uCvlfVsh1+xlsi0mtI0UgqV7gkP99cKEo8ojmie7VL1Z3s
vqY87HNKch4EM+zO6IE+2fKiVIc3lX4+DWqgL1+R8IheIOa2xaHeOxwq5MJuwR3iGoB49HHpr7GK
8lXD+HeGAe4caDGDtZsBxKcAxEQWa3O6RCxmbErW0J7GGAAQiRdnJQ1JzP8An+c0uj34OBgXGSvF
r7Y3dcDnPZ16xGjXKhn1TBEkA8a4eReXfjNqaObi2opoDA9WUBcpv8Gj3jm4muAaV7uyBYgHt0NC
h7KIepiwJ8+MnTqD2AdoT/yaq7XGH75eAwK1rY+ULW73iojdYTwU1pUsxl0/1dqqkAssY3Wh8dYV
uKokzPpsilElMf/gzb7kwAGUpcRPnmrOFRh6vFV+Q7BUe6I3d+ZO0G/HuXoMOJOHvDXuS9Mj6QFq
HIBa/uTG/J571XipuJPYIt5oFPYOv+ua3DVIbpgFQ97pQrb6ihK62PFn8OvZiB8XDNIcmdJyM9QK
Un5qlK0mnYWHAlfZW2n9YIv48M4iwzN140/PfCoFP/zVk5bvfdt0nU4cPgec2KnuAx3L+AE7Fv/w
+VIf52+yrfd6hRdXBYbRRHe5HS5++499HkmXMW3STFFFJScHz4B/jp6mplg+nTxduznRnox7tWJw
PElnZQ+hCYxRzU9DLCTPwmqfsIuYeuMLn0pkdD61AOxzKWdX+dPLczaUwUGScJeH1BI/hAqa3Rs6
H9JBdVgxhmBWQAfhpKLuor3HHlH2fJcK4vGAi2JzpdIhSrEctO7LnLWBjhOxI4zNZFP3EqGe6MLI
miCp18x1m7y9R5WprPLmqPwISSikMmr7ITFe7ESd36905HRbXeZzxWmTU0lQU37dXpM08zeTeLNC
Z7IQAe4qwgb30csmbk6ANahgr5FCE6duqLr6ZxgumWdAnwaJI52Ny5+n4Cvh8QKXSwlePCTwiZZf
KqpczNsDSuxleLCA5pXWOEAqYC5myECO7vGPhvEeL+cwhH5cqmpDxEk3TrglzOXYuquaQUaVRs9s
OmJKGWKaFlBwgJOdVCaKOgvpyND68GvjsJ2dsygdQ/YRUOjvQ2ceOrK9T4iHRqVFiWMkKit0bGjn
7YkNQTbv62vap+DhTISKmAyb1ohFjIfkGqhLBn/bDTzQ9iwuXRcplUsp5fxZEKLaR6N9qHuDhOgh
pcrcIWUx8VaAXDYrYCwqf4yUzhwCPSSO+gPgre8fsF/6ftjQrA2sxXS+M5RKV7PPUlfvA9s9oax6
X7Wr/Y60DJ/RuW/+VxbtEZ9yHI8ISMwsO/iZo1a0dd9oi/uF9GxTCSJvSGA8mV6fkIx9Ton+/Awv
lFFB0NL16BnBYMzfjeFFqteccHItPw7ge/n8RgmEupHkkK0nN2lq21I9I7WyB5QVUl5RFzu70Gz+
JLhrLQ0QCOjcMVRf9ZE3Nu/FdxGImvvVf2zDTMvTh8OpLPMP1IG6/b3HShTJpcGRPJsvnfOjPJA9
bC8w6lxuukGOMV9SrZ+jgtWXYw1fkJCli/BuqqMy5yGwkL0maEZAQDzQ4EC9F3VogO13Ov+ezo3N
SRqbFKFREIQ0/UPnMnn1NN3wcsqu9B3YoGYPd6C4HpfEHBIjAm4GJPIXWQBzaCzMHUJzsxXpdbHY
UbcMj+WC0179tA2ZcGSl85coOwmaY1TggT/8otYF3oEp0lRXrb6MOVp90m43AJIDUfpcp8yGP92W
q0tzJOnMSDAe3Y6Hvh12NHoRy3fvPDeM3NIjWlkb6HtFN7ncpK3WcYfP8KhMzE3bEds2pt/cr70J
fdFwsZtZ579ZHnys6G/EQ8EAh/8T+lRSnsG2S+soj5TmEDTNrI83hzsstghihZz17moEbdc6DXh9
Zn2nmyggM+da2u4FQkxux3rXWlQVL3Ejy2P+1sALDRBtBw6KkoZiSvXl3DlaKa+PKjPyli6Xgv7B
MD2r4/o01yb/vTJaxRkSXn51AH8BbrJaH7Q/3osFnHcWZ4IvfeYaX+1R5YT4YUCwZJn6A02Qca1C
PMLiPEAhPOYHYW1qu73IFts7muTnYOG6aubPIBXB859sb8QdCFLQmcXTuxJsyid6XgzG0Ghz/F5G
2u65nFp7D+tuSlpGcmjASo0tQ45ChYhtvuPuNup4r7Cim/9CN743z6yUIyDysE8aVUpHe1oXKSx2
rJPA6KvKLgX9/TgwSfgmqLd65/GnkJjStUPGxvZl5/Xd4/+REbggxhahPrU8CfftNh8s7L/+5MVL
wmd+uToY2QDb2KS6IZ8bLlXrlHiE2UY6hfLPSurB7638vBlLYOaBqS61dtsn7JA+oks1tlcq09zQ
INSr6w0C+oHthmrxz6vHNF3XhNFtbpRHUYXVVMuyu4w70RKJUGFEixhnK6EN5IsLfNwOTvBz5zHm
8hV6dXzGXzn+3RdijZInRXtZ+FIxDEybH2ELIiWHftWeMNJ3jvVRc//+gdIIj6+0wBej5ODui4us
e8KNN/EZpKgMv2+mtEpqr8YJ6oaqU5o6wnLgtdKLuWXCSUAR0PIFiG7tf5nKf0pxZ/CE3gUKNMuh
oKeO/pcasHENXVwQKBwhRVJkZ0WSZMB67vSP3BcGgFCLBcN2WqAV5PdvwAfYLyMQDDafV/bswNOh
aW/VG1gYzZaXEQbjAKoBMUuG1McfVdjM4pv/aauJry/DVj5Nc4VlmCZN0gNw6x6hH+Lywe4BuW84
ruSvCjB+u9PUdFzUM7CyKqYOo1lon4lB++owWpXe1e2mTxMY9VPg9xOr/vaZPrEps6J28yZj9QFN
EkxZTZoVp75mZ7xcr/suxoGu+mRzlThdgrgiw9v+pLccUrMkQYGzyVE6VpCa5XdjMvP1hOFjW+5b
WdsgNN4/2pls1Vm/v2UYjlqlsDzUFPADrB3mj5YeVkic8mE280EVTYS0XpHyrzNpeFTUMf3o/3P/
QsOACbsqm2OwTK4k5b/H7hgje1a1eugtHwsAyxsgjAJNAfXvmJ/3AXgr0NGAS2LBbQMJZRpZGhn3
B85PEgtSzfVm6tsKZCWdwTJTlTV8VRmZWaXIKZd+VCFqEPQQGgzG1gkZHSBDsFZTazGyji2P9i48
qciVh+FuCn8ciauna4QejvRootDJ8dSuJBe7qI/T+cDZQwbxqabTkEMi+cAj/GX2hR2DaH34FXRr
hYQqL3EXxYjCAbHPDKkmEcPdbSBHT2q3RLrt03gkgwOxz2vEHwdQtDes7CF58/pSg3xQGRys5vAU
1jmedYkPGYtkJxDr4UMaP80/xKIKmfNfju1XqKVCz6KApdCnqNxp6KzBCgIHF9rwNTD/n2mf/Xgc
CdDmq7LEfsSW5YwrZvP6EmzrCXS0cTRYrA8sGal477Hy7uoOWN4bl/dnp5gmrH+ZAtikBZOXA/iw
pA1DxjLWuagQFRFS1XMKoYiHAAFXn2wHB/9dIRqMAQ8ADP85HrpJz+tQds4H9eXAckcTzUQH+5lw
qnj1N8sEiDhvmO5O8C8q2rHskbA9kzz0GrMhzsfY7VxEoBICx9q5eWT9knrsem+j0N6ob5Kojtcs
zehm0RP4RSZp6ghRKIdlj2QkTU/NyBSw5Mzu+Jf8RxkWRU03tKtslGuPf9mz9UTAJ1O2q5aVo4ka
H76htO9g/pzP57jo2mEQAwoeTh23pz/aA2s85tRahG5f3G8YKgK28rVgH68XC9KbtiFPASE4CMPV
QIWHY0OQBBPf6Mea0CR9FRQ+KquigoZfkPt1eS2tiRTvd+InyO9kaNBiD48lJGASEOMnJ8iy5d+G
MX3K4DipkFsYLVogyqf9FsbiTY4UQlBIjTErY9ZMdsJ5kJ1OmSSybpZQvWMNcKy9lRMcacrdBTmI
FrJx52uvEzemtx/7/VUISSJQ9ewS0MavUwfPSknmauYzrDq0f4YaPYS9QtW6/nWptL0klEvEqwEK
L68H/6atZT1lz1fAFdlkS3wvqVbjU8piRt+ALWRxeK9vepFr+eQrI0hvtld6MV/JXnOM3ljQ2vxp
Mp+KGG9kBwGADwFhQ7BXrZ/9yPB1VWic0ni/eq7jGJziJSUpNZhZXp1iQwBiv+GSsGtcxSbFmKZg
mFi2XfbbfCffBN/O2VY+jCqcXcbv3YEtvr5oB0hTgv6V8Ou97K55GaKW62QubrvUq9r7NwnesatM
9cm7Y4wm2Tv80HpIdlheC6GWQlfv2pPagpaw3LOuuV7o1WC6+6HderOx1I194ZofSf3Mw+S9b2li
xZ+pNeTKmeOjJ7x+XSJn01je/2Ipk93Jct2XY8rY/VQ5lN6EsK/NyZGpIW96lY8jxNAXJ2DMgUT/
OM3x+JtJtgYXmFLoal8l4D5Dxj+lICEyScBiF7rHwjPsHame5CfEJzT4EBNS8S0G/RdYEYYsdm/k
KWkiPV9n7vSXjg+mANGzTG2hziEgH4kYe5qMBpqgihApCjtwGiu364cgFfte9+E+0zvWrulRVHho
RnS0F7nmxXKfKGfxzqnU7GMNqJrJDgkMerMDxQQM5YgdlN/ePl9ABS1CiV2DjO86XE+ss3WDwWnO
EZHR9UH5SPd3V+19h8796udBe8ecQZytPx7FYyY7BO03TCR5Zv0oQmu2jOOC2nhjieEBxETAxYrB
9+EycOxC+tq2BKiANqNmubzuDIjLWjOoEdyaKLwIwDoz1phff2OzNmosI5TBAQe8kLXMW7QTYOYF
SpF8hsNfqR8CovhRCMbT7ftrTyHO0nEUntYbHmoaKtuMiP3N2dOVMa+K2YbMYcpcO+sQyT1vF6R0
G+FdxvBLtrhq+NdHoarCb9sPT94NBkhkIYoHedd2JVB5Ew7qOJD79Clp0GCx+wmA6MfKeCvqCCnv
UMcYZyKofQnjNdYBkXMhqKe3KCxAAZi1EgtxFMLEqE0oBMInJvQgCLr5ih8P6d25M3crS8fWsZw/
UeFXOmLxQTVj3MksgnJhnKs7wKmST8MqrcuRyEM+QVQCoxbY4Nsy6XBBseBTLcAVno/nBzk8SaUl
dYvH3/prtdwOnfbmR/uR3w6JUr7roTfLdNkqSXpdrKUk8w7ooYZoW4mI5PxoyBiGVfRjkcf61p8P
vW8S2Bj3iabxMMA+QEK8aCLPZ8W892oA/k+5LxEqZrwIh7sbBNSZvT7l8/jhNxRCaxhLqo01Th9t
qos4YINnpylu5tR8riTrr2ZtcpJEFf1BW4sVvw2mkDhblIUCS5V8gUu2zH/K4TUh/vnWvbuPtH3N
UUyeFe8OUG5OOZXif5noZt2S1dUxTU9pMM3Xss1fUgwB7W6ArOJn0He97M4q3sxe/3GaYFTIA37R
tj2NVbGU1VyC2EBlYcZ2xBBasejUB6npFiqOuJx1mpMTI0Zr2hUNpLlReci0HSXdxcrQlVGnfrP+
R76DSUM2gkpMaEelTbTY/mf+LXZUlftUxedwp8M4GQ5/9dTPuGf10P4v7sVHyNbWOCUEH6gPDOeG
8vdF/mOypSpO79PA1mG9Ju0Ba8f7erbJ7kZVbBLPA605bCGnTxKRV7DysVChrLgDjuWOacvb913a
2ozEPdoL2TIdLfV7I82ppCj0lG16SqaHKxOt5ZlCrAUOoHLdnv0B0r2voLA0/b0/RAs3dC2FH8Lh
bVAUAxIxPvVLCL+eUhGNgoFVYEQIFwWFFezjqwsIkzOMUra8QkUmB0LiC0ilauAP8Mhdn2XtNdcj
I4ApinKNSGTG7PQQVG35ub8KzuFUU45R8T6L+/EqkKYc5Bh0FnP3573SKhNQkJ1k6yYP29qYOqnM
XnlwHjIC3rlu+LCWT0N/yRlwRFc5xbUPkd1jn8sQJMFMsT5qGtgtd72l4fFNiGu8nQHWxS611Vgq
lgIsFrf/T6nooluVPXv1WqLeTi6mOYnrFrbt/PYmogbGFbgxJZ8muoXJfkl5i0susI7wZRZ8vpj/
isvPk7PmE2/sbpvJQT/qBH5mbJnjj26frm3csn/WiSqjxuuwc9fwAw1Xqqda+AZRXDXYs3iuSveJ
qt3Ga8Ff/+bOc8TLf/Bj8rNXlLBhaHRhp2hkv+p6IuHdk9xcZQSXhlkTxX6nc1K8cX9NLmXwRD3Q
lN+owYVGcQ1qIogSb5zFqzRRqhTYFvq6JW8Blzxu34XntEU7lZgvc/RhBIAq7eSo11zxBqG17cdC
/1AYFSTPajQYyNnPKRDvMM0blLTsi7UvxQen+MYaNHQnZ2PqaDhr2CyeRf7nADaCivoqhziKf3yA
rPxwAQOU8eUvEog158ZIWqXgt5UmyB51y4Z2r42nfWvZAbr+sFdfXhTepoFKuMNzvi78LWSGuRPP
OHs7xp9cB8YOGBTnxK3dGKC9LCYneak6a24ZfQGIJ6F/tEGDD5yNrWPKe6XzDsJt0oeu2OZmZo00
rfI4gEr3bU8VBje/DmVaV+dDj6p45YzpmaFSxlsPHw8bNBfS368BmBRYONVc+Ymf60oRoq22KpxD
xtRaFKOakt0qKi1wQnrG/YHptxbBwTjXbQIwBoC2500R7FNrq0jZZ9RLCy3DJQcCyMVN+PJRZAE7
cYubiD7f4Tn7RnxWAn7D5t1v2NWYFk//hiaiNygHAy6nhgxfqB25xXvwMMBDKZ4vF1GkIVfvk/tZ
CBR+TtGupLl3cB7lupEnqv0az0EAwyntukNsmfOeXDCNhEHRvV32fYo+sB0APhpzTQKva4waQ1yJ
/HIcc9OdxA+hI7JbaDRxhljvFbRBD5YR5v4WL9WMfCp2pyjB/wTV/2ZLptkDqHwOFgB5iKcJk+tT
yaLsijw1dHKIUd8X0XShCdB/mUBVy0ygfsaZtIx96+FvvaYq3to4tqkwMTVZvioGuFHKrT3lBprz
e7fr1LlczddTSpN6ZJB1EfQwYrqjfCg4WjjxG2hEKBmo/I7Uk35ElP0cmZ0LuizJ6nEAI19ZhY1N
eQkJ1StlFP+o6OTGPN9ud4PpWX0N8ZsU1/vWSxuthJxD8W3jhDcxHPR3JtZpLULr2ZFJgi4KQodf
viEarD1Ap9BBPhLEYEYLfnXEyKPnYYGaE/s5tvFXiT/O+EDiT3qoZdqwNgYAjTxHgli8o4wkP4ms
mjgIpKYEryteimQzZkuBPZTvyHE2dbOmKTT5jOG4Sl26sVRatckIRiywkmnMRcGxXt6BRfTi+Jzn
sHnQ+Crbtww5KjLqPG8vDDXWrJkLhIRJ+ZhLzqZMR3BZ9eNtndKmMfk93fPfvDEPU9MUVefcdlIr
r5NmZhmhl6JaAzRGp8tKgatbpiaiF+lZDKBTAbXvnkfJJfawWm3sVYhQTv1HMMlLQYXNuj+rsPQH
d0OJjjj2lQ0sYEI5kbmPgnA/1q9/DXz3+UAF3+GZph3iH+yE1HgOwRlY2rRgCSqvqUyhGSoELRtC
ZufIb1RBSaJCJNxnPKI0ViT2alqHWK836yegKlmOXh5LyA1pkRVOn3K07YP3qwtcEkH8inZ8ODrU
zN/W9OP574znIcR6hPY6/sfyoAcCjz2RDNCoT1L9gY42xCpHk847Kx1Pc0lszUS6LaVbISqwVyrA
yoe+K+V78R7uqkdriG6LhY8Irx7IXWr1BR5QufjNUSQ3dH+32qhcIwJ71CMwnuMdSaGyeqgB36mz
kQowsuCp1cCwe7kpEelI1hv9FzkrYWjcFA/ot1wBtqNqtDGS0AaUK0fNLLKfSuttJS+4736AEgIK
vylxstQdZkismTLZ812FtcoaQ6NLIECPy813rpj/tRlYgpSzqzPWkBsY5mmDlvkry6oMvPpChqCw
ZX9hUCgK6aBT2MB6N1lNTUUfKsuy6JU4bs2UQ0uaF9XJYDhi446M1jsbDRYYs2FCGu0tGh+qecvN
nDbnMLMFamELPMeehe1c8fSj1KgMwGffxAKOR1+UEqGE86ahjby9QHP4112FvBYDdmj9kHZNOMZ7
iWUqaKg6+2I+X3kcFzZ0r9IoyUs/EIbdavsabh3uFaLebOTu/dcUtgU36Y2sq2GZb00/9HfhyMdQ
wYwRLJzOqTp/9zFEzW4RFvEZjR+rmkK1CF+7U6RAzZ3Bgt5oStoPEq0AdGjdojxt8LXPwIVlGO5B
vKQ0PKTwgt3ccxjtsx4swtWF8V7BQM+QoX+ypOiYVHRrCXZxjMN93Jeqp/+t+J6GkJa+bRfSpmsc
XinJIfTzrra7irJu091L4WYm6zEMBd6vQIPdtmPHKKoKNfsRHj/n0JDDdqdoTG+GZjws7oGxppRw
VG08scUU+OvGDUoVCAv7UZZJR6W4BdOTiKqATYNqEhHRpbSPc//CDgVQwJsqlSai0NW/69nPPUJ5
io+MBabKdhDwVd9EulsCBGhPfSI0j3/z490LbCCLADLhAuMg7fSnbPFW2qLypTaVn7fwvZwNyiEv
L6fpzwbU0PKrcHc07EuRbMK5ccuj10mBO5Xn3ziHteycx2zxX/e2AgDqBl8LnRa13bxIECbErAxl
o/h6D6fKf6g3u4N7ZoUnbhq3PtBw+KlkpIauDC/lIaEZoFUyUfJFpttqk6Dg7neUl9iOrJ8DtIDj
VcgbYk36SOfsrpYLKtFmsGmIgWIy+UY9iSK/hqXJ5XRTjKskGPEgPlyHRBrnrYuNYB+LwG/QbqCu
h6/a0lEEzw22qwfanl9nL3c5mTEdv82qFdwO2mTESMsHkmfYfYU+ChiMAqAZ3aVqRlwdVy3i9J4p
E74h36Nueigsw45n085eK6T1imujRzFBALL2nmjBQLRNHzjxqTn2TLptjtq/gwQAatHfYrW0EZDK
xH1T/YCGH7oMpZwl+B+EYLc6QQugO64te5hiYHWYJBFYvLlQNxl+JA2ztgn6Bp7bybEvsJNMia6j
ZYQA9eLuXH/EW65uuy8txoiLn8PTseJ+n9QJaUxXf3XkXAlyIk7Cl4K/tKEEbsRcRcfipGBTs0AR
90r/69SGRN0bPHyPvXF/LqHrwg7FEDTJafPxPFoCwfn9/GzSNUYJYNFTgMwtkQvpLs31BPNjm/6G
n+MvDpYEB4UhidDdNDG4+1evgtBUU/wIeQdyZMS3eLg6FRbYgLZiQEa2W8QPoW07QMT6whQDZZUy
hEeTSPBYqOWoCJ3mOcQTGjKaJRaktACtAXUTR3AryeBUuZY98kyTV8OfrLFC4AwmQzRkVQKYUz0T
qkOCVTxjyPskL5tdufYo2LxmbvYgYT8SwYHNwPbpT6KGYxhrfGR9vEoO9+Nj9yoWs7IYNYaIjvan
zH70w8r3/kSemh4fJgmUku0/VTIia6IMx5Syc6M+tsdghFh9HaEucU39VyvHd6S8uvdSQA9MjlFr
qOmvNvtvSu6gaxGjqOK7RYyT2644Sm69q/UtD8yqI2RCWI7w2DtOj7ep2O592TD+1LoY+WkecbPZ
G/G12tq2xxFcwHfIcGjJsGe19oeURZouMYUI5mtTlai8yCGnBdJCJhuYuvOa9ONeJmNdtwote1wB
i+DQNHzgrFAwwZOZhOKqQBgZKo3LNxplURxIYLwXRyb/YF2+XPXe3xojFAwewiWFDZZCiHr/BQIX
7u/a3/NKpEe5xdC+nk+0kDbnknguXialfcrPy52juk/qLPXQ4JJQE8tkfHalaD+3WAM9fthosFKT
Sj2k0sraybXsf8iRhc5c8DdoLlflpuOzaPUhV/JWNjaJxnKcxPuJgq4+LmeBa/MbA2A5SfU2wRUC
YgXgpv8Z+v/ORKG6zsCsgTUfBxKCg7QU3JE2k5aZRXNiNbmIgUPI3xWVtBF7Q3xG2QJvtgcZq4qy
yWvCsX+zmpknNgvD5i0SdORHgxBoCQmRH8cK7JrHQfVB/60WQx5Cw9kJcqIIRe6kOpb+qzd15Sx0
MXjCPOP1MMF7GxU4gj+2mXDatFabGPr1AKJpFoI5RcS2C6Hh+oTnLrKMtituJAgkxOS6c05urygV
42mtfRJ22qoQHIlRV/shRNhGjXc4pG5dasQ/KOYEYzUN9JDwA9VnNKP3q8uk32rH9OUgyvnCpO+6
DUzLTmrmfiNr7Y9Ox3txgFn1yr5GdmJvuY8tFZJ5/DL6R7MM17UvrRcoYCAD2cgx+HGw8Xx+GO3b
2QpcGK4+RHp4vxj4Um9IHsRnFLaIHpnf3vTaT8wdwu6LtDtkjaXJyrFwIZILNt94B/hWlO5ghAu/
/umAtCpcB0g5aYAxbcM93JZIhd7rauIsebJ9VtYkDX+DUXP91vhUEklFedrXofl+jLUM1Zkzk+Od
FGRegEEH9c+lHqQZ1OKr3I+jOnVDBA+SYdqjMbJb7lYHQilgPYcivxNHIzwID7MKNNlf1zg+Sux4
eEePlM4nFlPs7/hM8nrrF6PnGuKNx1xmeRP+iKGEgceCIsle1tQvdFMkeLnK7nKwfrj7diZCk6Vv
I3VD8UhJGPdFpmornaO2/pHu9+WQgNBoq45kStmsj4xvx1ZtLj5/KMDL6LzHnUoGKrH/8eeycZPc
TPfrsm+3J2PxljzQmtaNrB1dKEcWQoWovHiPPH3pwGjeQyi0hbXrkaTlHj6Yv6mi0tsQwu7HneZR
WRzmYr0DLayNlBFy7POug5cnfD3/ye/l7nA22PP7MFAvurOddsDTrlLxki9l3v3WHMv/DHkSXHh3
H1X9DCBi4di/m0VQrg0mauClN3VSNguwD1G9zUh0Xcp0LtPBZVEyzH1eSmuNp4APQ4m4XOpFUhUA
zbZrdmq9YDehaRUt8ZAie3xxslICFepg+PFHRvpPCNNdatLWffb+vPUcEuv2br/awgpWnnS3F+n1
kZ4uKiGsJ2xiVU6G89mSloZ8ZbCWWzR2JH0gjdC3ONptKYauyCpN1w/IKkDKWIbe5bPuOOTTOxIK
tPbLDKmDUR4EjYCuJxEhHHKQrC1m5jd61kTvfpHptg8j6zluex9SHvMUIuWZ7iE4ZbgDBSNpoxCh
sfJy2gRofTeQebHT8J2rnB9e2j49cKJt6lDQ9v1EzoFuj69zbW8iut07guV5/+ySufL5npJVW1BE
95tLO1tvcIZhTiNw61Sw7Y+lDSpDZ+RFZeiakDWHTp0ly1mIOW6CsW/PlrL4UU3l4bnSBLUI4qeh
rsuF4O2qZrwGIIKbFFSBddkB7mNTmxObtHs/B8dKytMyubTKUEU+dAfQR2vwry9CzRvK0BfVwSZl
mCsmgsQojepRp6QoGhTjDTKImeBe9uvGEHuLlM9KY+CDyg6mpoh/cYvJODbD1BBHArCCktbjgSMX
ooM58RPxGxWE862sNS/4zKhaZEfT1T7W5w49c0bxawJ2IhSxthyjP4XNSkQwXaC3kgo3XlBFSYSF
Y3xcF3oEra+HbiM2bhsoH9v9fpYxRYgvTuU5NmxC26pqCRaiF73HHTUugxotXkGx2pJylH2lL6hv
bhLX218w282VzQ447NWpMzscahCG+hQh8ZLSNUpYl7UlYETIK5CW3VDZXz7wu9yFcX0zGs8641sr
kg2eXRtLH22Ng+owJ2opy9/kfJLrzx30GOWlgDBslqZ5Lh6+4+d8vgysDdMlFfjXcO39HBEFadqt
ZtORtllRS5yRP/VakPhfyqgYeypnumrgZrnhecEIQA7/Z6YjwEkgaJtBCITMSN/myjn8Qe4HeM6X
5pl5I5eYtrV8CMHAdqCVjxsi3QlZfdruuwJ73yMWdC9+LnSLQqyKmz0XHsbFyz5jSsFc6prL/NLB
RbkrG9ggEILqxeBClrtV0zfMibuo5pg6JcJufqwnJvc56Y2y8zxjFoQMW3YHpLY4kmSAqu3pDQ2f
9SXi+0Y4/ccdjDvZo8HxpHCGMwFuJCLDeensFq6gg/7mzxmTGdI2DHllVt52D7dAOVvxWR2SLSIy
CpqiErIffXydVja8RI0lvdv9swMQFoYcFTTP5aEmWhSiE5GNDVDRXevtMKyIqFRcLCejx3CAlaZw
19JI/4MCIwOXM6cTo2Bx8Y4CorzJQHdyQGQAixUKt6FDK2YvZVFSh3bwfAr2UTpUc+7wYO/t/G+t
rg1E6NL09SyKfCznm9rCo4h0hKkJFnRwAg89Ny9+4g6uv6+c2Mzgz7qaxlFbWWdpnFUhfTfmtfTb
tU/ydAA/f4NwyB3sQMa6p8tM1atWD2MRHvDh4pcFMuPQIzFWD5OZbeZvhUNdoERpFI0hP9TM/E3V
/ir28RKDiBbD5k8ViXEtsZZNBAhTkgBmForTH5g2q6qkpWW5ifLUY+RnYzTNudIeV60ce2EZ+at9
bOSe4bNUG7iT4QtUmHs5AWXtEAsKCNnlKO3uVE+Y4+LNiA4oxc2sQ7GZvj3jUWil16RLgsEkKs5C
bxwt3IawQhy0kURvMJHbyrGC1/lrForm8uWnh9Td0rnFtztpur8ofBMM30j1NNvxaH8sx+RJC+5E
fk+ipUtxTIr0UMpw1QwqB8nbMzifp/Md7p6RyHnET2M5F7XKkZ/lDkyZuwcSVWFPAag+L3D1IUXs
9J+7cfU6IYIPTTfAoZX0v/0yxkYdBG2lezH0kzFxzoNX5QCT/spGrH6HNHnwKxrzV4oSy2U0B0ip
pQD30ui7tRIRYDh5IOEqNPZxOt6QMWSvUsc06xJCOHcpvc0QCdA8I5oVB9knlhG/VSenjwX8oxSY
NbL7jqzju7uFmqBe/pCFevW0U0jGofh8UCLykb4tqnLFyYicQVSZAagZGiPQtiAcvI5yJG7g2UVg
9t45zr+Qga4MnYTB+Udery9rj4w0OjOjbRGXAp0vpR3awGaeUNrA96MnUJ0it1FCN47XXP4haLJu
NQxP2B7+5FQIl3Jy0j8AXwY10/QjsANwmR1THtIgNtZ9qWZKcsE2pGUdfJ8OAew/zueTJ+ti7p4v
2eSeiaBH6qdqvhOdY64msGOiAAVzSpvV8xLzNIJqHl7u/e1adNQB8Fe6uxPm0HFIU8Eer0MBHZjY
idWwURSnNysYscG5649Uqozk1WzSO+rLi3I2BuijVvDNIqxoslIoJ39QjxB2sX029OaS9l++OzS5
VIYRIUqisssCkN5ESL8LvhRYOavxy+NXkSRBGkwksvaYqgyyQ2dqEpSeflA+geC/3BLudC7FEq4q
THlIPNqD+I2ASLGjbCtxWeIrpBeep2pJA1W37yZO1nLBAYvd5qdPsc/UEIFG28JnBU8LpSDvEP1r
oULvIFGXPxPHu8PyanwRvzRjePslVhHyzR4fi2VbAr2CgdRxOUs2AIsnpg1UTZIhQpaPrd+CtFKb
3wYHsGtPuhiil9XDUvOiS3/0o6+5z0+Ij6xqBoRjK2es3Ztqz/O1EbiokT3QDoyD0pWAMfyS/7rV
H1EMP3QMOfM8BOC1yJGx8HsNWstm1wjibkqmXRdL2lMxYYQYo6ZiFj73xFcs2QKHO4qU00MnsfXA
lWk0tGKkMUo7xqzzSNyptx12w46QqY39GstabRajgFj+MhHbJ3g5ASO+zAaHDcQyrd+iZ8xgu/eZ
W+lpJsaNBd9uQrJcM8J/eZG+TtIdUhAwmeVbd624s2TN/VF+nqAdyCxhmtO0NHwqZnMjwHpH4gcu
4RgELO+8lM0koK5lqPsSAk7NsNuOgZq4nen5sXNXkysvMC749fLkAyZyPIOlj+GOe6pK303MnRUi
9gNq/905xn+rZauBeXw2WyTSPvwyDyANhEsaeR9Yj5wxmmiq2/a2Hi/WfC97YwMCCXmTji+84Ph8
PfgVQWck/denTHPFNktK60IeQ9W8kNW4Y5XrUQzhF10Lqy6SxEGgDTAZY8u2iHgpor5DFiq3QwHj
W53aFP/qKoBOPdd+ZeMLNhdbtAg9CR+ymUPju/IqrqtPOV/KLS++2AMpc/zCFo9l+0A3slXCvDDo
EEsMDcR19DTS48uXdiys2Ctaj7rbubPoAAmaTymyiGGvyg/o1tzVCuosjgHDXbF/w5J6XzKqiEJs
sMHOI06F3iDyqI5eAF1u4ctUYNm9HaDgtmxhi9S0yVpfLPYatAsYVInqgWKqQZIcoVF8efTg3sqx
L3tzE5BQw+4YpMFL2GI1OjsFxoCGcYSh+sAIauDsmbN7rDEsBT6+jP78jtHr1Hyg+Q9iH4UBIu63
xhcKWvxWPb4WH0EmEsB2lxGV6jzwEUpx0b76tiSO3ieQTBqnaeOSmsuZxl97sTg4cwfUuBFfh1rA
UBnWOjgmg2c+5OnedeJLK1rpP7PIlHTQ2Jx00GJfDcO4gqzIwqlx+PUXDPuOgFyFWKl/WW/HdNMB
KDekmda8iDjNtkP6X3ss+AQxOzqVlg4fN5pA2/Ywq5NkWQtLVdWVh2vMZJGPFVg0aD80F1VjfU0m
YToKBT9bDsP3vtL4SQ12HyVmW9XVHVNywrVQYeBRpWN7+ORSXoTwFnm8aNK65uGQ7V9tcnwQtbPJ
PIErBxHFy2V+h5sQrNuuyPld4z/a0J9Kp2ajjZy8VYzxbEn7Cjj217ndpA2bsc77z6JC6OO83Bnm
VIvTi9TtFfr80yugMvZgvBX9GcHiPTbvqAhygZCFrAtRtVePEldvYnS6vL/0a/zsOxTHlu5IIpRt
f81UsaJ9XTBThPabRY9qC0P9e2s6zTFgaqEtOxkDvn5sITzOgzXNPfqeXBlpViW25JAwMNIuTpy1
9O/VKC/CAJk+NijEXvJYLvzzsCYkrn8NTeWgDr3CZS+EkBnWDHuVujfocaOtm6HPntjdifBxjXOn
OEFb4laXqio7DN/xK6abkGvINVpSFSh55J8a+iA49TKAhcXDUoIdlfBbpjlRnCPwIRwXox984ePZ
xeTMEbRLWUL5VPTl4mg9yd/FF1hDj1V8P6DwwcNhdxdTg5oNm35WSxfRGkDwpxi2DYBD7+rUlNil
Unu/Iqry43phccP10joUlpUQ76OAnvbrUPPkkAESVV2iPE6muR18/PaKBUvemdnSIIugDzVuc1/e
pMfJKh7vPbWnNkUJ1RxgCsykH0rFSzXdNOnnPo3RFG316+vw7gGyw5cTjM1QvjYxOdnJQ5QO2YTn
4kkttnS9SNP5Suh0z4GEOTPqeUqxh/tXlrn4bc1zvOi2pe16M8twRXrwJwpRS+HXjMWVxrb8csR4
lSOlVIASeO7LILje9Ai50F77QscmsJLW07ApBUAUT0+z2M4t+nDZ8TbB4WGn7UUtxGGw/by/C/K9
DzTjJYq0FJoSXMUg50qskDPJWR6FiuPM/sKaUpGM94r0CYceAxwK7bqlKOyqZzIIknXD5g/w4UfW
u2AF6eG6uWo/mbWlf+xKIgMWMRs6I55OSAdrW6BamHEUUsyEfY7fdZGm8EurAghuaF5xJiCfHjnv
MnnWXlXyMYiUUvJ3rTD6s2xIZHV/TjFChQlh00DR5HsYghDFphTHbyGawdWQJR9Sho3h7Dwdkh01
fyv6XXLviORD5Se7KHQxfjZtIaWiMeFJvkXAqcpRw2L0RbOgW6YjAvt+hsNIy3BG3QqPhqg1N1mj
o4kHTDPoYrfo7Frj11ZDFINNEXz66etJUzkmXh3bZLlrhuNVVEbfs+e4D8UWIlW6PB7GbKc/clAz
sT/Bh5pR7VaNaPWmJYLdo/R0kJUnBVoWKnpif0VSNoD82CY3r/Da/OwCztSJrGeVoeDnhPhWK7m5
BvZrvGy5iAbd2YeSfj0OYhR8AFnBjRLxPTTMrl5w3ahmgwyI1LBwKbTBgffdk5cWDHWeq6H/NEWU
+Q2hYJmKpXySwXOWdl+JNnRNSC4nP6ZwF0UE59QrMokWwkTiMYL3n2vo0Z/WiUZjVyh22pTHcONg
TWldIbv8jcygjWQoQkYWrBOf3HEj9gUTVPY/xOQ8UtgzJqZz+nDeddzDRz3tGdsAj2wYnF3wxSLQ
0g8K9i/GmJ3upGy8214UuX1GQGpPjyVSTtUBPhPfonJ3HeAuX/+DRUySl8wxOHxQhTsUh+CcTpjv
LDUD22K9TnvcxcHcZPzy4JYEH7owiimE/6yeDRPiGHE8qWYgXuiDNpDE4yoPC1mPfCmPS+v6z7/o
IeBECs+W5kM79lBjS/eBIiJ6g0IObzlKgaFzC7wzUH+BWYIKfVLOpxQ3BYAJXOqSwwRV/xufeWY9
ptp85yENXPJgP7UaemONLHx3niP67YZQX/3rkATR0mNn5SKbLGASTO5LmyL1fjicdJP7Vj5WuLsW
p+H4C2LDjOrAmyY+aKAhy5R3HHntNwn//od7wP3lO9TFTJkLMzJJsT6yqaqrNFVWagqRi6wXtwwT
+X1QjcvU58XvRALwQqKL/UeZ4p0iYca8Ace7DWt7QqG9Y3WVxC1Mzht5ZgAyvKJrWbq8gMAFmOVq
g8Evmv/9WP4v3pG2bYtk7sYgXUhpV0YUylogGIf/nk/c1SHIG1173qsVSEa0CLJgDSp7qYEJv2+j
T73KRjqQWx0G83FMUybjrL0awDbZ7M4J58vZM620NKMn6Nn0bSQ3fv6BvXLWIHaQWTINh2n8/Hb2
pZ/0/oK+U3jaV2Cw9fXJIAd9zK7GK8oLlbsIhb5qzoUoCvSa3VdYy3NRcPvv2/ha2Z5JJl1RZhAv
XQeNnPRJimiQgT+5rYDFVNO+kXVwPh7piY7VxZ3QYBlM92UmPqNSLszXFdvpwO+2bkOW5hM7hxsg
FZ6mDt1P5DdkINfqmSdaw8stI2u4OqW88Af3jTcTVZtGeQka8MKnG/0TSCRzkEsZNfYbJ7hwndqG
CUKrgRPLeORhiKy+JbQRnThzS0j6ysHqR8AAWR/XDJGKlSqy4ULK0Nm6YOGl4CmpliSdRV5ntdpr
e5Cf5bzS83XMOf0SgxEgxoT01cb591JH6EuqZhTv6DCYGV74Qd3nS/9UwP7ekyvrFCGPf9rl1yUn
cpNJUrF7CqK/d4hkE2MHOv4C5pPwwIjkDO8tffy29rk0RQxaFwIVInj1chcLLMupNgWpinuty5dI
CvEP/8aQTmvo9b89HCFRMIWQ275nL7zzjBiSMW7Fo3zXYQq4G2tkFJcFUcvaPOQzjAUe4d5zutx2
xYOQT7jHUdXWZiw3gWgiz1hZ8kftvJdDR/EslT2EjsWyWFrYOM24qpHfEPFVgtKsYGHFTcmS6fEv
yRCzKrVnlUbDgvjNFu1wPyP6KTE+6Xvm+nvyv+wGehQQXvfcItp5kvKWhFGnoREX8l/zpKlK25lS
pvb2vteOxIHEuI0tAKoRGwng6jJutyUlISILFGS5FQ4nbto45gfAA/t6eS719Eh0ij7R4QCvVuG0
W8bd0njbxg1+0Ya1KIdvQG525WQfKuQ4gUMUc1473+nY1f6X0cHVzWong2IuxEelMO2gbwsHSCRr
ad+IM8yucdV53b88siwDs5mxVAQ4IYAAF0hVxbmxw51JJR+2cfT5DrYPuTE5Das4zucsm6Rt4Bms
cp7EUp04ihsm5yZ14PcNTTiGzpK2VBkInBTkHkdNRM2k89wtTBJFiTqTZJRKB6FXKArwbjf3+S13
tdfKfWrBlYpN2wQjNwfHPlUKP87KQKEId0QxpH/1L9RxKbY4fjv9Vv2P1yyIg7aUJHU9xTMvo2vi
j0GOto5asya4n/KHc/QT2omRzjLx3JsaZGT71E9mU3FxeR/VqyXRNboy6bZjOBrfjtBMXfg3o69I
/kc583qoUYm/8s+T2wP6XcntFbQ1Z6v6bHS/meYpeLzj9TfNzjTYnWqRZvMW9/qXr6V8GyX60mQn
h/1/xlehk3Me6ajzQjOXhwWxKBWlOH2ngGC7VqwZU5ojZpY5m+AmkpkwdOGTj51uikdo9Co32QaV
usRNcrIkU/K4+eGvcnwSe0tTBFbIJM15pN/zZ6hz1Nn1ur3bHJ0i0JAC94mviymzXcoCPobjpXir
bImajh2rX2H7hC0DvLfEru+6qKxYhQPg9MhNqrRw6U9gWZcqi5iyDui/s1cFDXrJj7HZSQzMlBsv
1jQt7yIrqMN14a+7tQwnr0UcBDXDw2WVUOMP+ZzMCM6O/ibPy68Id3ZJGyTm/4YM5q3pY/GnZdHS
mw0mjDqEfBBQi0UqGGHnq6HwL6uzHs37yMETip4w0OXMBFZgSONT2ZP4reT10t9CdMVD/1L8BLPh
+zTDj3zpnrlXsRjzZHcQwlqBsywhV09BU0X3O4N2g3Yq9S6eneE+6oQ8pi1MPzUmSo/iUsI9yv1N
6pUpKvtiVkInbaWrwDI4jBYnAAyLutpWy+EYfOIolNOmh1/J8P6S1pqfV511+TMYt0NRDyAc9Fp6
y9JvOHvgMKrB/O/9Ddoob2mQ2qbndW2lpasBussAxn4TV3s8CIcHh2Vr5c7zH0NeKVmZtkKG+YoR
lvHOoco3CSWxu/zxOuscTd7EZAw0ARxiLeiUqxyLffqhPSV7EiIonhR9KnMeEVm/kJwWSlVVnE7s
Fgn3Dp8R81/4TvG6AoRlANCRl71oOG+B4l8+TiMoorTQsZB/VQN1ZsO1bB1MYUd0dbJAZ92slVmC
io8e4IuBX8fi1FzB0B0a3dCXPKctqcIudyye37E1cVyWmT0g9ABGdksIk3YlKdShJhxGkn+VCisR
R1EbbKnp/FbVgyEDzJZy4f7yBPJoFavf8vfweBSjdR3kmao1Rt/UauWkZknVsMy2lISaBUXylLu2
CuuOzhaLepZVN4zcI9fCVIz3Y8A8QtpFAk2FMzRSTh5QyYwhnv+y817/+2yZbHeWgMH7dD9KWjF7
8j5hXNoXvonpEUo93pu70q45ok4hs0bvZnKci+7gPAxwa0uU/2mgQAXTIw2Lo9+Z273g6gB+K78b
32v77vg3b2Xlmd2PLYM1dxF27ypPRMhdXDqmKqSlGKY96vNd5LOVUWUEzj9+fSg6DxyrMXzHK6Zy
zvWsvYnaP63aSLjHiLsAGNM1zMjs/anLrRJbsGWhdeoqvhY6AFTnvs9XISvrJ8uK/1p9StdRr0wm
9R2KdA7bH7T/tbu4W7/x5ml8zguRl8V5irmZk9APno60orOTL95olrwMI0IkElgEmg3yeCUEnRz0
t18Bv96/T/rAhYZOTo31u2f5thCxiXq5+O3VdimZrpn0cPVd6ueclqbSgJnR3Wtjjo9D2B3RCOte
NMBqYk8oslcFZu4X5w6HgO1GaTQ7lBHkZuQXnLYcsu7vB4dSSxCFM3Cb02KwK/Vm+gcScJ+NYdug
dOyinVNjjXbATSK+7H/Q59ZGCB10BzuNVNwZ0juOoVQH/Rogcd2m9NMH07u7kgngNUDhdiNpP/c6
WQiMK+7EaTLus6VVVeC+JUl0FtJwCaRyPuYZLkZU0tx3CJZdkySn63CHBGWuvTcHlUNtJH0/NVPf
Ix8wcM6qzKX0xdFwhqrwX52Hx8tTCyk5eBYNN76Xo4nMjBnknQdkpQITSAxbbNhKyTNBYoij0lov
pgVGsMS27osKoPD2HFRDJzS9XPGWcS5IbO9V1njtVuB5FCIjXt+QL6Pnwin5td8wF+2LkSubOADJ
Q2LWBNpY6X8AdEVHRPEJ9qLzbzfnO7RLh0Fx0/xYpXqtDPpH3xJsbM0Z/tFplNVhW7mNwp2/zeLe
Aewo+giR9sXImzaj/BoienkiS68h3ZO+L5G9FZ6A4vtpWbBD7k+d05pBygrvFzd21z85FSFRCpc6
rzaWb7i/QTWNkM3AEHWpL0fGEJ/zYV38bhAQ6vv2n7AeSYAE0Rp5a2fyrjH2P3vJpROOlbL1XhZc
SlQyHG76dbWfuJMXAJnXH3VT7AlvhamnEFNi9psIxroHf6ZdKRyjfI9wDVGKp9LoHX3QW9Npx1RU
feiXSttUTlEcmhuV9P2g63jXoLpttIR35RhIorUAiJPZNonVj/8sMl5gG2mCzEPtuHqMV5Xughkr
nJDJSIQl2BEdK2wEx6nNgT9Cetk5hKxKBkvX0OXRPkw2eyhVaGEEF/XmVXHpVw3DsCf3cTG8yT9u
qmynJFMPxlTRxhGr9Xd92wlIS2hePjlYrIX4rnAbYjCgUpHoENkkBvNDqvx+pTWtdbbpPqG/ET7b
6/AYNh18/vLyhpFm/tH4VkGpz+yiKtyeBZmMXKRp1+GfNKNsvRKQVGJ2+4Jp+qyLv7TVA7gpXnEF
XkCk5RUtfjDeey1+1LqELpLkAOiAivUUlc6oyuUGJBCeUauwX+EkFIjIl8d8LfiZBLQ2U+lbKaXC
NQNmdxM704ECWuLVYwSMYNNmI26reGgsaCsJtG+L5IaFj3UytFfVa0W3soducbrxX8oR23ILB05S
U7zJRV5m7io+H/c7M+xV2AA7HriTAZZmmW8SgOXS0A738BCKx3ywm/SSrULBcQ4Nx31Qj9DdRI6+
hZtfQUqfYbbjyoy0K+u9ZVTEKokOCZWxAF2Cp8TC9sRF7ILKfSL0vArVdkp9UUzP0PboPnerXhnq
juj8qNtEh4OLee2u0XQAbulPi/2VcReAbAhDQ75YwISoJfHtVuzPMMQEoCiBktcfc2DdWyWcwSM7
8ZSDIuAW2Rvx0vc0ooe97e9vxZyIQmifjgdn1QUbaY8iM7Z09TQuPQF/7PukfY89cF64bth/BVuD
GwyYR6nzvsZBnJlDO0T/5kO4UoXO85aRyTDEPBjNyItsFzUHuyPTy5KelqFujjos0owP9S0TyhSf
PH1OkLcXnU/BfRcf8cXttaue+Gm6IYpqJ6blgPUu6U+wAAElHhWjIs9lsHX0anyG1hz9LAapeyhx
d43hK4D0rfyHuBJsgOBS6LkgY03kYKi8rjjhmbXtpgtdWbossodvEMQJeOwCPsu2gS12FCb77I0Q
YAb3wSROlMaMF5cT5kUHeD8cNqr4CHrtr1GHoTdUgElnM+pYWI2OxQDFnkdpp2U+6p453ziZGwiB
+8Ygj2qq3craVOMCrHk3qCsA2MPLm46A+U9ftjX578Kglv9AmsW5Edg3zTXUQXkTUQispepc/TjA
GKtmfAwxIMk1lhsrZ3q7SIJByVQP0hSg2KwT1ce8GRteAcaTFzMOafFY1xl/nRkta5XVdifNfrD3
iOtF71XSxDkOmkuOLidEglG7PERPfdyryf3uluImzOeVpJ041zgySZUTruMuq2K2RTSYUAfGSvQK
kDRRLzU8eXw5gt37U5QxMh5sDLVZScDD95baLjQeTLKZNKJziQNYWfUQ3DsRCNoUnCtTjwOiiQZz
tNbjFGNteyH4yO+1nZEoB6AY5UA4zFWp9LmPJtq0wde180qcK5capKMhid3XD+PKx7/lgbkjU3OI
O6ZohMFsLCLpatoWTptvVTFWQBBYAlHsnez2I00MasoH57F9IWJuT7QD+cTe+vdlD3oN1+QrRcB+
YZKqFbyFthSqRaj2yd9rBoy6Skx97a16FIjznTsYK+aVh4z+Qlq0XVg77DuyQ9xe2bDNJ1PEHOrw
tynTp588xwY6waEZm5yg014tktQxDGL6utzzDqyMxCydnmt2uw65ktX6nNtHb3JR3RJ+/DviBj96
mvudvE2bKa7byPjPupknJ1ZcNbNoa6uvPkcotTkGT0Z5yXdSdOSp4lqx49TQzUWvseltu+g+mJUL
rnBI9X0/Rpqomlpv2f+Gv+wN9Cn6U9d83PjlVEEzZxq1GmXYH/RXPmkjeaCLRCfsuofGeyvgl779
JhMG5cyIpFcsuVPurmwAs5jp7EuxD04w+70WWx/jOENkqo1sKjrR9gpHfxSpH73idYFuYnK0FwmW
6JOoPUM5kxxmwRRpRXLwQVkBFx6LnYgP4Ctv9884pazHbSdmuDloG+qgPv2JtHSHA/j36Xud3oDU
9vjf9wbehgXxWBJiIGR+007hNIAylGXsSJbzr+0/4Ahu1NszEZ33Z4OIc2Cw1q0aKhEOoUbvsgL5
kOUMwRMELn9t9Gjqkb9QuzYqblCoDlEGCvhgIFQqr58vBOlzktWp56Rodkl4VUosjtbI8phg4Kft
mNBDNG7lyVDIalIIvafiQbgObfxg7obqlHs9/kgBiTjhwIaxuJWH4+nmHmuZ3eSEK/qnmfE6fmQv
1D4Y2Z0tcFxY4rH0KCoGS2wN9JNYGchBxyNJrcegmnm0TojenJt3+OTC+3qj02Bxbr6HlKb2FkY0
ey7hROxx2dFHGsXvMlS6mvol5RBDJ/3PT0U767/xtf7Z6geXDt8I1FV+6fr+lUmqeLxwrgKwPxkB
Dx/n6S82lADLTebsFzpYsqVmzEJ01MfsHGcV8p/3uOqUeMLjRtBK/PfimZifxlfQXJjwynoptLWX
1Dqsjwd9P74G2FtLiZR2zl4woC4AJdAJV4QE8/eMBUb24hBuaTTTHvdcFKp6kj3pj9q9JZlLBVtm
bT1QhpnHkSlhHbMAZfF/MSYzzA+NqXXqxPe5nzo7f+mtpJrSHeGcDOWah6foS7y02Q0AeF01kvhS
LqS0HFkuE6d9Yp5ehhwUEPFvXz7Zw6zqGx9Zq3Qxu4AbPTjcMBou7/chQxA8zPsh9PYi1D+1jWQK
SgyR38jJ1Ws57OTrla50+t18luX+rtyT4ybWx+S8HBSWZBOOj/VvGgEw75qAdqvJm0oDObpHWa+G
YunreLByfBy01P0FlvlChoyzpZsyBzX+x1J7GlFwLdo7TemscOBZ6xeRiOFDqZ5Uqc7sss6BwL98
KzcBAY7uUsZgZ/fcTPv6TgDxrCzdD/ZGwAVAl8hHnh/3DXU9bEf1LXqSd/ZZFlb4qHv6t5jbMiw8
B3oZpSnZrZXVJkYHFzxFIKNkcP3imPwP7TeR8V/at4DoXt4zJQRpDLSvLbptVIxZX7SXEVaLFY0H
pf1WBL0TtWDkCxcrCmxnfu0VZ1paBEc1WZ4YACmsyCBWUOgUnRpu57JOQ2WddWfmang4VR+5uQmk
Oi64XU/Q/fFX2dBdWrrIX16FcbViGRpeCDoLF3A4EpkeC6kp/khABZ5iVeo5eC/wNAoCVNjS3FPx
4yqJZ8g9ypCBk0x7Y0Y5yAAFg95w2LXRsc1YzPdd9ImlAzOcf1puP/p+KDHh3Hyf6hcEYy4JY9bl
HGMqCgYPbhhEfbD2RiYhk/luWBCBtbDPXUGs3+xi+954tYCT1Hu1tJUgcet1gJXE3LG5aMTJmcfl
0GGiKXie3mf4GHysNTKNiQLTV388JZ6cr3JDwM8IBCTZ34s5a3m/S8SxJzkM6NvoofAObsPsjKOV
xUfYuCb5yKzyghJEy4v6BAG6co5ptoqN3V9lOqMSVcH6xdH03wJiaukm56VVCvCkB4ow1og2+uVQ
heJfWfB4mb4kPxlljGH3PvPVRMjze3yuRZp2kHGOKzJx9N4oG7qSOduF1kVsv4VhCZluVb1PEY5R
tVhHyYLlDVIev5v4byX+n6Nf0x8SVdaaH5XLF4Y2d7XwKBak4y3SFKIvmjla6cha3VudRNFAhUNV
RWsr3SaVAZXnUODBLxGIhk3z6JrLtSMaIxJURAm8fx2deZmPRmAiBWQRIgErE1rayHq6rwtTJNyZ
tBw01jW1GTYwmOELr23pgWrPuM0zSjq3oL4Q7710fBoHFZhqj5JOs0iam9xzK0BMJo+T+Y4t2g6h
IpL8r8I8XmGtVPflZ+eFDofxVEqkdUv/HXFzxY128df8jzy9qObX9EYb26F6nutF88fUg6pfYI8a
5ndEOWPJgg3MCfnebtAmXIVfaNEXenCCTs0Vnaf4HXFNbrufWIX6rgIZg5UBMjbjHXQDxjEG5PNX
nbVNVGR+SLNLuOCYtat1a2EVDmnexvuoCcgB6VmGJvS8FGxmY9Mb+LU6SJrXUHvM//p9Gn8vLrfq
eJ5lWnfz9uziTpLaqEhHELQC081cqj7LWfe9VBONi2qQ6Pki2BpcRlbqm3Fyo1gNidp5QKRFm0sM
M/NRnBjumW0w4U2e6x4nRQktWkRvllIFdGtHMgbMK+0+KCYGFIGmqqJOMV+fIH/henqGcAfEBwwq
fT0kV3SoLdli+mxvbyv5Am9sV4f1t/0k8/o5LbOVODRw0+M59DXWnXJZo6YGzFLaCLjwam2CFb2U
30ODqysgHyHoRXCS1UCGtxPx4AEVsdgwB2q4qxyUI6FdXLAfYF4bYsSn7gnmuTo7XpUBIXmdG0Mn
htwkUHEymtvlFc4Gs7JQDrCc8ZFfTsR1wczF8hACm701HzOwBDUWlteS7Ce9P+HjSpUnMtsk1Wus
LpmmEw4fL3ZKQug1B038mc+9JnUOj7B3wZ5pPr37zM2IrVnJ7AaUw5KeHjNt6kEFXDudFuyz/NgN
9Rqjg/GIaifxBmMS0NRSdVO8rvj+5XBxs3NIktG0eaDWi27lvGelHRVcqwGpH+Suw+xbilxQBvyY
jEN6Os1pZ8TsAbpYDdeiuPs85sJ8cCaNtJu8XSz+GpBSa74J6rHJklBT5Hxs3UkHeSAZ1Ks/clrx
Wq7shDqaOeWgJ3tnnw27v0SgIorCv2O5pyZAl6q/pfFfvUHIc3LKNuecPe/dpkOl88nRBUAtJQnN
oMvgkn47Fi+EOShNY1WBqoFEHrY3YLbLLBqJGoHBWnHXc53J/E1OXVtIOeDEkjKAwj/joOjWHRG8
IxEKLYRM0gHiBVZE288ITfox62znJ2vbFQXVOCkEogRfonKchlgw+98qdRG3kbob0MwqcaXQq1pr
pSYDSdmVJwg+tWTJcmmfhz3Pt8/hj0q/Cs/y2SUYQGUmC8yl1LBdnVhWHafJ483/vgxR8S+BGKtb
uGnyF3rFDj6DxvdWQMBB66q6gxLuJOUft5S4d6ZdW7lvGQteUW/juvTLAFBvLD3475Sf9yr+xP7A
Wv+qRaAHs+v50pR+rKeP0J+cRpbrYjbuRlQtIHOPJoo9aJLIM8mSxPVxdQwWz4VrqxdLzs2rVmAf
LBrGPMO8E427fLluDt0R1oD5fX1uq/uT/ZIoFoiw63sRvQzbg1MXVT1GIbDmABF40Yz9YyQUjSIU
z16582/wCPMpren0ud6NSz7Vq75A/h2y0kro13D3h5Llg6qusT7ItvKJs+vNQ1r7Glda/Lsu5kkQ
Ap6qRmjSmJxnQO7RlN/T4OOs5Fitol/NgFgsh6AP/ANrSw0xVd3BFb4/yHsQSxWMQH+i1aXCZb/x
tdfmV+ccAkvOclKSDhKnFv5LHXWoGR5/9wZ94CpNZ9yY54oPKuz6y9RScamKvaG08kAnKdvfFFug
3M2pp4m0G4TK/buYNDj7uXyYCYObLT7TziPxIZeClX51PHVv6lXk0+Zo8OPMD6unQQA7WWC5oF3R
X1kdmfZhb0bnZu+oZ8RMzU0FWLbfDc9W5+OedvQ/o3SzrFI6LrnnovFSaFFgf6yQhwEPo5WqgK2t
xRz/JsytH33CL606rQAk61/9zMtLaX451dLZqFtQ51kMJa9K5/lg8/1K58tmjbFCKV4EReyW/GvR
7v47u6aWypljP6A/Z5uKHqQDfJQ6FW2IDpUXO8jMLBfFAyTaiU0T2Qqny+MHbTi/kVNeKHgtU/kQ
MgLTCdYgclhWa15gF9qz3/SO8/7iHTIUv9tGZkclWgJ4UMeHk2j76ovYbBU3qn/vxX6zKfGM+VlE
POyyKy6lK8tmxKYyal5i/5EASQfqujr9eoehVt7fonQZTFPdDkI0f+W78hqyjSlWzW0+t4ZjIlD6
qvqb/LLIUb+Qm7s2ukQmjVygRlKfZMAuuFex66U2OXbli0ZByDEST14Trbk7S48Qu/Go6msfuqB8
SwmNH2RlKrkCgkblIVW1tuHsHrQfebN5nGb3XL2SswIFLts0h+wCz8fkx5Zv0iWvTY4XS98wwK6O
9aCa9yUGz1VFZ3dIPoVOsV9REx1hHIreQjseLUMrAhWU0qq/q6xt1w5HpAMyB+9PbK8vbyuRLQmy
KSOiJS9a1283ft//I59yBQFOWD9m8J4QP3vlbYr/fi5fGgDDsLejLkG3uW/aoY81XkaXJMeFDbnP
9hsd7xmHM3RhZPthFkPpSG9rzTwz1YdtycjezUKxaM9Xa92SfCIG/1DX7R5VIhCqnnaiyGjgxfUL
vgNAB533Lxk9eMfP+PV/S1wtasgtsvgr2DfsmB/P0YTOqy24iJGclgIcM2upGk+BCtXzXreFjMLN
s1Qpa1wrGo1KYL6AzUPUFhH+OMsQgLR/J8g0+nrfMVRNr0kQUbDNHa4y/oIM6RhXNPrkQQpn4Q9e
IhFiJtJXFmRQek/PU2aksji5WsmFOHrkock961OndnWEkOCTfCzOMRqtjtVNGHej9d8U1IgQBju7
RO0oJ/w+uweHiMeYSkbvXj7KMsW3dvJr1AVOJ0L4wwA2Qb+LXS+WmykS90E3H2LM8KX57L0N59Nx
IM86wyJ4h1WVVQCFcLrlrcfxT+O/c2GVf0FZeX7SRrM0/3CF1Q33QIw3qTOycUJfW92Gbfr/uSNO
4DM6VUM/yYq30QJhcQCRTGmp11XuEU8+ufY8FBsKQCKo2/Vl1URugzHyTvxAwHZyQ0pXQrdl3jsh
rmGTzgRz4hyIiSP6lAC+WHSX8mOn/i8D4LbCvXjbCwekq0PZdlpJHn/nzS7qjWXmQmPagajGfsOn
MzM4THM+085nikYsnBZACPzW8/rjhSx6XSYJRzpGXXupB6A5PTcz6mR0HbzwSRpNHheQEdl10KbQ
qN9jBs++30xcFWvmH97qtboXgFf9g9qjTFWVR9K2g+Jg+gfOxGiaV3Xj+PpKiCpEPE8dUU9EjYTI
yAur4tNddobkK0zFEQAIohvSM6ZeIixWh27XuqA/XsM3SecaUH9m+BQQ9BT7hDl0p8NGve2l0jbG
80QnEf/ApFmqj9TttVHv6rU+3wRuVgKNuP9KW6W7RXRnI8gWQETnic+/PeLoE2vLG1S0oIKeqK2K
yatibWusEPnp0ENUj8jF7ST8SVEGQ0aL6VpymrchuTLc0mCVGA4/oHfPdzgyOQHZWksfKWy9qNoM
huSM1CVI4CuGB0VpVmY1Xpl3IRcno0D7ZeOWBPmmNlkY/lBXosiVot5M7DcYpUpn8zmTptgG9yvH
34SHZJApFmIlVSCcYWRzFZ/UV9mg7818ovdJYKf+1Fv5i12DfdmVgsDDZoFNLf7EOWv3UG6xTp0O
uFl1gb4GuZ1gkhPXgLVuy/QzN9xEHoWjnVrRAwsWwDaLjB4tsvnzuRRJ7Bp9XqCebs78L1lNOmDk
obuQNb6Rlord8aeV3AU7cd1ITcUsrQK94V7faUmD8RPpPufwFSg9ef2hE9uxmRORtxeAmyVB9iUq
u3fty+/CoRT2KsIJmE4qC/Wwtl0KGjjPpmLcVusEkjJ53sGHPsy6cnBL8dUrjk73HfE63VkOEAAc
jvtasW61o0Myrgzrjr9QREk0I1lYsDbOjuvo7cWdNitRksIdewXcmn/X+EFI3WwSrvoS/A/YKcKP
BNRE6un70MAF5RZK7WTELHHzV6s/R58pOsHSiZtPS585zUh4f3+7GZhnGBuB9neZGqH4sn04ep9l
5goOL7GpJOTIsfRS69DdhKkQBRgchNtrsFlagYXyHckTPZgYqf0StC3rKYbRh1vp0n5d5c5Egk0r
qWPc2QrlI/lV1+MFHsIjxDqCzmQwkN/PhHv2+zESktQIVjZ4o2IwTz5bHHwbH819e5LFaDLhi8Nk
sTjKlZ9kavvM+fddhUUJbssjkS5M8LoOq9jdbVQ9EFLKe++vjodz2HO3G1lQ6ilDoLWVGpzLM14P
oEb2ctJ1OIqFF40DcYJbP6kygnX6ioCxE1QvAuixXsflasi3NzKB8s9fagoC9+B4s/l3VOYssJym
DPaJoLNSZ4fSwos12bMBezryfLPgKNRLR0hEHwDfrbFMf+khSMaWbWAd7FZkxearMgZg6wcAf4F6
NVjLFVRWhObVRVzoA9KOlsIaf9ib3l1P2+fDBXKPr0HZMqUuXLpd0Y8EdjQLhZ62NKUjutgt5dpl
pNF/E14Ra7ZfzKidbQeFIvhcztHgkF1wW35I0JhXCN0yXE7GaY+TGBefFg+hP5wwHgqUkYe+fuzu
aL4hgScIlXc85tiSKqGf9s3Xz6VGUl+CzkuZ7KQKBHdS0z92MWYXmkh6LE3t8CXVybbxlUw8U7uB
tXJt1I4R/H+421s52JSWFBrB5PAADrC4LKjvB8JjEBWzi5wbPIHNgQ0w0ehZUcB6ZpNdLa57YvfV
ssFhIC+e1aCsxyD6a4hJRSZAyGk1EfdtPYX3tHgw6QvFsDoRmj/EVE+ZmicvVSKVvf/agpGmT2ia
gpcyGDf25c99/W8pJpFaYJjcnTEMcVTVEYUIaQEzA8Ap3Hgaz/H+OQJ1ViG6LUR1kEQ5+9PmOWLY
L64j6QLhhsEptp4A2bxH09hZ9rllG1OniApWrv53MWvRcihJ1Xr12KFIIB5QEzOEhwKEkigDDUE3
utkwlhIrUeABHvwmYrhJLIlzlgkhfrj4gknI8H5MG1K7RRe6OE3hrKs1cEgLRZdp3aULTfv+jD37
lK2Qus0uDGfcbyrA8uSR35oHI5XPXK7ydUjQDdWRGBzJHk4cGaJRgtMTiNkMN/jFKf0UTKc2TVrx
8nyNF1Irbcxljdjad9BoAjbAJwCtRkwYf+DZEPrAy/02h6A4TC1zJ0r8qPbS5CfrOox8Tj+XzcCC
vuHwldSP4eN0rfjXgOg2GkDEjMoMdsR1YqhXfc4wykb/MR/BiCWzVPUfAF/0B9ey32za593ADkG2
8tLRK2HHQUMHhIK3LVp380SNMKaegRnC5/QFceRFFyDJWjoszjWLFHR3Uj7ro8a+nNPGX94DcpZU
OpRTfQJjFmUb6VSZxe2lCgebfh1avQ2LlbGyjoZmcrGiolokf7+zxolLYF+h7YgxpE5D3RYs9gom
c6skYGLPCPJLeF64K41DXkk1VtPlAnOR2w9vCnrF69sAfdvu4frThrl6es/tG/TNSeXDnPRP/tkW
BdLXIJ3T+V61MGryn15SFYgj7iv17pkypxImOgZK+tsXQMLPIiAT9i6WQGXoXuNyNFaVrfKGfUKp
QNB7kmhr5Y/dz5AcZauO9c6hTLG48HDU7isNz926w5wvBCaTotzj6d6rD0yaNplsGM6CUFM3bwB8
9zzLaUO/MPgf3Vijtam6TkzpYQyaHfCGynQ90NIj3uHljEoHoa2Z+zJTLK6ezr3k/LUmJ7D11Ii8
jefhNWWYargZg1iXJhwLedYMvzzvvq1brQWDPccDpCC09rYIiAwpnB/zywG4PKOmwPfR5sU5p07X
aM8sG+OJcXrDETUDiB7d7CLm19uPrzgARi0bFxRGQuQfdJ/bTFwiK2JKQ3hdu56mB0WChwjU8Xyd
IGaGXEeoeprUlsXnhv80IPnZtreMRT9oMSvC79uPo+bNAMgbblfhyoFV9KwWZG+xV9zGqd98fFVe
ImFXwND4EuqC/dztc/k4GOUUNFHvmy1oDavpG3W+qt0EczJJVuaBtiaJlfWYfPkRx8iOFz5em5vt
FG1PYx66AUAmUBbGWSUFQloZm4UnQhorxlIGcjggMRSytntfJU2m4QtnsQ6E868kZB8O4N/NPkKV
dKBWe+6aj2zHI3z9hqe1p9iqohSKLcoiBIw2r/tkPSG21xDRpU3c5Dw7xFP0adtEwvGjSuB/eSgf
TTj8L54bH980BOHbUnmKU2X9jRC9E1a+hui+t71xEUFfrd95S/wK43wkOKZqt1yNQEI9s9gz1qeV
+H8I4uP8FXfMny6PxZlo5MN7DNR86gKncVa7hla+PrTB25g2jkU/r5+hh1973FThQNfhVS2QedrM
sR+niz4OZUa8FjlgYCwsaJrWrmQlAWD+hoquwdVj/WAKsOOTq9STbgpwLpsHKJRIp74YBg1U9Eg0
eNCdYCPBmfLxCyQglhmxiiwV4R9xw2i0WKQk2pkg/u7ycQftMxMJLadEVtYJtNtSbyXaDbI62cXG
nGvpb9iBliD9IKYX8WjhPA1liprEYpky9/m9rr73VO8bwtNfgq9pPd/4tBaGfKFUe6Lu6zv5adn5
aqgsM4aY3KJofOkTwBozMHR2RFbuQPt8C1g1LJzwZ+K++Jg6ZF9YKRPMc+UZYnsQB8t49sJehUXX
Kmue7ekMyg2hMnKElT00prD+FtYltDLwEEQdhpKK+YZetqyHAvxPxKIwiKtWKYSZgwHksbR45oHg
YUS64gzqzn+s5kPRJ1wOc3Z/WK2UCwV9R8nev8Z6v0Furah6IEiZYp2Q5Mi4sWLHCqELCUrea2hF
2OEyunTqIM2OqYfyvkvWB/ebJHcDAsdUTqzVNqNM4G2FY4/AviYesF2jrBBMuYu9IyociSIa7mYh
gHktbxPWb+aN/rQFBQfS1+ZNDz9kchlo4vkfP81TY2jCGlTag1p0fBSHJxF19x2nsbkFHq/MadXp
vuJPxm1FmbMfdRTwJ9/33jKkjYe2t5PmwmqYM7Gb8qCc6r5hQmPIzXW+VmzWJQmxpjw+Ro2r2ifz
Wd9+bs3Xo4ejUk/8UlT+ru7o9lmXHlNDZCo4AK/oeG+3qI4Thr0w9G3XYgflJgm/cj3rp/eGwn6O
pz124Ij3UVjJcnaPZJlXOGJ/ZvIkvRgPTmL542z6/GSWJlEwqrskapOrxOajkTT4E2VkmOZoJlKJ
ySCInJq7W3fWY7bt4hnhJxwGj4zpx+becLAj1OJZJ/PSl1OJBqCt4FMQQlBvMKEIBQA66LlK8s0a
o2cYQIUZRpz9L3LymyoZ1sM9Rb2of+zIqHwpcy4EG6qsR/DTwSpXKBbedzYYQFEzlpW2Hsg3SdEG
18PBeiqnUZly5HiBi0QxCejwwhdeWfILu0Nrv4ReRtnYzE8pJv/N9ySPMmtqOUEoUZsRqfthA5cE
5pGzEAdh7y09QZTg4D74tPHf+4dP2W5+EKmgMedDOTZK5j/TE8Ur4TruwqGkZsOgi+qfldsW//oa
zhI7wNHe0ciYl70lrekczCroO6es2iDRd37OKI9KppMETI2lCJ0K6nvnxALBG/djn3ZXbV4Z0gQm
vLrxABzTKeJPH6oIQ6ctHQvlK9k3MsNnfyGFmKS34U1EwBWjHWAn/AXdY1tVHXbrs3eBM4b4GsTp
8V8qAkrPPgYks3LaCteca3CtKKqugasvePx/5kMAkpy9mXJwpGR46+4XewueRRQVx3Rv5gcQWjO/
tF9JoBtXg6fqr7yEBrBSYbrDdr1dBUGf35WXcyGGpalYFF3pjcZtPF+5xANytpd7IVJ6E4PkMbZL
uzwvMd1bBzzXqp2ygDfK8J13orJFn1dxHKf5tYpV42etdmaSRFxBy3ciemQkqL7JsP7FlDBkgin5
Q5k4+1Hrrk3/oPnKZ3p5r9aVdR+KS9SUxujoC5o/WeUAx8QZtaV6388Hxxoyt4nmgLawJipkrNa4
FJiYYCMgwa4v3HCBuxcATDOAPee0vD+JEOliwodHsQ0DsiF8oJMZ/9t5V3d2r3NP4vx2LsCOUTcH
67TCGqVBIQ1E7RZEOUbt+mYCntgjOLfkADq9eM2FsIRzsOOcFdDLy20rW/jtzZZp5Bi8dA5ZNFyF
h9I0sQKeAwSId2WGSj7TPaKvgMHeopPMcQxpg8uTZr68lq8a+K4Paa/77pZQiWI0HC4EDIj/g03a
9Oozstfu+74octcmH6AUT5kKnckl0ZvXPPcItL7azLN0ctV+cPuJkMW5PUUfvhPMQwnBeoSlJlwV
RpHlvPhohiil71XVTlN1MPAJ5JRCxyPFXU0RfbITs2hGeOFDbtzhu7USzl5uACaoMwyOi8Asht5B
M+s3rBaRWEywucppCkwAKFoPGMzMZxdT0snQmcNtpREXyjg5qeLcWLlSF5ugAiDZZKfaU99fLrZ5
/vcDwE+E1/+BH2mjPbsMhzeBH1Nhso4pzPgl9g6y3zodaPIS0YbiD2BPUC7VbNUhYugEae0tiiUX
mv/V56J8VBWQtiBJckMfmWqffdTn6RfVkoyHGEZTFK8saYw1q0705LpoqagEgpbgx67N5pte1uQs
/6Tl9m/VV9TSIyhJ+vB0i4P9iW3au6mZniCkhuJKV7x5+jiLbLKwn/kkkTLy9oWul10lglJVpI2H
Hvxe+qPTWZGWUy2vh5tkLFcwPcXqrhkOV5ReQuzOqGsoBKt2OkHYTybRpLoffvS3BWyS0HMvUGD/
r7fcwHqqIHJ9b63L/A0OWSztlxUIx2hoLHtorowMgTDcyJ85k7hT0osGY6oaoC7G00IpLpAF0ESi
S8ZZ5ammZLA+Q6+I8vbqqJ2IcJj+qbHWl0FgpovblsP9TmRQM9hUD1kjvxzLevX++B8O/OUIffGT
cLAtt64hrWO7jWQmxgppHxSHXqqrqb5IkgxsAup1QcqAoWN4fWaAlNub+3LXFDoVCgIuhjgfqH1X
W22yBOL2zVf5VKQgnRZlyr5Ovf3lGLhLgt+nVlXkFXgsCNw6/Jt1v7PnhmRHCv3RkxDgIFGMOiUj
5RqW5KEFNRxdA4VWeqQlmfSi41GuW2RvqBRxzVXshUYgN/jOurs60LuyBn+PcFrwF+98TrJKP5At
P0IugVhEjo38/e70eLcRZ8tojWUVU556XgNf6FFFp6MUUtl5kPPMzL/ZDkZEMFsEFLcMWk/3msi0
qb58ZQ786SPnPljjKQczPMjDsu8UWalIhek5GpCCs/TrfjDjsxoHWVn0ZKRqbiVk8/GUWkUcespS
big84q5f9oCNWWt5fa2rUy8bUJ9NRi+VXohG6DaPmHcYhkeuYokPEEWp9fTPpn7BJWYsMbFLF3jn
Gj1JbeRj5Z+7Ene5bdqRdikRUAl7hsxyYycGyrxXP7d2/xuSWSyOYsw27W+wo0+YkWq8PFN7u3bz
hnz4Nh29mTruQSh17xwMYmXiinDCINKCzrpfUYf7isyG+p1n8pzKptHAYf+1ntdXyDNfcEY33ckx
AYjOC/SxdDTPVGhCHbnDeWNFdjLXz4iLkcuTgqx1OkAF+Iege27KYkqKYHPAN4pzmb+TFpfdqiX8
WLeAhojYJNDAGfjSybHbCF9UWM/+EAcjnWOw9qBmTXLACNLTgLVkKroad3uQ1q+pL8QD827JFpLV
Hmv/bUOrULC5NCzQWcH8gARnBu3kzO3f965uTiVbvRbskS8Qh1vEMr4KEZYMkPEfmYTSp5nx/jzM
7ud8IfGPNVplyjhVPG71otMw7X+Yzy8ffDb2cWqTvCcHEC7JlAq0SSXrgwcYoVJ24x12ImPv00Gv
5ardP5oh8ktclbAc4K1FUDuganqdCw03/qhDYwbyABQdZ10uNSRv9VxSbws/E2gcGA6c4TLGn4jz
2vdJpx9YjwfI4wu41ovbvei3d6rula6A/iovzIWfTubfyWycZsFm5D0juYQqy8PPT7Es4CxFxeLo
XCRpQBRvfXelgtQAlmnx/dTYpeF6ulYiYYROJZXEjP2Pr+hE20aQK8Mtd1CIFYzbZdFzL59NbQik
GEaIxSzswf9DL4YjNSvDXANgYYOVozrMRvLJVD/tFbJUI3573OBdEYrgDGrxbacF/DGDH5AcM1B+
7XrN2slA+vOa7dJTf9QPqId5EJtdnEGlwe9fA4zfYtoj/lW69resaInQaa8jvMgYg9rWE25JS8bv
zcf1S4PGF6rGrPe5+Xtpb1pwSoN3FkPjqK9Y6VbhKqG94chHrOlCr0tHrNq6mtR/ntJsjm7RpQ+6
UVh8Z345lflZ7/0cYz2v2qb7rx18A63xxKyLRfbGb20XZycBMq1RW7jBlVgiCLyGPz8DVWii04yG
eeyiqvoaHdwMhwb5I3WmZSKgg9iXxhawJaNbFnCJ+OLrFMpQSDayPaM/NleRkxgojfpNjsQGAxgJ
kVDcVWb9h0NSfPPyzbKIcjypHOuOXTek21KL+78kqMZwR+rXCMe58fFGvJrqr94Bp375Is0UcKlo
r2CwKrH1Xfh7vFksLl9utB0vo5uDNbkK1TFHI4xdxnGwS6vxZqJFVU4TcrNmabZNg7xKbNoOGHu7
VbxLKZPX9KJofB3EmloeI/qY2UmTNcLePZKV07dCO+QYI3LZ+067mxrLCMcKt9S2oTvmUAQ4mZH1
jHM4bEYDmMPUDRHJ4FgZynBvBQYP/LkCOnCzZjsZOFdBTC0VeIha6eYASwYlZi5o3TN9+jvTJ7dX
AALsn6qqjAMDV0TpVbTxVWS33NalE+NRBUyfAyMyef989EpXtXizLcjrXyzh9wD35KOhZkTRhJ0E
iqJVvAyXIb7l0+YzmHN7c+KuGgvBY7OctIBi1E6uCGHcFBIXR5IsP/8smnIKglmhqsd3AELJO1uz
pneyC0qZ8mJeYEZPzrZx2wwjvCUFxlwjRGsMbuVF4Z1ypmS1jHZFZFLl0L5ZPGjE0h8f0LVdC36j
rq8vEascc5kOcsAQUdq9VOlsEy+Rgi8epVJikQxVycpCsxIWS9VzUkP3jdJaIXcv+xzsKmnBMoSX
Rm6JyHGEy5vRCuAP4pR939g5Bo+vRt6p0GbZC/+aF002IdNvkAjwmVLpmoeuec0CNeaO20hrz2nX
DV7Thryq/Y/D/hXTbqzM7s54RW9ZMtDaVePm3h88UnvyBo2sju3h0otLeaU3I51ZpHr92uhLWf50
dvXJAlVXN+MyLRZeg8o4Wcq5yCRNNhKVDutWM2YY++eau1JyTBJriEzP1zYcymt4NOncMco1n9cy
NvzDwdpr8ju9OhMRLydF2Q2M+mumMHGt187Pre6EHm7wfiZBSsu2Ve281PkR6ogpG9ptrb1vIgpL
zh+BaCC+YFIG8DAmdAFWsAeTCtfWA75WksLfT/vySNlEY1sAO9edGsboJoC7UagThcaOkdhmrSsa
Z0Yg3cNE4sbPhS3qWjon5PVoxM9x7PJZp+3/U74rPAPe4X0e60PoXqsnxoVQ4PAL16sSliKU3lBh
gFSljwaDZxqlrPHtlmsfuPaNk6VTjQDtH3VDpnpQvUErM0DlWdqjc849YytB3LMTGJBUoz7zqwmZ
4+I58E32mlPo8UEHaKpoWtE7BCftQWuvPQpcHNnuDCmkr5w86sykAD9uSlPizXTf6n8OshgbKlqQ
QBoxBGZjs2x5nW9iydUN7511DuWHP4LxpS5DQQq1/XtQvU4GrY4J8AyUeRBZPSowJnFMRVBOMYRl
ay/wpl/QvrUsFSSuhaUwFVp+2j7Qg50z2cVTGiZr9gnEN2H2DEXSVwiyOzan6X5UB+K4140hGVqj
R1d1enpK2cHkRR4OHe9iRq26Eaw7uU2RZQyOfE8MyTgBhdWT+SrrXwhm8v6SRFJaM7zFLezixBXm
K89uOlvDzYlCsQZ9p8ayvtvGw/RZ9Q0NVVpYttB2Ombyi9JpTShew4AqM0VoDfz/8ZF6MrQZsNcY
P10MILnL3Gu7VJehgoUn8vC7o1M3ns2lqgj9oC1JvlNCMfYZx9mIBTAHb1JLZVpaRl3429cEHmnW
uSzP63adquu2L19x2y9/4wjYZC0g+ejBsdn+KSnnr+e+oLdck2dDnr3QfAtNv8++A9/WGmyFJpX3
mEeXCUspdXOfbnXeP1ZJQQuTF0dkqgmo8uED9wl7kwL5IHsuLJD/5ZyISzF+VRVrOSeqwbLmJonp
KnZiuasuFSUoyuiJuFqkAcUf18eNX8iNHl1/T2gNDt8mDRUvmKXyDd8ztTF3uT9/l6e21Jf+AS2i
2wrQR48HEF+f0f0wMSxYxR4ugLLrMm5igRY3+iJnl4Wi4qrunswOL6qwSF35wnEwvVWTP+krvys5
UHavWTmpYkAW+yyXtIx3bWQCjwJRGrsA2XLCq59I60Y4ichdbVzjTaGtdJU9+zOpHoOq8JrQKAII
wBs3rWc/3HHfrE/sWkoB6oh5z6JXCmI8zqkT05MLWtnxaW3j3XVKM7znRNU7EeWiZKHMbJLvnuqw
pISYJFUZfeCwZhUd9CZcOtAy9+w/Z8H/TcNZ8kj7RRhLQ8AZYpmNEFdswaJq591bKhcU+hy0Eqe0
cxMwE7VVw7Kv9R72vaocSxFHcYnBTjj6F90K55QD48sspuFRyXOJCn2G/CAb8LScIdVMyztkdlcS
pIeODO3F3Cj8Wa/+DPdeyBdW4AV7msEXPuTxndQpohXK27puen+akjn1XPYAq5I922s3wRhwHqFk
w8rD+vyAEjZTRIb5ATMSIFydFCjGrObuMAvDCGNHvk5wq49rRj5XlxoTZLHEH79PjcpohFX03pEb
fwpcdZDzRb/wcY+qY58dnmngbHa1M8Jr1Ssc1fxm6lPCaXGl350Z+G7ZZ1235bnJ45fvhiFterwG
a5IQ2l/jKXVRauMTx4aJXZL5rrlBRpW0UtfGs1bZFEDxDakdRt3ULbt+JNhkOM4d/g0BzHAaK2Tw
ZU9IZGRlKp5tpQVquFC75knlBxNi28NNVBQo2Ep7fp5ggimLMAO3GzOq5P3zKy2qpIfR93pTq5++
kTgGXabktQmUQH2cC55eVG3/KJjmOmvTnc0vLfeKBrqWAbC3nFrE7OULq8as+GJO/mjdofBos+yF
ctcL3vAE3/qmyAdZk6VOfjYrQf11vKJ7mG3Fdsb6tGh4U2jgHWUvCTcS+gj3yUAH1QG2ppV/C3LK
uiSB+7ij1nF6l5d2JI5V4OiwdRkmEO1VmivvG/g7dHUDZ7il3yOX6NkK3NYlVSM8cndQ8PUdW6b+
kQ6pqsidLZ6tKoyUxz1ggOxooAm5tbAw98fgL8lBhSpVR4c2zFN318v3LUG5exk42yXUvlWcNCog
+1adQUx/SlaJgZGcAB5MkHmYIUFVKjpbg7wleA2P3Z7fTYL5ltRoHFVZ9BQYbBHdSeeta/QqW6rm
jlatm4z2J1if+ftLd5RgpzpoU+csqse1tCeFvNE/ye2S2W7hxbwfqZUiUY4YcNwtUzW8gUCQSFWF
JVU5fvkm7ITBDCvk8ggrgTZzGyMxYfrQhY4yvVOC80nyBn1zjsneP4NK+KfXKaqsgTLFEmXIH6SC
RVUgG2yQ95T2VicZcFMokW4N9rtxYHYJPPnXnuo0wQJBH/81Fwj/Q/Y3GTa/5RDFdRpARqXcdxy6
DKhY5NEblgo2jjJW7oFkajThySRFgiUihtH/vzIqr6xQZazonVMO+659bZmqaJWEHjPHU3mgZoyH
AMvIphTcx9nT6msJQYMyYXlkr5u8zDKJOpfJ7BV1DRbNyZWfMW0XnPYewe29mONarJiwOoTqT/2g
Xt1l7RNP7C3DYMEAQ4+6SDkNJfTFBnu8tJLJ63StPhaC/7m4EMcBlkw1YjqDsRsVAxV2LAhruLPM
PFaY2hnCDshu9HXcHgAIBlLSOHpGlt/7YuiLDtNjpkIdz/DoW0tTnN69JWmP9iS92zzMKU1WCLiC
VAPMjz6Xe1ndFtSsMFRMKM43U6+XdSEj0/1jpUsKYhHU8zr8OfCxxUbdo1YeRrmiIGCDC4UuZ8li
3Rd97u55DLs6c09L8iu7IPKC14iN8PfTD0U+8+pUnlwYd9YMU69VNT91Tt0oWSnpNeOBa4jHTY+A
yE62Hfz6Ib6z41iGYhVvTNMS8AfM7LThAk6/AKak+zByQkHZSSdxP2FueZ1w8/6KK+PRmYQOcmeT
gQitZr8vYuMvSmpGYlbvPjpoohUCSwoXuRYRbYdCAEfg6CnFPRCSRGWLr86oes6AjIl05kLJTUvt
T+zx1ScXTgR9/LZtgETJuLwwYVKR65EPDxB9W+h/IH7IsrAKb07NmtAKAk+md6korHIvdJQuuJBZ
yoAl0JDTFDXRlEGIPJPvfLn/pj7WEPvFdtZRIR69yjpdjr6Dm+/UY64d5dYV405rOicIA7BYrkCP
gatfXLTXPuIIsQ4vag0lVSXUCrEcd2n903cVZ28YkCqKAYWlXPALfrL7do0CTo1hwcletiChV1Ju
pX2wzrLCFTHxNl73lLLyBbzsP7XXyJcbnJf+5i8oyi/q5BVXhhNXSKHS3o5KRMYKpWbROWD4IzlV
CK2gvZuhm/9f/rSp2S6nz0RB4GK39KxUj0WC2X2MR4Z50wnamVZW3vQq+hc11CVPAWlldY52f9MT
bdYXdn+iDNLciKgKOWP9s3f0R2Tru1b/MJAQ0+lsIterpoF2duyo8/F+rlH/f6IcXH3Wlh/aK3o1
IqtRV/il+0HM2tmCec7HcvxgP6rdbW3N77ptmwSJg0Ih4cxM3SpvKaSKeRn9rpiugMH7Z5aJ9fUD
ofcdHp3+BDX6gLyor73dpjXXA2vQ2irww/PiNvB/ORZcmMYXgfd0+6JQ/UhdbG8r1S8s8lsQdGr+
d7O5E1s32qxYBFSFPaKLylHIDJXqtkEGB9uaTWhinYOn9nm2JVvUlXwG5cMZwsw6W4x1IpN3pgoZ
L9P5ERdiYrwN/7Bl9c1FZKqxxYutD1ayzqBRnJkJg/iX+tIz6xV/eTsN8J+HfYfbAXZMDpAAhXFE
IUVXc5svIud7adEvJh5/jCtz5tlGqthPy6V+eUCLZaV6QEWXr3jouTAQ5h4fX91ougqSMbdJxiIR
yYIJk2EVK74GRrd64cBupanWxtM4MKdmRF78MYGv48oedn472huU8TK22vdlifdOPzYxIwsFG0Pn
KqmzyMZZMhscQJYiW+HBlMJwPCyJMiOXCnCmUSvAbv7c00YfQ1uM8V9y/TBjWWxJEyiJLRfgpY89
x9gpYTSTptzUUtuuE7OTz2EYDitqvzYGCssVs37P+fp28LhKFiyydxa42Njwg0lMqCK0F42RnT2Y
AjqRAmz+hmo35NSwmvuJomQODulXK/65XxXIeZrfEqW5ABqYOhoUp5HMxVzdrTXvluy3NDs+0EAx
Y78apyMi9ciIufCKqCLA/Ykkio04zcBWJ84Mkq4gxUhDE7XvYiuCtSf/RNMnx+qbBNrYX/EZbW7G
6TLPcdjkCNTvb1MYLAAixIgbRzMdHimIPQQuppqumZia6wFFwOX1fXhmVjEC528LO4MpIDCaO1Kk
ykxp8ot8BcsHMR3ECVegdkdnvbVAhj4dguydZv+HdwIcP1kmi/vXS0LU+/onMCHmIFdqWNQKcZ9b
lKE6nU09h6wVaYJms/5qaLpHWbdTAOY2KyDBWjDfAn86ZIi/u4kwGCZ1xtr3/vi+jLCIF6T99zR0
/k0PgNZUSUdtVtqk1pdjHpnOL6W/WrpCHeXQcO+kAHDjtAEmquwyMDFiBLNn3VaWgsqM94Iks18c
4ABujjRDbzW0s2NPjI06XkWOuVzwLUC/G/EBaEHtC2RFcWJSfgsvdlJp0FFhYbuNCGZy7yEWiX93
IF/5FhG+GbdJpTVv5kVKLorWwwKC0626AnjEWTSJb0Thfsyo1FNDUDDh+wfPQkyMcK4rlOUfLsLA
Joe0F9jGiHzG7X9UY4V7ThUXOcdd/z3ZuJP9LvvImIti/VL7ouPEcR4kA97MZ2eMhadkivzd0tbT
NQqUpC7ryNRf92pN6VyElbA9pw408b1fZBF6Tajv8NykBhXtFZg9p3tc/ZLA9sh6hgoxH9c2ZahW
ef5Lvuh+V7ss65YZLjDZqJeMrxMtO24V5rIJoWxtIBpiM8/SmQR+PJX+uM4W7GXOMdJxmV0miyeS
JUtr7cb8XEEmYYPjzjuoKXgGQds5qqvSpYgDGjA9FO09CgfEQ9qBbb0pwVv8fjqt355yXY2bp9TE
jnwIEHnS7lw1y9/2pdZ14sfBkHX7iBZ0qFjXtzTqckmcGhumgWW6a4xlIH23Q+wleUwBCYh3Eqzz
9pihreLdG0zqWt0bzqDoYraCkyzRgiGU/2Kqo/9jiBpmQtliQxzUpU3WeBhAGhWGXoQ1NL0xWBJ9
UK1eFGan59SA7CfM91mwQZKGIBOao2WfjZob9cefR7HrNFFLlgc+5+P5KClCemR3DuQTx42ZHx1D
lYyFng1mwGIrFC+V6NnBLZ0xjx30J89Rb6sbay3Lnyss2Fk1JFwHVvG2N/Ki5E7lIBrDL68d6uRP
LwFAeVTN/3/QfA7v3nVKYkN79q8YZfE4EXZPsIA3ZxG2YYV/GycpPezQEOuILVgxMueh4VbWxXWB
4W5XzTG7jC1sBqfRZaVqrWxxB0pu3yeYGD9vB0gufkgMLIeiENu64Bq6awkX+w3xmovL2EpH479x
63uiXUw2RKX4WXcgMRVJBwAdtHlZlRNOW2Ufledj4uRBGZw4zapua5NM3hTcxnkaAuI3vyv4q48I
9xY8vTVrvM/QX74Od2joZVxGdWPoJKfsSin0BEfKC/evbvdef219CP/a1Rw/r9aUdi0Aeic5qCua
VR8iQgqWkI6/aQzsB50ap7KatJIR2B4lEiwm6zoFCSgclFHaaKXtwMeHJKGoBJiewb7Wa7sDUS65
M8CZHwIT8zQn1NH8JDV54kSdAqllWWn5Pi4TjkkB5Wuo31j301wHrMY+RSX2iHAPSRUvtvQTlHEs
988Cj6Wx5MyfwAKTQZqICMYpstM9V5usFuJ9Nq7MP2vcaXLL4pSOIdOlaF0FROXE51lDoxg/c7a0
2kFIVrCFbFfzOC2pSnpMQi7iKXzVYdC8kqVeYH9U9AqCSdd0X8FhNoNBnPTH1YsQqTh8nDQZiOR0
cK50lzbJ+LGF+DBBPtd2rTDFFbRhcKvENIbWzvTt4b/dzHJxw2A+pKYQUwOsH2Y8iSsd+OKXr7X8
oKOg+TYmXEfhxfnXGcy8PBb4ptpRm1d1OCNuKkokqsECc/x2+R+Q3Q38nDx2E8yNo74JFRDs8sVk
+uh/GQIPmf3pqktxZjF9mwidg59LcrNIn8ZTgG64o/k7zYLOWlYk9/7I4LffOYK54JRWNYFXqqrN
BG6qwQ3y9aNX2rYQ/dlrNRuIScs4pkulYIzfvKTZgnA4DiXbjmFprt12CKlP9LigHZCLsA6kF2Ia
LlZ9doD4IMrtx6ED0+Fz/HNDofN797+6Zer+5rNu61UeuRtESCdSTN6zz2DbG6gatoGoG5638k36
z4JrEzegHrOkBQSxrsO9GETZVpTFNZFTQxs9tBksCk/XrZElmNN62lZC17bVay5T29Ikpn65xsJT
E01b6Fna8WWJVXj1SV8D4aV+Y107LGsQJYXnL2ljkyk3t7V/wi891YLpf76/U8w1rMPkwGWJ8my0
BJM/iqZJZ3z2yXuctKMPilOm37JlovMF9nfcNXYBOT9g8rsAoFuNxRqosCam87bZOFFNRYghFf93
1NE/uXvR1Lk7clLYBc/5VLBPe0tS8QKns1Qipju71y9T/amDwMuuo98e/e117h+tfdCoCt1WmVPG
Ce0yJxBoU6kW98kU309J98eMpghrzVOKZJ5k29qdfxsRjsjRsb4DOqxZgDDdXpr+KNo2mianFVFY
HNJ4BH6QqOZx533ZXSPca5v80YfFxxhDS7DQLG3kzsdkf8x6w2o0HpD4X7Ura5Jg+ZQ7MnhMCXto
UOx52ziOQituLN1qJqshha5UWgOsKM8H2eIhORgVZf3EMgMje8auPdh0luVtE2hZifBNkafCIcR7
zgFAbQYkVt2qxOMjf4JVGWF5ZJxCNKgCIp6QV18jqh1RzjqiI2jwSzsVkZdYwXXhWd0CGCEOxVFc
rxiki6h6/tae0xzJyyrnEmHYSxOwFY1Idx/ZQF2ngkzENJbjJNLA4x6PHDfXqxvVoQ8o0h+MoSQj
2aPS9cbtd/nxcM/kz6zjDhhSYrqXSxY4rpVVKUkHgIhJrGdEhj8YG5eeEq4daI4Ip70yEa4IMwlJ
cRYVTfZh3vml0LJA3EPHOnoqQwxZauR6UbD3qBP7VQPA1H9wGLKk441cfvpott0JMVBXvgcyDD5K
52zi23d3rwcSTkp0CW9CxUBLF+wFvTJ1SgOYvIGQwQNfFgdRWXFuy3D8ETiod1TyzH1ayWiESHiq
vvPtLo6lI3buCWtKtC/bfhUTUb8QCe+RGfjNcTO9WQUPBgzzhP+aM7bPaBf2ltj2H+yHCA2m8+rP
iuF4c2g3m49IE54VtXNK91/geI36YvpNZhx/00Ux6rkC6EQ4aqNKKNXc2mPbpuUr1EtOf9jkv6QU
Q+7zO7dIamgYvKhbWH7H5egX3jkNrSb2nZf9yYx0Ii9QKmzi6AKxJLRwNagVyz/goNaOOy4Rayub
aRN9dXeS1P2SzLUeDG4NvMYUG3ZTZQU8B9DS1wsIyY30Ybx8x41Pc8aegQu1BcVZH49AYeHDQUQC
htpQi4aAwwlVUM41YoIjAuuw7ValhkvEROgLkNPuvVN9aNEu4ODLMUWFDWl/Vsrza/0hNXTiASsz
8WTCv3l2ZnlTOgahZWQfz8bFilwiwHyXlAogbN3ofGABP9/6a5qK74gUtDLXoo9BNto7dt79sasQ
el6n7gVLjRoxOQs5zjjZFQ3GdlxHiY3rcn2+8cpmPRxEvIeAszIFWz4OdZjtTaLq8RoMhtAb8P5f
XapxDh9y1yPzaUoYsBK5EGMEAQEgC5T9rDx9xZy+J8M49FRbwSNZ+oozqCwNZG3pKDyWElvDNlGp
DrSFYkFIZG3M5KWEjMxTFBcX+GF6LJde5QB30LJOPfbIadgs1GNR17h0bo/AT5sq1Srr5dSBJAaJ
s0l8u6eh7bGW59gTWvkx83EUupaV5c+RZwDqJxmjee3JYUiQtvdx+KyFxtLCXDYPJxhmXJ5AzXEp
MS9hGcuFesPd99ILMyme0N1RIGKGR/+lrRFVcb03nBc6ZG/wpsyQxFxVplZGCKiGpWSv97P+0sz6
pew4oceJsJclHXgMOvO7W3X8lyfeF5kd5qsngdHPMCAj57lb1qRFhjVoEWJCxAL0ucx4wxFAQfyw
y2r5Ck4tm7S65ZIQgby7Si5r9gJgzTz+dNxrS6AIrTJy89/A+r5va+av3CmlwEvIm80eVaxXqwsS
Yf5NHe6JPShtEQv1ltVcwslL6IDHOB4k+BTnvqj1AzZET/QzSaFUaq7adFye+rczlCn7UpGxVn1D
0aVRHEh3DIytLdHOGpUPziKZkLycnQsL5lDMsEiTFtAezCdG0toc+TBEhvtk476G7Vy+MfU5PKZY
H0rdzeBmaCL7h0FqsUf8BtSVIJVP7v071YiE4SkZTMDXwh8TrOOJs2otOOFBqtI4X2RlpeBl2Uka
DigKdf2rsWb0Nv+W1rfJZqfB5BbpuZmRA3CYaYOa9jKvGk3JrYCfiDQ8MXPc3ht3ZHI5h7Oq5Pww
MaXcS3iiZcV3kVBLbX5UoYfM/1w5ffMS1P0muoPUHe+iMtq4CdxPIDTgiY78lNE0uVXtfe4WNXVh
NUMz0T7PL+5NelbvHnsOGvPcAvzH28QkE9ELZiO+Qef48Y7lgn9TaGUKbWSyXCeX6GFC6SxAaC36
9OoNItbz8fRYXFtvMZ1kce5WdYREB2oSPplrPYD/tVbLnw+Zex8fAEY9ZNJY2Q9nTJ6keE42GE48
W5S20WqxJPLJW6z9YAUYd/jh4/t/xPRtFSuosdv3vFPNUXGmdi54xEn//9CdkRgn/uLhc9UzirVQ
8rxmR7jEMvSNTF4n/4sJTIDNTR6TllWB+GdUTlYiKIM0w8pEtoR6BoHyop75VEwaO0oRnjnKbnzB
tYfsHYGNhQLwlA+K4JcBpbzmg/bMaOt4jrwyUSblsAjS3d9aRrMJzz2wcCPoNmIPLSHXBrWbD+cB
hFk4NMEFn973BPxcpqNl9fM6h1jjAvmHXzl3S/cwATHzZOOMSbxqsfaw3lcJMz9MxeVELxGsb9My
dsj6icLY/jfipfKKtplP2uA6wnAf+fUHLjPaWg0DJNoaNptHihEHZgxVD9Z+uN7sJXtOF/lSISdj
7HoWNZBf6QUcNUT57nII79z3/nFrFa96ZITu60gbKsQEr0QAX0YuSs0gstooDwUk+xv3+vp58VcS
El7sFFfn/MsaGF8UNJGStg3P6aopdJEtzACrAoDl9sf7ToEq35ejLFRzgJAq+cGCx32JN5KSH5RN
akvU1pYqIW0S09z5SGdbR74M7xIDidnzrZ1xeu6JQO+vMfqj8tZa0sP0qflpMOt6vpyiKjjhJ6KW
d5y3LQqOAohvU1Ix2X2Esq0Szp3Yz6Y5EH/hK1SLRqGnDkQmdN2GvuEmC6jJ7gG3DFBFcX68lIB1
yfUJCwD39kPL3bxBP2WsDGuFvraawV3Oti8sTQcqe89Fk+gdemFOGHp957pJLAVnkWcW7c9+uZeW
sXP790DD5z0v5pOImsyIMK5CleC7DKkPKoQyVUCKkkxgBgsmVSQjCjRcQV3kDz2TfGga59yOye4/
P5dj60CDl68p2KB4RrE6+COmeyQ8f7pkZgJzdkWpRAzGd/z9avAIckFmpugzO4ehK4s3cCoZEkFG
CHNzGINdDjOu7YnKhlppGcS6j0m75WytTiccM2JYE2pWKzW08B64Efqnw6gbfKhD09BIsACdrnkM
udc/pEeMy9N/v0OpbM6ov1O3cFgbvjcp+qU412ylrIrKlluE6n4RtNQfx7qFhmvudxJTY7LJFpZd
77bUWIdtWXadorBA7FKY5PahJnQlyIRiXYu8xMXE+8+1vtdxwT7hBMQPk6/HdhK/seg1XpYqWmZB
MiLeZWUvY2CjibL7TwwoyuC8rOCqQDMqDeSMpYupZikhCpoKNgRuuyHRIUgkdkQ7QriSDUmew1qz
QQAgI63rQk5qs/v/2oJIlF1EfXn1iz0K9uU1jTGNtnvQoCp6cn3rZ0G8JweuHuB3NWYZXHH+2i+E
BHabOcGq1+BI75RIv7l4fHrrmDavV6khM6kbydmeUq/r6zjfEO0pHfSkvpLyauC8WenhAx7zRgv2
8I7zyEcIRkFW7cf476/y6hG1bSG1nfdlvq5mv7+hIgXebxlpqShlxd9heGdxKGu74pt5E3xTDUKV
MgXd87LUcIGiWhQ+Z1FSxPj3TgnfXe3GWyY5YN4eJNrsaUMTiEfGHu+9kZAo8b4xKhwnkx45bXT5
MDyM2QMC4JJExLpGd0vZAcCii40iENApcuW2aMWNpwu2pdhc44uRhS+kqalMBFbLrHwy3gcLMYFa
z4BMR+gj9AoK+8AzWlFKCp8ZoIqnjQ7q1IPpT5DJGYlXst36urLcOp+C738nyjezXvWHeW9hUP20
tCbyQ12xrKwKy/qkce45SDvG0XecqxbLLct1y1pXfuKi3R8NfDUp54H3H5nUIgtDEpNuKA4DCpn+
2wW7so1ZSMli3SDFaU+xnYPzsG8IxPWcvtuQ5Z6ykCW62g1nsARyS1Qk5Tf3zz9sSoGGHsdu3KV2
Q7pGRJ0vabmmWgAkJ8sQeyXn5gig4b06htgFC9iMEWm44lnZJ/37zDaKM+vmUiiUqSikYFytULso
iKEXulS4923yFW76tkP7RjM4MgSfGdoHS6LeisJIU4l1jeE1SSFvcrpghBNfaq3D2kkFNXgte56B
m+PhjiI94nEfRJQCxoMSdyBUwPJZINuc7FOs1PsMdbjnF7PkmdWCKnBfTG9e8gtuGUHv6TCwdY2H
lU+3+tdEs7KRSwPimQfQQznSek5dM/3EWQqlvpyTWII3byFz01qQR/8WYkNmDDium33Blw55/a66
e07DTh6L06JuKjhFPe06rmmucMyDp8RM3NyMwtXGnrgf3SYFCFrXeDnrEqs6V+0CeJ9PAjLnl5lO
F88vAzlSaly/ZUA8dUXl5AwSaQcK+zeu9o8J3eIf/TTCdBIs6XxG+1e4em8HeH6fvfPWWsXMR0Gs
j91l7aVpfPFF0uvOKXQ9vbivt6gEq0Hd4k+d1IdKAtH2DwXGF7UVA60Drulm0uWvzLsWm7k5n/iz
N9OBrmcTQiArH753swDZL98LP9tLRAb29fYwKleXcPV8XFNb1j47jcW7tJ5DkG3RufkCMdcD+kAY
6ANqrB1vK/1lhKs0KwcJ2Xq3TPW1ZqqWibZWz12PxgmIbgQJ6aV+Z5ScbCLpqU/uBckO7EhSD14B
3fG9016X2oEWISTCnDpanKfJGu9Ht0J2Ue+ItOprSLH6k4FxTeXGUCN4F4PSrjH8RvAQaitHG/mf
+98dBIFDUi9FOpns80RNwKI9jmG0UhU/0Rqg6fjX5hPJi0sCRO5UdXVjQvzkvWsvKT4/+SYMn5Mk
T3pnYE0S2kM5kFCHOuuKOaocI/6sHGnNutZa0O208rj9LGVQ1c49FHYXgHhlQ7zu+9AVK0ap6yNQ
7a6MP4wWTyH/MoZ1qvM4xpi1767CZ++YC0aQIht1V1OYClMbJgbEP0Sld7WagE3olk3PKvs2LBt2
QMFggCQr94D63m8K8RpQshC2FImqvDvNaLdOJNj1Kv23ac4TTG1Y8cHQCaxGEY1AwopQ+dF9C97y
4/bksaDwyLcy0IMQgR+6kWOc4t3/ngit6d27nlcYKBMPCBPK/15Z31t0X8V49VNEB/cYzTLaLpxv
PNSLlyjmIxuqnDpdNV/opdeBudFh/zVFZFSR1kRIotfKUR0DxUzxcxjSAQuoABKeeX/yUGSo6a0f
4TKoXaFcTkgbsDaZmQqDqBYGFrtEid+Ru39j/dgy0JKk4ojsFuNnh7L9Pm0w722dB2eWt3rwamzx
z85naWRv3Cj9Y6N6qcIKdZm06aX6NSeDbDTNDBjLIL5a69b+1ury/nKKNkTzyS3DjtzL/v9X7sjN
FvtsRFwWnIPBnkR/G22FA9XpU7nLnAo0w0gy+phl1Be7dGQ1clmhN7TbTkmqpfaB/k25Ne25q84t
BMC8NJCP/eaKIkkT1Y6RhckfwYQR3ZZ+zMbSRGxJ1OO5BsqMxl0SFTewS7tIM1SLNz7hW5Qg5GCj
XJb30KWzY38JvEm0SV9JoiCH85vCg6xNckde4COZq9kpt9cPDNfkf4f30mdGLW4Ddsm2RFMY7Mlz
01BunCkY/bJwUiktyNAdjWT6DoxrRqipDQM1qJc2sQhBnlcut5X+vYhuwIqexVWSUsKFJhCGXMyw
xh767jN50jWs2t7UZb0xZowYAVBhEnnPBx/zlsJLc90C9uuJLMDPoeMmubysdUgWHHBsV2K2zFoE
3bqHFDIMfCvH+8JROZOsJxehJnqBdHkdthvhvJZqTtOj/28FTBEr3NuFXnzLyWVgYWY4Oiwr1av3
BfksY7HjTcdRReRceK/bNXG3fChjVfpW8LOiM8trTC2pvjxugiDx7xb/95TAMT9d806NCcgpe93j
gRWAjfrUAxI6OKUg1U9l/zCAkuYmW9f7jBg5FGaCLgZ+n02dYu3T4ogIcWeVEPyFARj1Spa1F5XL
SAizhB2LxZi1TZlXyK8rtmK1+vo10BrTCgDJ4OJ1pgBwtMKUWreLSx2rhgfL8j8uP+1qR5aUgo0Q
FlQU7hYaSDEmkIuIzYncIALyF3dtbJY/xhul33DLxLm8cjHPHt6HLbt0R4DSVJoyxrF3uX9i+c2c
2NFFq4xcQ+BZErFa6m/g5Ef+PgNL2+Fye/4GBhpG6AXLo0k89eroHwXlBrwmWRX69XROT+IofBb0
1cUy+z+TS4WK0sOqcvwXERIrfhqiZTDmI9/C2K3PdvhDkuPej9dWSsOi4v+0YqU0WWHTIPS0BAIB
3wBgXCYCyvp1kTb8zqO7LK001dwUvlaMKetfAnGnJJosvLCyVz1XcDYP07YxrraAhIyGG7KLAKl+
7TujEBnEgDwGRnp8RLw9pV1NgMU88KT/bDuoS1NInZXbNmaPMmr1K8OryQPRUzjgOtHgsPDnveZy
bPgfZ4Y95tdo56Q2wcxe85ejelLQ2g0I1r9c8UEwlTDPevOJQGw2z4P6D5iFPRCRPXOdsbq8XzLX
rMCA2zs4mZIX75GsxVMjg16uOmleMLcEA4qxOUO1RsIHaw6D0kjJGqpldWIg69oVYygBdUkW/Nuw
r8uFwuv3h3Ed0RRGf28nYZxVRe2EWCtmfQisIlHIB6IewDgeyO2TlWchUFRtPyriJbuMLoUJX0Jn
spLzb0vsLrcRXrBi1COmM1LeAPU8Sbe4h3p44Pj2uBDsgVN5dF0Db/sS7DUG5I91CLxojjGrbN51
zdSGoT6/GfaLDjUxEe798YWgzJQCJR8S/JyEetk+Ctq6+gPLC33y5Pu7+7CaY9o22ThKcKEuzlvc
30syQD7bLSTqDDkO9zJ0ip+4+o07js0i6DejMiHD4damLLWE73hxsaDzojueZtjLRsGjE/ZdquPA
9hChmHCYrGjAl+OuqwakUCFcIkhv4neD+t6We0m2MRe4tihrTI26ynP8UYm3nE+I7e09K+ZVSUtl
Tn62AFva1IbsB3HKY91UYvJnwVyWsuw+WTNDAs8CW7erlQAPwnqZdUMmv6X7gWNtoOXZFZLHz+si
Qi7bi2qm1jcS0zqDNhEl9Dkzp3rjWXDjy67ApPxxBbJzGC/nPo16zantbYlBA6gjuXd8YNW/7ds1
x5N7f+ucqWtTKs8r4mM+D7JqPa1cFhNemZWhShuG8XipFc0a1i9QJ/QX7oMcrkwSuOCdBSOP73FY
JGLazsgLF4xWUS73HQektoO0KUTvauNS3XUDpRGVI64rXNsiZzC2UT6paS03MEK6j6OVxeD8SzJY
l9SBzkj4aDJQU4caVIvYIsezqHCbAvHZTRUO1CMZ78MPbPI0kZImqy5kF6iGkKEZvtYP2PnuSFTe
cVbmoJJLFq/sbn6335kG26naZPWp5CdzNfE+EDhDLzsJYdMrCeCGhbWnHfJhsPLSWtK/VMYDh/48
cBB6hvX819fYlsXMYNK4I5H03Y55fepQglGwuyhsJxZa3dywjvFq2A/+vH5zgQB/3ycu5ZNjSmSu
iLxuenVnQMN7Gg8mpqsClXK2mHppMY156Dm2BDlPxRo/un7U5wld7kyhyE27ayct1YV+e/cgK9kN
+VQKCEcSoP3bageC1Fk3Zg0W572AUkQkyEJPmKm65cacdyv4EvBjOCYAW9NMzmFehqoWds+ZqjEo
Mdheh8LJm8s9UkAfSDF0PeqvPtnzFmXolAngEYsKMNOWWKdh7uAec00Gnx8H4/MQF1kwVWdXm38Q
4Pt/zcqEw0qRqhP2/QdJOhqHCN1Au9CYVR2q7SwwzKtI+VHBRpCIhXUml0yT6KPt5NTIXStT1lXv
hFP9luFRWDWXZ0ou+5bdSyNOiREGu8C8pCz51hgbdL3aPdWpuXVxE3spiuAB8JS+HrXJ9pEky28i
WBpChqfM3oB9lD6KJqC+reQvekL8s5DD+5dtomn6WUNoMF6h9RODINnc+X1OnEGAIjGeXqrw+t8R
4Xsx7DEjL1+S+TWcgOk2qwaSFC/1Lr/ppHzoR8fe4PPQzZkJE7UlCzDbnYt2t9HNLmew7GrjADUl
kiIpgF4RwfkD41XqMRphCNMHsG0/IEe0Ia9F2DMDSPlorkjEOumebVHGBrAWRLbXk7FCyukBusN6
QpLskLw/Xy2GFsLG1UzYcO7SvdovxH/pRSmPvguqzR1y3FrN/kwdONfrxrj5Mi8dJj6bYYrNKbIE
2TwbnK9kk2iPD7m8SgD/NXrYhk8i/epRSPjtOK3Umr8yod05h5OLfRBdkyxLJVlsISJpfwhKD2R5
dfXtUFDgT0EExyv15zVpnUadnVPI0ov31PJzjywskQmvu04f8BxLpQlA0rrSMAbCGu1PW2xlDyk7
oqq5PeVrOQnl42swaJ59uc+y78BZqyDrpa2PYSaywa6lVrNT4sEjRruNerffHbIl5uGzfR1bpO1O
BIE1qQ/JlAIfgIv4lbPyjfKfzdUo44cgWw1AwGx7h8toixTgZZu70KkJJ5x+9X2fFvajOCyq5Pc2
PZesInCSu6VV17qBr7ZFn3dSYnizK0zQ+7Iwo59m2pC9/UwbcaDTl1quAi7rb+o4QYeaxDMYXft2
3zFSo/+6NPwuifAvCuw4PDJtTSAUksY1HBG4XzjhgTzVs4Z4eEO+2g9tZt0usy/1lLRRQIcgQ1En
P4ux5AfyCtWJH6Dz0RsSc9iM+bCgDnllpKdT0lirTFdow387lKUgEJd2uOm3Hxq2tXMV9Ls/bY9a
0RLXlNa49ipj5xIXa8wOiD6doCoF+gUo7KMANlvnf8yfhZs5yv111HhFIJdcZsUZn7Uwd1Y25KQy
Q1TvAzUrvF3SHzfsUeqZA07QEvsKmoCXD8Lto/cmmHRekyr1B29tsUSGXC2NeDiS0coJ8ordplxp
KntBB85KG2gNJUIsymSUuEnbPRuc0aQc0P6s1R4NNGYvazg38LsaIVtHIeZ7PguOtGWuu1CDCqbr
kjWMsrHpDB9Nh88uCIHd1BV63JIQNnr9WKgYbfdNZ8vo8yUydcuhw8W8oLR8o4oHDtnhqppcQS7V
W8C1xgmRZ1c+3TKONUH+anIQqCz+9q10IQ9XP5zPVtUrVcEviZRv6+2ybNpU8Pr11qpZyMd+7ReL
yqbcqyvDbUALrustK7MbuY7yG+PCCL7BhrR9OqMxBwkKuRrNo4jKeHOA+JBB5JNnsfaIItcrIPiO
7ymCUcmgl86uZTCiRkwWWlSXGnpvJtJDA5dwLsZSDIjt3v4ZJ5KueB3TT+hiQcXDAH6hQxwyaNee
dKUJeG4kybYA/3TOTLsWE76+DFe5dwPlWUD3eKX6CVCidFC48z+qeGatsY6OGcwVvOQRnf0bNhM/
3iMB+3BL5IHXUtZyfUi0YaSJHZo2NiexU25KRDaOYBrN0AnL1sWaJ6AgDui4kCYxwPNbNmSICdgY
Nz+0DkaTPryAKGFoXKBARyJhIszsSbdW/6QsThaxQ9LKCnN2fhaNMAIPzdffiCoWueVeph/YQ21t
jJwzWoAtxAZyj//yLllcR5qCCuBkl3WbdK76/ClZ9DvnS53GLcn4VAGk/IiWCovaK1q1r+083fpU
M3B03hRnheEJcJJUCuUAua/Tt/p85l2sqYJSMYuVgt5ncwNVnkRDt7lh9R3XVH+kH8fBY8qZkNwY
eS1jzb2+V4CUBR6hJHMaBDdo1Ruj1KLdIoTumzDSa2fOjRMsl8sGF0D2bauKUZFX+sLkXnIrPpAW
ER127ZqQK81+Jy3dsSbmDSMqYhLIPGNffqAg88JA3FAhoCGCb1jG27it32URvxcdK3keXTqhMTiC
vsD0xjogLyU6NWYbQUg3V+YwIGESCP0repXZZ9kmkRC+OFeYSf+UzkFRPoGMna1Z6/4Id7KOWLKs
HFrUv625ygmDIWJYPVPHlc2CvsJeY6t7tJe1wzGUSIHixUVK5yTz3irecRUQH+uj6zYGWBrS4iPf
kUhWgVBOjltj4t1rGI0uZFcJEnvTVKquXsYckrcTVQx12Su4dW4HBspr34qoWEEYPsqo/osXlngY
Giba0KiJuRj2fXZgll0uRqwNDB88E2goeB6wt/xM1dIJQgsClO+mlrMoChSoV0+q1j0b2WkGvi9v
7/wj0w85K3JuALy7Ot/xWrweYv4BB5WxMhVEV6Ekxw2JRsT5hEIM1Vso5aQcyngnJ0l/QJBlu6Fg
EnMcazb4lpIbiAtpYfD8nwgzi6Fqev8ze2RO/3eKrhXUYaCRSZi87iL1p0oynDBO3fJIS2A527g+
aTP8n3igEP4zMDFQNm71GVob6Nw9mBjPZLR2ahU35x5OE2ozciUDI/ahNCFjm2RSvdOdHzOsanKn
RWFzdvei+GKS2XR2rUmHHBKjKxRJxSywzyXPG49thC9Dj6NNFaV99tGmls6CW0mMpU7+0Wknupbc
KcVZoCBxNAr83cH2ifmebAZXDck/g6/aErDfhldiPxUYuupbgi/gxjvyXtlEi933UG00GiwHnbrP
KgmHZrQIj67V5FsBe3MO+aKu4cF4BBmkvMneXmvo8dTLzUPp6lDvg8VZ0au+avsLINqzGC83sE/Q
VN76TI2L+DRE6QPWSNJcDqTNgTABqfv4mzk11A8HqLAhWuJRX98TpFOY4H7Ixan18mDM1A/K99/P
YNhgKZamvMn93I9k/lncum7PpJRLHBVLhonpN2MEsqlUoc0JnjUEsECpvUGx+oQV234nzyguC9am
fB9SUzypsh3poQE00bzWBDnbIUu1R2f15YQ7cTjc+uC1YFgRQn1Jb7zXMTvK4kxxp31wlUUhLbmJ
f1RusCCDuIZfUozXXbiVaI/+7oZZEgQnzLiXA0jXrQ6gtlNlSbKsl3uxGGhFPbe1hqk8sYwdKp3I
mALOs9zKeAf/Nhmn2nTiZdgezzytbBImFU4kyJ75MnJtjjVhazvbjQ3RfWWg9a20Ek57ug6sTymR
DQdsEvxP0U3cPV+levx+eFVugkmxHLjg5m4S4kRDRhKM6ByV3fVEDslNQw//BLTUqMgGTZ4tQtqM
cyhYXZwJ4QMWpFUUgo39Bubhk1sVXRWIqSTYJpuFewmAjQ0ht3auyxUaTB9YHrRKhlgI7V5MAruH
clihmbxSPWkiYxHAzUfa3Ifvt/59G+BFxC75DTza8UVDa3mPJVQxUjSZvORJu0tRpPBJFsxO4x3x
Kw26tv3K9vHl0sv/CMMIgiwzi4gYhX+TDaDbUQsGCmkTeRzhvOjsrPmyq4nLeqmnMkYDx5vA4/QU
VVZZh96Lj2XBSgPqWlAZlPM2+N3+/66OZ/A+HwXSafWGEWhxKvE/iSutVQUnO5sLtNK2CL3J2WTx
F0UW9m5wbcAFX217KvsAqTDw4zRODUu7TBxvo+kKpC8BLTRSvyiqSHmgc0ZZwKzEACgEhG4WyjDj
+zOZvNh04EQ/BZC6e7yI12/2M4pW9uqykZ49LpYWdlRwUg4oTlLyMJVK7tV4pCCwG1ekO3oUa5h6
fIs/MYGFn6KSvBXaqK4lwndxybiw7GuzMTqVBu29gEVlTaR3hcva9TRNWXyjIBCaWrf40P4NejWn
Q5ALrHPKaojCoVVwucTwr2FtxvppG4AKxEaQeUTAk5Hz6Z9pUV3aocNJbFTo6en3DYNrGh314HTw
8VxlrmRsmwS2QYPNV3PWPfDFKyvRydqmwlx4wJL8Ub6S1eAAcTG/KfMIsZzwHjBWqerJpBCu61Pl
YHXUiHArES8kvR5TNsIVJPNVU1AevwPl8hHUvJ5ks8CYB4LL+/JsXT/gBhUDJn8etxC50hiRm45D
iogM90ENiZvPQ01xeBCFTLU/6YPmuIb9nhQSokFe+6jEc5c921Bqa3aQCjMc8PbxHTA1/IEXYKTD
4hmJtcef4h1OXugTb6ARNaKkusuVvX8jJLSeLilP6CkjIq2HwhGhI4O3i+4/ROpF4xNobqNnbhXn
EPJvjCQEG6sJZfOTDUm8++59Pwy7ZGx/HyahPZb9B6A84fTqPiXkPSTpD45U40T+plK88o0IB9Ey
L2MgkP6RLS3zc7yFtxE7RxSwiUl0p5ngQ2WRO49dz3E7vl3L2uxZAiUnGwGOqqLe5kI2LqfU4om8
TLTFgfXnI/tGAqQBfKs5sMrif3oYe69nRVP1EKHjFxCMktpZn+ZNe+WS/CmXTzCwreYe3kCNPtal
rkMxhXvrTbI+zkdEe2JHO/PGzn3AvKRruw1pUrvsHFRWQupfqUYhWnstfK11ZV7TqtDR0rYwTcWm
NJMW6rfpiGp7MXo3X7RJd7i9+emEKQGwnO5PZYEQJGI4xVmMfBuejQNN+tNhCmJ7mbhzZugIw0XM
EwS5phj8HbqHBTE9M+4YdjZhDl40LWVvY+4QwP5jaWDhHrqzunL//iieLGQQckZBxm8rGDy2Gboc
/V3LcfTW9C4FADsRgKGn80cfPXSa7QiWkyCLacbO3c4wHJdyG5Ckm2DEPIqxTlro1QTY0e3Tyriw
uFdW8KlLRGUzn3PRzqk+TQeGKdOBHNSYXoOITGMLLJ80HZNkBl2aVcRE2yW1t35AmfwXpGqQfhlE
nOdWkTfXILz86RG7PvpRfLHdPCY8f57W8ezRxYQ4unFso6Ma5rDzsMPdMGQyo4YIua2IknrgxZWB
7cLaLvTzqFabZ7mlnZKAYOKs+kCFXMA0oZHUpMjIKOdgzezgERc7Fj83PRuB5+k7TidL6e792EY/
ATXFc8AAT3gxr1lPFXfWDPf2nVaJpkEqeHDNVNTi0m+bkpP49QV92vWFtZlHQXFs+7REZmdREOy3
VWSWwANWEmiBsXs0umvkUenp2WEsHyBum3b/Ye04ne7IGWtjR3cZJGlePfkcU6Wujn1U4tssJWjH
CO6KSgLwejSNaEBX5ionYlX4k+J/dem2leSNCB/DKOY6K/2IMSd3kgrc3KweLtTb9lATz0CJiUxO
n95qnYgdQKYh2cgeqvh0LJCBvIc/8wSBYHChS42a0V/PgdLp44ZFaiKyX6uebd0ZWpm8RLl6l9SK
JDMyFrY+l/lZfl8SfmzF519pV50kGN0JjJiewmbuxr9UiFQ2yT1JWrPxErutbJv1gyEwju6BW1X1
FsFMYFnc+bARlw+c8z4wSQy7NhBlNOrm8P4vH6q8a6zZ4XpBhwjKDntLsucZzT26Mteo/zc0nTN/
4wqdK1r4gt309hXd/9ILrsLkdXLg4yWvwyNI83TiaBV+7kSIuc842K6eSN3JwoY8XI37w1n1AvIU
rdNHWEdMp7tlEoTHDlZrQzV/Ddx3GfyJwisyiVoTeqAdqABPKskqrYot+fBs7115A6bgS1QyqMHw
zwIV/IQHyGSyrI1Jvtt/0RZiN3ze2O/C154NXmTIns0VBVTObeSTFUu/8VBJhR0uV3/yUbHB6W7P
7XItUEJ3Q5Mu4tMz2xmy0pciwkgGELGw/MapWD1d6EricCNpJdWA8Q1T5sxTy617rFlyd6FBKSqv
8aZtOb7TSSMUc7Z/swgXtrrlTmXbHsA9A8TXW+k5EYktsOZQTcKF3NlZa6DXSKeJotByMfTjcYLm
RkoIQB/vJoTrghGku3hS8reZRvTfcvu6aszd2dqc8QvxYrdKlOu+GAdtYnKjfBjqlkxjwg0JmR9P
IFO/K/zwX7yhGrCOkdZiAr02mPXOWcJnexARqXroYXJKOlpIMDHroekJUOPhVd5IAoVHNdU1ebWO
31VvO9f4B4wn622OXXXA+8kva2gATZJ6bYg3zUoG7/5VG9CIePp08ZGqvRvd97EomsKz293aRBgL
hr08zidfeYAaX9LoNFejIBxlvkLWiWmXrT/SHvH6JDv5+MjCn6TGaR3RQpyNpKoY1fSS3JHvvA4D
PR7q8VSQRFmJsIC73QjL0ysH/T/EK3TFSnZURCdHBBuGvIsTMim6bUzstocOf0rjF1Vu/l/m2uix
VOrreyrYSfqVl39LvMfW2hYCPG8ECzuv7nGvDEIDMfqzMc36H6QNyvaMjcqqt7U+tBT1asrb4L/Z
MKz34mSYubEN7nH68FnXAsU/B3cLa1nv0y3MIellzWTq1vuV6k/3HPPDyiTH8ZRo96HUeRE8Y5gF
BPBvMorV+JYWQx8WEVa8zFjotdan+68+M+DXwfNu0THyzIYUNDBsTl896OYTxdsKmmtMo/jdTro+
kuyrJHOYvGvpXcG9ehC/mTVpvRRTziWlYHf/cv2Stj3mAb1lGqdZX72B1AUc9NyBnzDakuBRRHu5
6UFKAdHpVMjHuZpZrIHOcjEVrBOWtl2jfjdyB7YkdLA1KXWCVDlVdRu8mfYcfsxXRfuDLQbSbrVA
6+X6hhFPILeHhixR2qcA66JsxeIoh0YItU4ZAJDz/+FzcQPan7w3zCuBIPA/nZ9P1KFB94nQFV8Y
WRxbGmaVNA+2pLeNQXjXXofIKHwEqwq4iwFvxuHU1elUWIopOH1IbpElKSM8VpTCOrLgBWSe4+Uq
PbDnMmj8nbGCjDZIpkMkSOUE+e0ssBCMBO2MJqVkY3Cay+dXobQXMJUGLPo+Vfn7LIgMCTiA165n
b/so02Ib5RbJdrwUFltelmJErJa4zK77sI0o1JxvO1sPqcwgLatt+PC0e+2i1tX/kNblx2/eBvnC
RrZ39ZBDTxHIjQHU/HPciMAeMnZVVU928GAYogWsfL1oDgadYa6T/e1L3+m8C+rvArVfF0wliz4a
Rb6XqW3w5OE55idTf8bqCUM3JMCxPIVOY3UBMuRv1ZhAF+DMnLDRacVL/6+VRylzJ1s7zufXTWcs
y/9fKaYSlTLeK8M3XYAgaFj6scQZGhMG0V6VXn6S8Og4TYTbKv/c0U88NGq7OfLHG6T2Mio/iQqW
zKdT4usqmRhBQ+d63GFYRNr1wwwDdHaIUPFkU/EOhAukFj0l1jCYYrJofD26noUY12HSPmxRlZw8
R1L6zAg9oxxl17vfzYLcJl08AVdAJWBrOTzPI+vVkLtrriqIwidODKw+rmLKBc33aCVqU+MbePze
APSgHNKvb69nT18glJ3sqnU99Kt+R+t3MFU4PJBqEMFSRq9Ort8zxFMQQ0/5w4BY7eOZxs1zhmcV
xOQ4rFZ3n9ECpfcSMlK3N3XREDAdrxGj5w3/Mm8HiOcHz7q/ajxYUQI0iNeH/MM+/tHCcagaLLn2
xP0oUpnh+D/irnZtnfG2GHJElEtxuOKvTpygIhNlz4jV69MzahyaeqEQAQKOj0oZk3Nn8dES6ZsE
uOfzKgPRXpJl9fPlBjITR71TiEnODDn4eF71jZIWntTwe3TKBH0ucDqqdWPvKwnJyczH/ZicsYH2
3n2hM4ks2SRHbk92BnjbIvtHVAI+DgWJf4YaIILGcTs38x7Q8XwHEjKGIjjxEJeAzqPswFp0tEDx
4InagxiF/XBH8lvD4vlq3qBnJR5FfwlSLzciUkwsmOsz1C3FnGCsd9wRHAM598tnqG+QYNlhjlIo
k41L4zXXxNIMSCk6bB/sHGvxoPNLtY5yX6xKSmVBJ5h7kqD++cse6AhYbNKFWa9yGP9yvrfKphOO
36po+xMUsiE2cMWiklQHyO6/FMV2S3ygvIh6grSq1+hlA8VkRncT8jovi6novhtQYiLWVfY9mUE/
GeWWUPf7+0D6euEWCBNoPIhzli9eOYao4lqohG0WY2wn76ICIfgfrpm6VQhShdrLtYpP4Re/Bw+Q
3kO59eawL3DQd5pO5pmt4/MUa2EMluq6U2qmHzP5U2jiL2aeDd2IX0N9KOUe5h7KcF/nL6VonV7G
W9FKLJhhF7vTq30yzvM1OJRHUPtqSj/zoeCEWPYdOOkiingJJDmRxWcVPmi5JgoJT0ANIhc2NPhf
84sTenV6DDJOgfDYcUTHgxekSGfy04yTf14C5wRYsRGei2RQ8CFXoQy2hi7H9psjhye4j8V2R6d3
4cGHmDtw+PSObDS7HPSW4Y8hDu8VBagHgTpOZWxheeNom2LT9+sfc6tyNdxm2B/DphjTxFXvkPhW
9dqlHNpopjv1D+ohakIoSOyW0zHBfouV/ZuFwyDHKXx0Pr9/8YJgJ6Ej+7bzw0KPjixHM69Vdzt4
Sl0D73TqIL2cn7rm5bJfJVbN8Xua1ZWUh3LYu+SpNSu0oS95ZEkKx4iUV3nwFaM1nS1lCiRijzzJ
9Id+my4Oht0BkwhEF4HjNIUgDCm49CyM43C8+YQg9nA8JXsEh7DmJ30vWwOxifp5+FM4SN+lZ5KR
10oCVH+ZmIw/uqhQtDrxLRFpAM1U3XXeqc9L1KZAaj7dZQYrPFJ5FepQvau0fbHST2vydD22kqlb
XA0Uwz7loRUu7yrd/WfVNu8+ZBgcNzk7OfhCUIT62HHeL8G/m1M+6Kz87HaPP99bk9jdNsr+hVio
0qG0DV8SkDqh5piAJjqgYXHD7dYS4rG4yz4wMxRWS4qq784WaXMppNro8KfXToSljbvpa7Km22Hu
figK7ExOzvMGLKUSTwDsQzU0Oz0MsfQ85VLeNDHW0pWQj3V2uEG7ja8KvXLH7xBYq2kCQ8OqSSIo
0Jy13BM40KUZEm4diw1H+n9dyHa82BAWNcOEeyr/f/scKaK+/38HxYyyZKl4cXylD0mHxE0++V9p
ey6p166rBOdE9R0TEIT8h3TjQvZAzmNo1GgffO1bGsGrRLUm9WqA16pnMnFdT8jAmiYh9Bg3b+pk
3YgM8YkRNlzDV5VTGVvPwrj/YkK1QlArY6pDg9HUGvCMCCwDMqqYaFIabwg0GPsSEnzGB4GyxiZg
GNNMVzWh/bqIZ4EtviyB3+lEUFi+XgQK8/l8ipND48KICgevOnC5TqMyKWndA2XtKWBlE86lBR5v
86YV0PlsNs8kS09Q0exJL5hixdD8fFT9jmWWIuJDwVHug7AH6wn/jDaiPSpvY1VVYI+JV3eHrY0D
tFo9jImsCeTulTtPEml5cMCoXncbl0ucPVqgc1Ynu9I0VgeH01i+qqRgKe1BEoH8fibX/26y83Cy
fDgtM0djcmGIyQeMNcxOflvupXIo+1shWeIyfxE5Y0ogCI/mDYC6ykVOhBpxUPGETvCGpGDzXS59
M2ZB8mltQe2UrWT/YyqFAGYBnUBK776vv5/JantsW4j635UDR+53Qk9stOjTtUoRXml78a+ULMzZ
GfEch9ZWlBvTu5QvWWFogdVChGhqJEmc6YK405tEqAV9NMNc0WCVwSHjb3FIi/4Uqut8BislhotQ
aYNPc0Dr+cR6NZnVIm/KuRYL1OTmLs1Bims8b0kM7Y3b7tIF+G0RiPuq2K4eRLhot9s1qDppG1c3
7N0pyAUcjhyMbaZFN9Sds93DWvtoCase6mblOZeEuzY1dQQtrcRgVjRPXrs0ZqAXH3VcjzPBPWjn
dBpidNkjSWHpEc9aCN2XYR15dcs+dkBRc+7SPokMOWSa4Px8VkDv+5xTEPav+4GTjeGOcp0+saiH
wK4D3AHup+Dlxy6C+aBBu7fJWWc97ViBBMYbGiAeIPCz2OvmI3tsak5w1mcBcwTjVJ0+PZBR1KyD
N+XOiBwRIPVqpaujoJ29gt/YTIsIOoY3n9lUVVkQSmnGtC3piB8Ki0yi2TjqYbTlU3dWnw4ETcE2
c/6mMR03dcgTAByVub9kHEZ6AvUThicamdMQ/WLs1w5taW4KMXopBR+8PWS4c698tG0AKtSjt8GE
jLhYxqiZQyiLWFFmJ9H2GpKBON78LfBtRGzX/bt+pqrLml/i64htAvPpc0NQzg8hLsyiZpX81pOl
qxQEvglxUFdf2vWsLGh6k2EOyKEv4nOm6rEd3jzIBOD1duHH4uYLWJrhpPMTk6NUxqtbQwR9gUl0
ofcLmmuWz0aq5rwRqsQEhV+Z8DhY60A2atL52BdZCwRrKUEX2AAtRxvJ780lmDFf8zu9xq7PrX0s
BkCRdWquzw3hqYEoXidc8+HH7bS4tFsb2lE1NV2Hqb7umqt+T1tr7fDZScUq9LU3mam6j/4ZJu9H
s1iJ22kESafviPswMbp3KF7yBMfP7PxlKfANFLqNpv/9OL221GxmsW3YLMNOQsUXj/96rfDQtw9h
RVsWKnul6Gd1EncgRbH/YQZVsvHGAhQVAr/o3B8AEPCEIXbJ2hXwlLCPvwswVfjgynRIZm+GR8OF
2xPDBhgymwK3IKquKGi8eHHZyzdX/pjwHgP4EvmwVqnGbTaprFpmNFvcNfGBCKQMiynNSd1N//pm
id4ysevJqC5c/8Hf0FIlLmTEXmdpQwSEi6sR++GHTpBzLGnR7H6Wwkdy3XA0DYNQIbLIDNB69yaP
TQl+lLDXyGgn6MxRU3XNSIAi7zQLZnch46eMSkr8ijsQFm4hxwgLPAVb2aDTn8zc60TAsS1JRnq6
GaQgRNElBkOp8v2cHRaNVYz1ggQBGkKDlzo9kUg5/wYe+B8VNIShwmhNBd3sKpc2w3HKgs09vDHy
oAmzXSHSg3FlbYcB7g9mgw7LwCUVc8mnexPYwh1E1BGaMc39Ri/Mh9UEGMn6sRA+gPEmzT0YixXp
JZ/vZ8C9TlkoJoc1Wofk6x9UPKnTNoEMqvozb9DsD5gQbgNMSHAHPiEFoF/LF7UXyYgYVq5NcXtC
U/xriCv4x64YDdEgOeBQPXFlVhJUK/jadfumvWvF81ZadRmPIirziT690bR+tajLeDo6EW3LJgtg
inyOtg37nBSaWswQwenpbG1HT4gL98mmH2SZug+IilJ2/u8p0ShI+nqL1Pl+T6+PCFzmcCVhCC2+
++nNbA8tYvoTxVDqbctHAHT1BHRkeMaAxEXVOTnptGwNU5rKlhGbKTqWfsrmqQEp9AIptQPE7PAo
gW9V7e928Y58W4wZW27z2j64NVWHQamcxsf8NRYo1FcVAuC2SsQcLsJnGskPvHtfR1mAJMgMHZ5Y
bGBQNOd54r5+cuEVbVXRXvsHC7N7YMYvbuAyEs7wZEr6qaZ4kjjg7DRsntlqRf07MnAQZmdJtPrJ
UKI1PaZwK4RdH89I7oXOgcIDejuaVePfnQgnWHIhm+RgpQEexaJVExDl4/W2rO2V8C5ZpgfDuQuF
LgLCG+88Y1IWuA5sOptRV+jjImpgIxZdHBwvVf3+4QAz52dZSWQ9oA+PzNvQqLnvV4zS44xEPaRH
K5fACGWRVdorxKu1zra38jtVwrE45nBYBuyPJ68Yx884bLdLtHjbf5JG7eITK1y3dY4Cnf/Lor9U
PsyWpC7EAZP+kxsp0BXMYQ28jtwP4kRg0zLtTWNuKjqg3+QMIgfXlxy/8V3LA984QzeW3wlpUJOw
LBdp72Df7k8E9RiXpZFdmohIiIXcFmg7SFm8/6eMf2GjOUoD1HpxGLXsMDlcKBRso7CqZv7hO47B
5bK8kJHHiUGIRPruOHGzFY94gbkrU16CjFDEUwL0gsvCrjVQCfgJi+oz4ZRJzAgICHefTJNhuvBv
c+w9WwFm5e8nQiCJDdCmrti6OP4XXUnnunox2nW3Q3DZsPqiQ3H1fL69pFNTil8xPr7C3bOz4SVa
6lqpOYVRT+eTTp7+X9yQfb9pLBCUhVA8RaolJ0hAM44V3DhGXqNnNgq/dX16BZcVIc45Q9yOr0pB
x5TJnMvUfe6J22d+wdFqKI7+oFhq2T49B/W8QeaYpRXO/nwQ7WXuRjijm/XMdtx/e7VBNR/uu1Zw
9M5es9aLOc5uPhExqn3zjIAqfWVEVdA+lAk467dkGGwl6ZmXsJYu22lhlVm1h/3U5w0jEZegJLe5
64LrRZMtu7OGeClNSHezVj/pa8KiS7LLEo6bDmSWqp96dmlIZQnZQIEZ1myk2tal9TCucV+62cyM
iS6OmQhn0g8GmjSpnamFq0ehIQA7AhjfLIeroaSB8tk8ZYHoS1pqEl5P4HGA8DsPEUyd8s2M6itr
j8Y3FFYUvWJ22h2HdQ7qbL10WJgcqg2swIxZcOZ0nXFcqyQQ6h1BczMhlYJSWJZaYH9QDs5w7etb
Kci3KgfNiYMEFCf7fk0qo84K8yOHW1UXNNBsntV8mIphFpZrXPEA9k9tTQYbZBCa1/lg8W1pEES0
Ka8PBn1ra9GpbPn7bEYpHeX5dzfatEqLCtfISzMzgmARu5j5Tz3ZQVHv0I6Em/k1IJpnIsFYglr2
oCTXzqlqRh8seH5hqXQ+gXDQhR1ZGw8mSqoUgHRLMoOm0p+1bnPTkHGKS/lEHcBcphRFs+K4Rkbg
Y+FLTkHAG55GXZ+acHVxeI94hNktstS3kgGptTAacHf7z/Eg+qsqBbBYQDFoKaRJ+G1tUIFKyap1
xBg4bLNhAy1QzTBz4YHhiS/olJmKuHcIUd0TFOpr6Fih61n9K4lYGLjxJxHXLa03xHYsnHv47hR8
2yVPs6V2guARIPpjZ4S5ds38fJlBYsRUlUpRN05apBPJWyP8521y54q1dGy5EtZSTBXLKn9cxpIp
G7mREnsrzWzOBevVwuYiQD/FzzKZtNSfPSUNm1Tb5Ntken6Rdekf89KSZKy2HEZr+ywi2edV8Cig
VT6vDug+BJM8U+aWBKo8R3diXgFuPh9HaamjqtHtTeU/eM9H/QInWOrrwOpaBPLbrtRv2+iQS/+j
8Qkpujy7dPmz5XIT3dCP+INVjkZgN7vG3Up/NjpFeoBAczvjjdNKER/6p3gAu5wMz1wut1YgQE70
m9KXUr/CXQ1mNkkjzgA8tz9QX6Z73nl3GPdDlR47CowDBHcfk35M4Hy2HwTkpRbW6YlbCe2425WI
ooxn17X6zy2wyrjuKVtugseji5att/Akv4oe7+L0C0lCBnTf8km3/1Vwpdop3C4vbDJnolcqs9P0
nAsyQY870Iznk4KCV8kQH57N+yqDLFf/DytfddKngwjDukoN4wD1cAgBZpQ7wCgWsksdYSAU3XVq
b3bcxUH91eDpHnxqQSSTqLZuyJXDDTIaPedVqisFJOmb5Rb4VSQOrR58vpHmnjAu3YV+Gby+UfmO
douvS4etCUyzkIkLs+HOFiX62xMItTugqvmeX4fL7JsfF78avt8CdEyanEi92V3NWTApWehjO24J
wEEvbYX2Q6TUzriWB4YLzBEYRBLxlYQbYckLUym3U9fWIgAJ0e9jwMPaVCoohFmCcph1lLwj1XhE
MOCR5m/rX9o1qfdWjdkSwLm/EwoaV386hCoGlMhmHoQ874A3ybCI2DMl74upXfO79SEtgCjmtW48
jx3dsgzoOmeF4iEqBWjak+zJucvHSCUXvda3VyBZSKN4Q9Q9peadCwAem2q+9dMcT0rmvU+v2T9D
qSgdOsGWeawxkhSqJQge9LflyWRoQWbO23nfb/XKuiBKb13qR08pWLEIDR/2KJrTfvggYx9qQSxT
fMLTfwbE0dCzr1soW+2pVB+8wyf0lQBXSJxhdDIXWiDbTJ+aThTtIVTvaBZIX23zrLLU2u+4s8RK
6GxofsXUYl5Ls7sK/KGOZe+rQLUOEqWBdVsxgVIG4kQizer6rH2vLN4MQuj1SDBVhwSclg10658m
LE2S/M53ZqRG2XNqieJsXHnJbpWR6KlVU2bJwGYBZ5J0ZMfYQ8WHw6/sduPqxBYRexolZdu8v2vQ
tvZ+nPCYJvV+DVhXZEB9ua5XzmBo8eIe6BT20Yieai84Boinunc6SzWUtfpZGHl5CdF553l1z80W
J62c7FQyeohoCry0qSmBXiDBvp6cqiyhQrqDXvRNAU7xnJnrpFyh6GQ29jcqtIx5XDBPDBhWGQXs
hcB4pJ65a1A2uoH/oeRFs65wFC4RSnYLM4JZIPNvn//6uadWn0u01NCa4aFHBVMOtpTT/lDs6kuG
7dcKyuwfwCWnIM1+JpcdXM5/uakJtACQoB9Mkml2Ieuw8S+XHvZKIG8uhwVz4JGnr6pwfYoHr6ae
cd6gvhiGoJK1YEMehAgDcLv/yoIN5C7+sfYW+9DT7FQB6d9ZRfdQISxU9ZFyeN6Jy1CrOYkjoy//
LD1NEWVeUzinIJiwCZw47ETJHXMqtYnqwh5rYoK0F+l/a8V2O6iFfkGpfoighFbBJl8ZcB3GWnUx
5bG9MRpeJPwdllb5UW/XunLNSBL1ZKW4bPZaPtePUPl8LvK3RRwSTcNTTLETUh0WbE8KlsZdMAsW
8zTqw8rW0Ky7BKS596KtXc23kvNYleOYfqOUT9+4eFjv842Oe5Xt6jQ8HGQfShcsvVwJTiSrjg1R
JxHgpYJ0TJnybQuGAtXMtcN9WznHG1ezQHej5fyGnWg9ni7tqyUIJ/Y6nRasKUYB28ahj09dEk5S
u+4sNbfwJcH2F8/hWGqIEHDRbgvH7fEB7r9R3qBhjvX793DRQ6JnH/36wV/M0katCBYoYK2e/nbO
pGoVtCyflBgDjPz+j7nlCRH8ZlLadnz6TtHrw0gvYtERusI8Rmd3beUA+HGJ+ukFk9p/gytcTicb
EjtVpE6DqdRiZ8RBsyFAZZSHfO2MfL8phthEYbhpO5gr6GCif/dPEjvX5N1SH1GTbJ5rye/Qavtl
z5nwqAN8hlEFX2CuJqpGzWZMqIQrTRd2gI8wgPVUNxMTsuCjIEz9p2OYOZNEgC/99AwxSl4EzDPq
Y1QOitZG89pYBONE2Su5SQN4Qy9rl37choOXKgxwB3Hqo/tiCn9ybJmIk9BAwk7Lwpxb8vuW7ibR
YOULILJ/+IRNtvkxelewIXt2fJf3W6zJk2bpmygNqsWICG5DkfIucx/bNN8zuG2WhCG+RkdOp0E2
3pB+z8rGD0IKen2scnPge97Ww5p+8F4n5VQX6wLbM8VN18ZC7dMrgWbg5EG2rtMaCcMW7Qp4pJDU
Lb60ZXTvVG6iUpnGMeOUIFwzSLhFmOuqaSMq7wFqCeaviOh6KWnqId4pu6+KX95nfUmB9swBo/KS
lgcC7u9a4j/duj/jNbkrpnDYeHhFfFznL4MD56kzwl8+hxflxzCZ2uGU4I2Gfz7MU6xFax3tGW3l
R0tXsYASzkYuwiOO+yT+fU3EGzhGwP0qKJrKpkvonmsmjH3nKTWa6u0Yv4o0nhfCMh0EZ590l3QY
rHtbYpS/9WY7PsrnZxDgutqqEhJFWCN3FigUvfKeLlKO1Y8efySddZgKHeczphCDl0y4HzCailPk
mKYXTS5cSHIZkKuWb8ANk+aX9tweJMaMATpO2P1sulRkfpdCiYQuUjPDC7DeCxYq81wH80gfwWAn
9uJ6xcw6RM200tDcBjA6PtLseRMdwdvVVZvYd4s5BJG+WEyMY4xoBRSmbeWmbewQ3z16J/TQMDy5
snEaphA3NasepUVDDEfk/v51h41VSNAoCy28Jk/9fwOFSZAikVCXXNGz2JEO4Coj3ubFLMb/aYiy
a/U6HE5x9tW79ghNjVqVQ2zn1m4GsgPk0Yrz3B6a7d/N6uMTD+MrCKsFmC6/sC7KfcQSzjp/xYsW
shhd5bzcoPVttoTsWmxrpXKbPk2J1VJuiINy/wXojIujY2U8gg3sPaX3dgxIF326a3SXW3xA5DCW
Sn2qBakXHrq+yE0ApKwu9DqPKkcaSbUNIJUZzEG+jCTI0wsic20bkAwgN8xNUe+fIGrMp87bF7o8
VjqETHx0KPtRe3D29vXYT1vOY5TJDQM6y8epLfIhlXRBHK4Z2jKZu2POEBLbA3NFlPIhTKJQC/8p
a3VLUtg39ioCF5fXdYJAPopGqBgMDuJt5ODI5EoXi9F7JDAK1RYhLHSomKoE63YCb+hT50GabjIn
HyUbnaXYppHs10QrfE1NBbcphdLRmaSd77GeZw7FrusTzVRwlKWiqLaq7oa315v28/o+bg5yTBvb
vYZ3BK0myWX1Ba2c6nAQuQ3xLpFurNAClr9wAWo8HVgETmDvFlMxgy1XduTQyxgpfkkEFF3yXQ2J
pPVXU3nq0Kt2ljfvpBXrd8ClIYAija0lCF1sjwjdgXaEe3oCeS86FgeBmvhgDutR8rqOxouP01TZ
qzK+Gp/b2KQAf9kJLGEd9VmFSszWxQQ/zjpLypwMSl2+CLt5SSodcxlxCKTWl9NFYjUBRWY7s71R
LqGQ3XDnvDgpHf4q0NPfrqwdiRcVHnVdWPikgFti9SyXtThx3b+LrEOFVNSLy1DaTPTuq/JmAIPw
xEPxQp+MZeqZ++u5YFwj1HK4ofd2j9hKJbECXp/WUdVXtdRv4+++5zdsFyVKoSofaTegJ8mvJmCI
0GgZIKjN+afX95TRrHutsXpv9JtFTYajLLY3fVwkHcVER5CD4/lWP0Fhpp/V0JEkWeCvixBAhaYC
rHGRub5/o9SHY7nhTMlVm31NmO1bc0brUxoiz2Bx6dhcGONjPx9fc7UfDVWTmGg6INJ3b8Mf4CpU
zgmrW9Plu0GNoQi9MApDfxdGDH7nUDn7xNc7CZ6G54UCq+igD9B3qwglIFh9u65YYFgGVIG3MmiS
IlVkx99xCzMGWgWWQrsOpWCEPfR+Ui4HQJy4k3ZwsoeznmcpBc49bhjA8xpEcO/ij5DEJpDCV8u2
RJbpqjiHcJW/kQgl27HqwkibNxCid8bl1hTNxTgmZBF+CNt8SroQFRSeAdDmTk3CxUxyqL9H84Xh
DCGvHrvCbSy4CrpH4kMiVIJ2/gOm5Kt2LQzWJmx3FQP8YJOGVAebcvxUKkUjpKziZgE13ZOWWVuJ
s0ud0mmYlz41jRNx/TGujZfxk/sf2SqfRTPFa3ie5OCXXNSgsRqh/TngZMhDN1UYvFZ4yWhaJvnJ
nkPp5tk3bfWQJoFqwMkk4d15DegW8HcDTy+xnODYypOVKM+Os6uUhymCIjJ+g4bSydZCol/0E/DQ
aidHqjcJInzwm1Pnc7ooC+mcRVTS4+jxv9TGoZavgCSvrcdo7MkIGPGlOb2pjmGH0ZRQ1ON1A0Mr
SIDK4DLQhxljxd/Khcj4PEA10BtSHjWym748TnhibcaGj5hxBQ/TDEn2XrDRQl/tAmbJBUBNOg62
rToh2dWKc8i9Lbl+KWkTXt+mIBvbDyA3QsPaVcKckCwS4pHqDiAxLvshUCQc5fcMz0W9XIKaqk30
xY20XpM2hGJ8MJKgHHjLAo2ScVbhiRcyZakg0MeuXFhvrLlH6ykYHK1kQn4cBZTu3+whDvgshytp
Bc/dtCXlc3R6hRiXv75glpB5e70v6lL5kcKuBXyfnMSpje+POsTeRsrRt9Bc0I0JIzbkCTM54qTW
HpgiiveVxQbKU+mKezRrulRAwCC5xi/Cq2kBCN+Uqq72D8lNzows9faUgyXDMR9XAJmr0MWFtrxR
rvLF4D5k1dqGbSp+ox6gBqFq9+v0NEc8JZgUbOJqQUG6FmmOU65p6dpmLCkwPnSVcWA7EFIAFnYO
7KpjHlcfxd8N6/10LbjIDLe5ACxrDQSv0XSPH5YjjsQoGoEPu5jcE1tUbmJmwpjFcJUMyE+354Ph
KBE1rmpY1HULyOqUfDIC9bNVcSBjbWV0ZVoWGOKUAf9v31YHhEDA6HgjL30rrsLHOLzVcqlxpNnF
XSRp9sNMj2NhOouErSjbVzHcWCIIJNgpsalN3vm217HgQum50XeMUN6hbaCe55ny/0oUjMNqCzR+
ZdOCn15BVGV7+x92HwQpPPpGxmrDm7EgUk83N9QNG8sxSF4upjrcOYTdfmOaxoKxK2yZUhvaDXqI
gkn3ak9149A8geuKn3L4/2Vi9nGgwfXwrl90q4KJ2LiVsm04r3Y5xvCR2BPMkEqLJzdTVmNN9o++
JeBRVUmHtXC6Dje3wt2g8RKZ7ixCBZfTLWA8cbhQttsEy/WVUS1URwad4NBSYwFtretXBrFCo/cW
0PSxr2f17w1+NtrQLX1xELMBTi2LKRMEvvwJw1QT2YET+VVjZ8jIygFKVrTTLSCfM+REguz54Xge
uXNrSFKt6otOK7UsYhVum/uL+9USr1GbVumTUhFKqN3nbulzeFhyLx/5EVGYZ3aTpjO5fN8JDajy
+3HS4XF/Pu6UMlZ32XmuE3yNOZ0eEm14OfEfSompLwNsmKOI6uCDc7Ppb1s2+2J2iTjn3nEWEsFG
2NyUEkhy2/GI70fxj6KY2wlGqu79Qp7kBkcRuB9vxS0+ZP620vflpVIZLVnHzJ82zpPC/Z9Y0qJk
4L0Udu2h2yO3Xh1jSgUoB6LbZXQnsCpr8MUgwrXuIWPIyOUaH4RxvO1m279F4i5Ut+sNhxNWZRYh
L9XH1BfL1DDaSQBGv8lbRF/xRDqPGozlvB75XdUcBzqozyG+c65duXqu/Z01+2q24RjoqgIfSuAE
bFbZfjMhhxEiA0vIaZG+OcsPsgbmwARSVLWOyGZClPCQx+EfsG2Xq1IKQynCvRCVHxiAa8koY/el
GnBijB31QlggpHDWavKTCgTXrw2GXZMRx0wPI7Ao1APfqqV05TuCAxj75gY0jkPvC8Q7id+UggHv
fyH514xqavaQxiUakjCLz4dSufQ2scKK/9wKiou+onCrKlp3i3eRfx1HF0gbjz9KpQtt3jCwmZFU
2f4CcV7paGkQTLe5qPh5JdExDd+BXJ3P3toX7raRh6/FmJkoUiyvIqwS/qlLT5veW/yP7XY/A/aS
vBwpc+gJVmPa7yEPVZ/zXlM1FARNrHO3akCfsL+rFQddVC9MxIqf/DO7ziymla/r67R2ydSVw/AR
eRltc/ALZ30dRW3PFBIDB3DIsTl6yKb2zN7LjYeMcQQYFxduHXCvovd2x4nYJREXg+YlgGWOmZ86
jQsJ0BxBwwtURHd+Vxjd4vpsQFlYxwWSAQ96TqhOOvfiv5MekVHg/S8qMFK4OdagjXgWfITtU+Fj
2M2wPJ8hq31ebercpvSvFgB5oXJUE5JutkPJb1XnoBU8nQcCTPhxPwJQ+/1Wox6KGlBH9kQVbldh
242/nKhuY1jqzFjNjfSkWLvawtQh+mJsL39Dh6KxPYdHeLGwdlwdOfdfvcUhwb2IJOWhM3kNxQMw
9tSrFB9KJ3DhYoXdlJNIXnMFwUD1NsLOub3gegD6+2eQ2sjwK3KdO1ZdkcBfySYRzjEqQJvj+VhF
7WFVvQ3nqZY+YR1NFb3CUkaP80G4qKe1RJvV00OUeiQ53qOqQrwR6vrc+31TeuomlB/zgrmy+I+6
3Vk2oMJ37neAhvAdaRgOIxdfZnT313IJqXeinr85l2KhU4odGksS6KlQJ1KT+N8UkEiJo5YuBAGu
4V10EGTUSoJkhaVIG+7mtUEfaoezPSuc49wFFyErpkywvSMzhg9SLEbaBUk7oGVySaT2wyyCy8Ik
3AoRUZ6RJCA1rQWxI4wL4tqKsfW3IsE3r42m7TTZ7YtIs2SISFgScrzDsRPMqmmc4eAwShute/PT
X/4svRnHiJCv4dd3iypWnAEXU92IFl6EtNEzgp0jDYpdB0nzEA6J63vyplBQPRHcyvegdoc6Wavi
WfI1gMIdUYi8wVczxjQ0MutnnycnVekiKGU6B6IVLiuvHqxY/zZAXkT5nfILn/0Q1Uw1L4BpGi7E
/cqGsxldu18ADgYZSABcsOm0kPf7UaCNpETyi4i+mtFu+r+tlzeRNTts02kAW2V3HhV/QhE0UIdc
1f2/f5+KBkSfMKLURNJ3sUdYVHDvsI0TG4JZqk+Nuzie6HjBDM5APfyArkWlNSFdmaM8vNz3ZHpx
PYKL15dquxyVdpaZv1Fhrzb0tm2ZDHJZ/tuQZxfpGb4nkS6daQxEMIqr1J+MtGVTeql5Fh7V+voN
qg7TYo/025ldyxNJ6YpAHjBPDKPkkAhFCPIe66zfmRC/4nzQBXLG9FOar0zQCMU16k7Ewn7aqNZf
bzIDjkdh9PbDnEJev7qDGw3CcGsMITOZpz/kbUwOS79sJ4tWJ6JNXtMJ+51nHKrx7kxq0xS8wjpX
nqQlZy6Jjtny9kK0e9O7vLy/m+FjpdRXVn5OqPA3YIsqkz8tbiCCJ+JCC8wGuLFhv1wLvPyuho4D
ooaDz3EHFdjdLR+bHPvVH32yNjVStxqyN3M5Ffox7I4aXckiZHS2vozbFjtgWq26skawHfso/58Q
K+8lo30hD7YCMBadJKxt0xLly+MlF7yb+aMrlRft6i7l+ETSTmv43QxLunaTfNiKy7r2htPxIPPR
15uehlfDK53EUbzwyeFMaO2IwXgd959BjPTBANDJPZTZNxA3G2mKszSZuCY5u2/9IVLplNx+rQbi
09HZL0bLGCQe4QYZaBVdDbZbNtO0vK8zjH35l8SfdylNQVNNX8fqm1SJg0ziwGyW3GIZH1EohZm+
j8w+4AiVec+stHW4nfoBHw7ujt9nJmQmzl3f4Ok6WpZqm9MkYQBqEj5w/nc+X2dhvIAbu40rFBs1
R5r8qTICxO5M3zS1Ze+g03VB/iHkurv2Yq5sOaoZr9FHXUxpBnumMwmZeE6mdZU0lLGwpl60JMWw
hp3cWwEOtMy+cuBIDSrTCc0EomjXc8/nQEEC/wzG7Mt6ozHCGU+w01PjgzbnU9ula+b38ixWkOAG
pR5/rOauRYVZry5ZQ8afZClK6Re+bpQtQMB6ZMWY13MXEldSSABwF5+lbsJDsY+sxoxmbrOPU+DZ
jepX4dfLwp5aJHCfKhnDCH6Bu+Q5ol+V18cEjECjmZvrE81VN3EOp4xtxqLUThYKrZgbj/AVeVjc
HFawrWVTej190wEip5va2BbyLmltXgkAF9EZVwr/m6FWmZro37FIuFYcJGVAevCWosGg1BDjvlLN
IvQcDGLvUE6vBnMOLygsYy4KCQB2Osu9GnLEEmRmrB+U1arVTyYY1/9yZHql+hyAtssj3v7y8CHX
V2eRXxptr1Awc4ZlpXGERlAALsomHiDV8i1x7UNZ3OX2106dMj1k0THLsuA+DrI8p93iIboZxPBr
4NU9wX/GQUo5EK1vP82uUplRW1h8osrUgTtKhuE99jy1wkdV7TVqacwAm94kQgPaiWtYOaHGdndM
oVoR0T+eLlA0PfX+0wvoajt2425L4E9t0xcQ9KtuJU/3DKn97zOzBWaRJhs7jcH9U89x70OGlOSD
fafrDQatV/WqwTTO9vUMHZvIiWX9Lj6EiEO8sM1HoA8KAoEtmHRF+YcuJeWbsTod3ypRm0QCCRnH
7H9eSic48n7ODF1Q/SdA6wxF8DKc29BqOG407kDp385Pvglz3ooJ+3HSCdq3EzfrFGwHizDrhaBJ
yGJRK4Np6mIyUwdPwLaI8Pzsz+dmVn6yFCeNUH2GR9mP4JMRH975GQSCd+pEc9e1G0Hw24rkx7X8
CktU1jZQ/5Fl3IEMzGNQrZ4QPI3mAaoBIwKKs/0Otp5uEgNvqc8lOghrzzAM/LxlH6Y+NDd22W3J
KHV4Ix7yKbBtUr5uvKGaiPe4eB2dZvjAa2H0oUudoypiSVVPw0d7eS+Xg2Ra6pLqhgd5S95ly61o
+wewz4eEUwPiNZ0QDYNz+kAApvqu4QpTZxmLdaOBnYtQeGzsAb2Tn4C2Xak4ky9IFBAjiME7+MwL
3jMqmNHjStxnKiNSUu42G7Ew4h+RyXtWNVETz2xTtAzkweHAp1T8yT+8fLTI/0lhCNdC8LZiffS+
usIE+aznHhgLC2HDYg4Y9WJBq/RFqRi6wb6xTjNjknKyYhP1ync/dzaBoGb6ECnd4h7NvoS+wtWD
GgedwfBzSqdLqH+YqlzA/CvTG82M2vDYByJ3FKXV+lsos7dj4bBa/wGnvI46AXXZZ4g0rT2H2/8s
J8oD/FCuVIOukrfPhnDc0auyOKBimSKyn36RKE38/AA+8ISDqNH/VbN4lmQNrQrGCwrO2BYXycgr
NEUtpwLdG6qDy0UaqK4m4Lhd4tsG+epFBJEA9RqO2DGv+txN1w0Lz/JAPvncgaovdoymfCWbyl16
PoBW1+EpR66LdD1F7lZO+VtLsbwzVTf+0WkjHT1BJRmu5L1OGRnAMYt0EhNkjGZKB51Aww1bIpxM
HzWAbUxtcZg9xcx0BQAi2Od1tqHEUOBsE+fY90UYhXHw1J1Tq4eYCPG46F9QguSFqQ/9cV6QMQcl
U//sITzKDG42uEoJpT2QTlFVzvkGP+bdvpLQt3kBdOmNplj27PC3BCT85AQNtHlOu54Xq7Hc3Wp6
tqeam8nSX+xJMTMQNkfxUvW3g+oMrev9gikCQwkb1/f78zsj0+cyX6GTt5BCco+ksNhbEy2ZUK4P
kK8iAIX/wvY5h/Y92NgRMOtk7Hw6WFz0+ZIpQUWe5574irAF2BC/NenpIZVvUpVBuSHd+uu27oly
El03yggvj7iAREHAn5ePK0gRwDqdL8yXbtPbhTa16l3xWTTBnPXxcLnGKZBUzlUwlDf4DmydaddW
jAknkyQV+muYCoN5w6/fuCj1m//YFVLhWbFrrVEh1CBdAEqIaoE4DCB+cbRh2kr8PYzrEhxVQi/u
iXV/PPdT/RDgryufHsta5qtLlWq7mqJHG7DV01ROCAqrz3LDLEtzu5H9T0MWWGqJNRUsB+13t589
buvgp28otDJRZR5fS9aekj0q8E/smVBnLdnJbXCRVJAeJSP/Cnmehk9ZaHP65j75In0Pg2Qsgcrm
1wKidKuPC3Fsfi7CeGw/7XCfCuGWbOMpF0TL5Y/7oCRqsypiQ9Pvzk9ZbnL0auP/hhnq7BURNZYY
hpIzSqZC6gv/B9AuB9aApPF8SRXSbVe9gQuZvXx4pYh7BtZidai93UYsdG2jhGm7Bs3J/RhcGgbg
bbhU85QO6qhSFEGppZq3C153Mzv8H+iBgDHsyOBa9ssqSO/R7xZRGeH3PIjOWaQF1MkR5p0FkB4s
xqNyku30Wgugf1Dzxg4LfHa+VQEKQsXBDXhoGti/R4z22rxIiMdH1i1p3XSE/BLMELMuFmpU+mJd
Qg3wnF7GFc3ebDbtsfZ7ZXwmLPMnooZwWrJe/Sx6+j0CYbVedGFhYqKnlpRX5cXx6uUe5CN8fvOj
qNcQlIqIuK8z9tHkbgJPD0jhiwg6VHXV6N3HI7iyJPKTQJzG6oWL3ujGDCcaK0qxY3fup57+QVZ1
9coDdwnvRNxwCVUfuiH5Us4OQI+mHVQAQDWHeWAef0FEK52xRoZUzb0DtQCoAXKNfBVzw+XquumG
R7FpnavQfq1yVIPLsPDGgDryEjRc6MSBw6tulFYyTNwzsQWhKgg4DO/Ct3FPXHFqzQRLNLbR1v/F
DBGUGqQc0K0o1zaF9o2mBAyYHo1/QGdM8gMQrIq4Y4gk7borJjsOuX6mE4FIQ8uH3o/vILRSmhRi
Ldgd9SdvYxLn5OlYjIQLmxc57BBeQ6vm4gGQkg1EFUIzucsJGWDyYI3ES7771vaRyyKpaiUR+5I+
LdBhE4bf0+kYBBQXtKBFImqFTeolqHVewApw/nfKRb2TInoNQR9yE4kSIvrpC28n73yEjp50d+EL
EMt3ae1r0tVA53/Po0PMKu7boMZ31eV4pOAJyEOB07A+Cp7i4PPoGzXEIl0qoKLZuEfFoUC5CySR
esLS57BOdIFWy1kCUdgo7fh9aZVllzutEVmi/M7VmO9GgWNjHUlM5VX8Tuf7RL9oxsKUoIA8AkI2
8pjed6vFlKxSgc+wmyNKr0MZKLd/G9EBjQyyxqnrSm8pBD2lOfCAWxKfnXkLcO4OXaBwQgQbwGSP
3NgrpVFcqQ0niRJ2rNy0LcfYPRLg2nD2qww1sfcr4xDtYB+1yqCv1yPjdPlliFTbb/bhkbIFJezn
ch0H/EuxLGPwm4kbsy+fVP3p8P2u+E72u5+cXEGE6XBpdFCWA5tBnxDtB+vor5hLedMfXgeBZZNO
Rl8uGzhi5D/UQFmUXNvdH1S04ZFcx9nB0Ph2tPFRabyBvG3kxGl5xEVJhdmPuTngSBZJ3VL9twZk
hi8EqPkzr/FQR7AysppmsqaP2xWVPRe1X6tAAlL5bkG2H++wVCtGt5ZuXZXR9IK5TdVXMpfGGWyD
61N10YMmXd1iN/Gq6lckGYpLOVIO4lRfxInc1KULBQ9CsXmz0mjz5s1GM+/lLzwYvR2vSqpq8G2H
du2D1GnVwQ/apP1Ds10j+mOJuydJD0fNkq3scTQwU/vHX7TwdFN/Br+eGBQ5gZkNQrzFZrX3tkHe
wVC0N4OBPHizuQ/g0LbwogsPg+mb9S11sd9M0cvWfoaYeCT3nj7KxJJenlX54odjSrfaFu+gLH5L
ohmOpx8wfXPVSmaxeWcNE9UWssgzuXAjJ5Hq8KIF7lXaf0WH5l86gowUDPGXtFDb86R8qBGUZhEB
g1Q6GyAGP+LHcNepWRqialxGC3E5/hE8EoW7yphLZp/mW3qGV4qeaGO729WxKyA09bDa8LZK35VI
A+XxRtaJ/E7jCYIxJHT+AxIeIsfEuVESz7yPKEUxapnIkMVZjtbpfU4rpW3TW5qa9wSFpgJ1ZZ/3
Ir9m9zZZiCucyL1kqEYRa5KHBDl3cV1PkFMUNDEZmug0fVpZMetq8leq/05R/BN71Fd1j6ARza+O
cHKKkjVAT7t1ilwGf9mBIBx9TpZ470p7Vvm7kRyumqsu+ErsbZi9hIY51lKjTzWu6SsZTXYxWMN1
v0IzpebnO2uPttqqHlaBdVAltISvNUzogi5rJW6YmJ/ScQT12o8VUuLMiSqQdsUXfhNi+zWl9Fo2
93zclBCebGH5FQR675H8P+ocrYjykjbqjXQ+UMDyzSHYc7EYUa7Z4K/jPvr1jF+WH7etIcL/QRsY
qmnU+ZWOjMfyps9NU1UlfMGJJD+qlhA8Nf/nz/jnEU7VYT4jMaC+1pCBjt8jhqjNvmGgD2UMhdCu
LAzF+h+3cHIkre6XAj8MYb6y+xhA+vBzf5yC3HAgaW9iQgNQkm8E6AP+gVSaQWp2CKcxGZvtwJTz
NzH72jn0pJpcuBYN7zHqxQQp11hP9ADgXLou2w9QpoVdilSlQeShM9qD9johe8ZKBSRgao1qtHG9
Fdx4aK+eJ+IZgv1Vxh0WlVdM54JhLXb7G8vsybMHfsNiQWsgZO3yEvRqpV66sMScDzkVOhxcaOvu
vOM6ScSxr4TDdbve3zyYyHazOIcLSGFfRh5fZyHdT6/JDH3hDWNUZqLrZQoUBk7v6HmCTWW7Zjb7
5CwRE90oNrHkdNT5uWwZGO1yVM82As0YiXSSlw7nBUHQZxgJdzUD7Mrx1g/GEf3nuYNz1GRnt1tm
J/zT7TzmFh0HkkqwZoqX341H9u9Ylwvko9QvYxNdvPEkLhipBuQzhV0TxfRWkCuFnw2TKTkFQaja
mSQKKz7lzqr36y4+1LFkcMiltaZlLXJJKmcYnO34IH5EuKnFA1AbVMpUb2NUaXR5O+9BhgxI17I5
h+tfhQ4xO724XnT0GSJ+SdztLBLzADhj+t9+PPsyAXOrP4SNe/tXbXQiqfhf4laLALDkZpQyVQk7
jZlyzfr3EmnN0Z2n0ZQiYstd8CO6pX8F5BwR37ay/IBSkt1lb/jLTRmjH+FPJJQJF5ZnjgsxLj7h
d6ujCxiMObZfh8KjKI7j2n7OuIKUNBJqJAKOlRuo/fLvqbUFdBIxDO/SMOdrJsuZLmoSp8PwAUpR
oEMipMnWPcoPCCV5YmPBY5BjAcH5qc7qhM4dD0fz2WlROo5C1oa3sl1VCaCKDTmQ/+pi2S/oTZki
7jg6qKwY2i1DE4rlxdb708nT1Ag2AH1GMcHE1kL5J/MU4re7KnoFj/QA7UthkZxYRvohRP7eW+Pk
A/KypvGHYSKG+t6kGsU5LHgzUE+SgtyWZ+PayN1TakIVsTKQvu4zVaOvm2RXJLulsmj63zYossmV
JSLFnkbvFxOAZfM0AsCoVVFXtehkQOfCo1YCxQ3Gp07wYNwKRnM1iNMerzKIM282dfaFZ2CO1MZH
lmVGcNvOKGF56jSY9r5ZRgRXFkJ7QOzwTQi5i9fWzlM02dXfIVSf+dS6OsOwjgT7mu/nbg9h3Icn
hZT808TvVynFj4CAcsWT1rT6PAwtHVQymj4HtYfKUaHPx/viZ9klmnXG6TjDGlfcPH6CxueZ/gLG
KGtS/JqfMv/0KcDlGQ+YYa+rUWbj4NXTvdqkLnUsMBu8qQqaXr+DG4wMRKUebw8a6dCxQIjBL/nq
xSvzrYbe3mIV2XWolXLJeuzMSpBebB5VWyULnlesXTNf9jpnjfxREYGRWQ/B0xAqndOQyuj8n7aQ
Kaxa81LmJESfH6MRf0hyrch34lIGvDo1wByoP9Gs92Vz+L5Z83aUIK8MarFkLDkmMjcvZShFxC+d
bvPOo1/MnKSWh/rtBIDCbbFYKsxyQiCameA++deFCm4eUm2pEkWnRf2EIgmPWQ8w7+JS3ZDjcPeR
uEqwdjburuuKWBzW584IeOKcR0bdM1GoMxSI29UB8ESo/BCYlKlbKnEscWwrQdkbtHN3wWfDSGZ0
sITMR9SQJTm9yJOsy/SOi6FglbrmQzgPHHZAQ72KR+3fpZIJ5LNEUK7gO2yC6kH5uMnwIhffm2JX
JUQAi1eDUefiV5p0DPXhKBYUD1vFHMO4ADbOJBv071wD0eXEb3wjwKJks/NUJyB5AXP1zVTherCv
j0gFH4o3ihKOBqU5Frjcp96jS7MiV1fdu5qNamUaIU3OqVpldB8E2qu9wM/a7V20fBb7GVC2X4gQ
YkGmLPVgh0Ktzox1SIvHANnfh1FNKPDNtZXi43p0S2IGKpi1tdJnQVpqgT60WzKCeIeBbgs6BfIT
CBRRk2NE4qYYdT1V4W9oVTnuAUxW5vbgfGGmrT/fgDViH85PJc75PmARCp+sKW4fO3h/872FZyE6
ei0e7GqLgoqjpBdZZDjjT5ZcPseoV9cZOCza4vH+j2qWTfSxKvo74iavBDlLHleHzCsPxBEsqu25
JPl0kj5qZ8jFde5L4GXu6hW6gUDgRIpK3YMciiMLFQ2ZgseDFlo6dLVz9XzpIMWW5AvJsMKnI1R+
KJ/B2XUKl2132HZ8fjdkTHr/IcRvlF7LlBD1wBIWnFrSwpDgJfcdlStiKmDDRvmezmSL9SjO4vaz
xk+KJFPBQlsO7JAcqXf0qpSTby31+9vvvW5RR1m5rlkd396r79K+p991ApB0PT5/mCxEPJjGy9Ra
ljosziTi5hgu6IdGiltMXzfg7szVdR1FCMcaSgBzmJfrB96VaVEV23bUgIPs6a/d8ll5LN9IrkfB
3DXTtycvGjTFo/ZysOaJgr9QS5WI2oBDDf8+pGhbiBFTyaqRSFso9BvgFz3LHwAabuWYRUzbUtVI
Jek7PV78gAqJ6N+mfywG/HivMePle5ijJ7qlKT+VrU/gTLLoH1eVYLzGTqGozjELZd2bKuM6JJq3
kiAacErn5cEZhOjEMor/FoxWL7LzUAgmxXglcFPzFxjJQsZqF6r/dViNlYTOJsSuKtAX6x8Cx7tw
HujJ77XjOFuXe2yfzS8JRNTF3M7iGA2wkeyVd84yXi1pYzWlEV9/6JpHpBGEoxfabbiFhLra3K45
EYZcRvaQGFvy8ZuOPq75dK3uAYP11juSwO8+wP0Ai2XCGKt1eRL+wjO10PExqWaE1B6Q3a+J15Lp
cu1clN6oL+ULHL6QBVuIhX7HoCa4tqtUfzhIjwT6438EeBr/ffBQamQWvxt5oXooYIca+pmcQ4Dg
XkD7wN1ASfCypeJXpjirSinG1PKL870iXtk3JPeunCkwnQdoF7BPMWMmqkUiF2+A3Mw6jXQzgB/G
Ze1dvCxFKedO3oofux61cdbAGzad8BNxJAbDNt5LoP93m01RsD+oM4KvQaOyHQtGt6oMmghiqoRA
vZuJQW1ztQXZoR8aa2e/XgO/gzHJaOhlo0QcE66JhaTi/qB5iVoGJx+oOA7MvaxzT7sIgCpv6ria
VW4F8/mnl/lB8Gmu9WXXTgN7sPjLhHKV6UsMqUyz5EoklS4ebOuvso3951q4jWIMEp5WbfI7u/ke
sqLFjlvUL6TwY7BTwRfIj2+qmsHuC0kCFN/JyTP4szafUqQEehn5Vb/BqAVu9qvNtJzqiwxmKldV
H040rQJDrv3nnBHxQdjKp1yrAmcHVoBFoQ71jHTVshbHJ8Mz3AG6NPASk0Dv3Gfbn5hBZrmwm6kZ
i6eN3ZqkAbPyyj5phWRZF3WwwTzJGYKaQLJ+CxxXECoXkKNhAmRgmDDp9Oq4rj7q024+gkI2mORX
ww1esGLMGWBC5eoYsAybfDDe1JYIHXa+gWlCnp8Ud4TjwsDfBAzGFOrWc0JYvUmbcByfQyfoW5Q6
MwlJxrjmeOdtAvEhF+kllP5KgPRPhq1WGnnhs7rE1Ae0OcOy5YcOsG1L71QMM6Fb1z0WZyecJwgD
rgIANaBrS2F8sR0tMX4FboesgkCZGBknbSDoUkbPzsDU5FesOXju5P+okttq8GLNY223eOh/C/xB
tIARJjEmZhVenobnn9jtAPvwitYqG72pOnoVHNO3RZk+ZL5K689ss8LriyXzdyTDF0HfoUV9kqKF
K0jMl/eIa3HlkZ/seVYTj2MuKCJsK6DYU6qBEODgtMAZ5Fpbih9z7wB3AdYtjOKH9NrasZHg0lCm
Ync/GzpHT4oCVmGOtVJIiOZDr0jbfYNnBj8BFjIKbmabP3UYfoYfSBgdeDlLRGsoDCFwQ8H5pCah
46wFQZtiI1D+et0PnNq6ptZpqpnai/iyOKspyJqqM3Bq+i5I/eE+797eIIGUgAncJ1/BucQXiCKY
5Mc9BR9gXFOoBkaKYBiQZBJulB1YGaNsX58VHsdHki2gO7XYR/tqAZ+MaKQOLkg23102pIPyZfNR
iltaMgCc1N7sH4SSgTd4ERgHuw9dk4+8jD67tI/xYfzdTF/LszWpTwf8b5uOChpDdVl/Z017uct+
J+kRj1TzAhD8bFh6EgEjL48Ja4Tot/QYAtJBIi+OQJIEf9v9L5Ovk+dNTpRJGLbgaXxLQqJKqX+L
fBgl4YVf0gxOvSQeRtfkkE0xkWgf2ll4PiDUvkCqRSQ8fC4/HR7qzxMfD9xTH7GxPx1TE79BQ1mf
Dd8vNoi1L4hPqkcaqWpRRP/XLMtMlOoQVrbaCP4mbatOomwtN4Bez7AO7YFwlZiJhsqP9/IjotLS
GHP64ek40idwz9lYvkPEAUW5svwvJg7IGkrQkRjBeekeKG4Mm98Z3TV1UFL6YIfZAmzDj1X0bijg
qtswrMCYsPPTDnOLwOjSloOe/VCBMKDRjZwuoivJj30oUxrDEFvTra/AHuMo7uvy+3Z8r+jXffuc
nYuXPAuQ+mNughJTCPzKO9SHBKXgPtn+0sYeLUGfHbdPn64sQtZrAeDS+tJr+HYdFzDyzutOv/TG
ImPFE0r6ZVCwnA6jmjmygVyn/bXnRXbEX7SDbm6qOvToOwkFgXLiXPHCyMMwkcMfZQIf+aGWA49h
0qQuciHN0vvB62n/v38qRZrC6RHGg2q3hCcg4s9VCbjIV0qYsXHnFLxo3hdQxVlAfsttOewNVnEU
oeHdEW6Dqd+aI1nIQCFY01Bs2yrcBbhOyQM9Ap/b6EGU2BXyHbjHSz3DgZLvLLQ6DhrtVKcBZHfy
akE7MXzo8xBN3iC/jPC9N7S7LMQFfy/sqUQkVbT33g1FQneWGyXRWEZrEFvn77OWdyqJvr83qEBn
dxsD7uOzcLrjBC09f2iDEkXwBNB5Wxymu011K5+cIbvH6qCFjrnEqN9WP8pr56mMBPgWmJJXJYat
ubcq+eNd+IkIpwbg4w2RUS2X34yxExvvSKQ9T8yoM96WI3KGDlVD/Upo0XxMnE7rKllxaiTS8SRP
Vh8fLe1JN/niPGlRQIPnZ2+DWbE81Ck/wuwpB4uD+272dBkDcDti09k0R1BnponIw6XOE6bNGgYh
DSe6xRZHvOvZVcA0ZCvcDObkkDmEhaL9llpuFBkfH00yCccu254excveJsSh6uJ7MDco8Oakr2Un
ImvFbyy1gX2qfnUf+eEY0b+8bRkKZcm0ll9n6wHRrcutljJBxuuEoIif+dJ+krrCjCQZgKOntRGO
KG+nLBVcxwLMHAMff7+KGxwjYTSnkDEGSmRswBJf0XL571WFo9Npw7aUUgfLL2GG+tXD/nR+55q9
H5Qiwk+rgX4Nee5lj1RXp1rz1twFiXA2V0pxy7iyGHZkl3l990LkwYTyeUQtuSZDD4w13OyVVMkm
Szp38ISdyMi+gXCI9UvHKWzy7dg1GcAi+ZbOfgezKztlq8aEAtar6faWM+7yZ1MK/RwI5CBx/MMf
uUz/ZWWkoslP33W7i5h4dIm0HiWD5OWCAIH0Up5n/QR+XSGh9SS9JGwcUhAfACn/FTis7uIavela
INhud7nWwQKOEhiKEf/aPRtKw5pfYhi4CScqIwDJp6xSo9ClZvRM9uSP9unQuVMXzH+DfXIgmsGr
mrhb/ncFvEQ/CSCUzzN97OG5m+UdnRR3RLOjR8oCpqC9HZqqoyFvyVq2DylTBG/8gK2i3Qs0R3Ub
Zie3AE5oTNr+kH8te1EQSDNqCFgnvzsDS4CJDgKQR9lMxPE8dkOuC8odkWTZWY9ewRbAkMqxvkQK
y2bQYPmfF2SVefz86skEWcBWthYIF4A4gjmEOIyvu16tN4I1TU2mfs/4PIF5k4ah69HVhZkR4WkB
R3FWXsdM8SUHfZf4ZmOaI6puR1KN+/5GYgkYh+GG/s0G4wCCA1wmiPw1J0yFpiji7c5v3PT/P9n7
v3clTrXJ06ZZ/+Kk8PBHAJ01ldgKxX0+5mFQt59kUHTOmU2vXIqUP09TAeI0Jpie3EKdNfIXeiKB
+ByErs2Izuy2zW/vXasDKj1ve0MOlFseNkmxdhbr19ezGzqJWK9NP+MtkFsvtrhfwulzMzbPrMcX
bU2QBeM1zgP2JORk11IJxtGqS5Y2So/kcKH4P5lzigxqSFyQ2ozM2P6bEPOcWWWlhjnZq+LQz5uV
zNF98i50T1tpGHaQcabCmD/wSe0KH9HKMYOcI4dCCuZw7/bKeaI0FhvdZZtr6EsWf8jqOUxoXcrA
vrzK8iahMOiFzXgw1jed4RNdRPtCIBD4VH1wKok8isBDh5+JEoRpAD9r8hdXQkC0RqxeXfSsack5
YWJF7Ju1FUBsm1cqzMXNPnP4R21zJFV8/il0OD8InoIquHUXjfAVyheReYlQsMKgmJUeSjm2IaTC
zMtqw2UJBglRC1uZCXCQsHMHI5oHs+g7oZo2d9gDNgXWqx+G7iqLIW2BdeuQ7OPl31OzEJyGDFSl
SvK+MzH1NnC/6vzQQcugoSNnpB2TReZXg+OddvQ4K9XMnxcYJdIeXOhIE3duDjCwkGRMyuPihRap
2ey9liSv6pZ9NujvIGK0yi0FBRcmKOsHJW2zwfFEsI2vqgOf/EKDYxBUV/dzwaJ2tS6m+AOiIUbc
SMi02fgQaqQSf9M8wabITSHYUy+X3Z9oGq//zZJr3BuFpTTSlmsM04oZuaCK4TiLcC/y31c8oK0k
kTibKlGm8OZvFkMwDWs6Uh1NRFrDTwgS0SAjqNXqR9ketL3y8+abe+v05FErzhleK1dlEv1bUOBh
BWyJ7ezz71YMRtgzeSC4axVD7MW4pz9Lu+xbHTD9pUAup/RgG7DNZSYI/68CplG+9uoG5F97JjTW
TbSlaEpON5hEjKC0dfE64hs3ABo2pJU77dJjTYb2mtP6xcix+SV9W7JEFgx/uHPgvURQyg6alwhv
jMGao0lAxfsM+EUkt6iHtaCDP4CJ3cunwt61+tDlR1l3XncSboktEV9aHOnBfSxn0ac9DX4Ph9sG
hXbrQMxlfH8JnZWHuH6HktMop5X/X2s05CFDPrx67abwy1Nxj4b6bx/VYVYdH7sUgSs/dmE4NVLL
8TQZSiGUe1EoTIB+2AH/3iU5144rz9XoTrFW6zmLeFG5MZfSPMd7G4txNP0lhvgvUJlNVbAJxZRy
6ZgEucv/5LmfC0UX7QuZoF4//v2uByMQVldiUvKFC+q8NxrWapFCD1RQjMKOsJFPDHBdR3UguVH9
NiXNj6H0/V5P1cQFdkXQlqZJYLZ/J27jTSZfEjCa3PrqV+b1AR4mX/H584qVo2bDUcFc77lHJQ1V
wG0QSL9kiMGdOluSLh0MoC5dxbBHRS9zK/cfgmPUHIrh0iZKCx5QRnbZTwkhYYy38/eAyC//zhHJ
gVnKtEp+hQZrH8ijyAhlsvrycseUEHB0xZsY9g+W/8kdMH97FFfn/SZIzt3QogYQJLSBPLIIuyDs
xPuRYclzd9getKSZSoKkZ5Suj+FYpIWPPeiUOxiX/ntm0V9THJLGPqJ9/wqXlilk/mxJ6SawTVYc
Ux2xRX5c89Zk+GYXjB71OZOJ9HWR0MaQyNz/Vfkyg0ViVM7N+DP2A8Sh8nksQMnKU04RVqEks3MO
RZjYfUzhOKCvCEHjMfKZSphX3rJHN6/15FUsBlnovCRdDfYS6s7iZJ+S7q3J5D5SbnWuxDNu3SMP
w4QTHbsZO2PEspodmjzCLcXumv+Q0s9Tv7s2jpIspyLKcweH3yQouWdIo1x4kyUEOM7El5wj9C2Q
qpo8EVTkeWDHnQ+y5tMKmlP0JneVOY/6AKrP0zQGXFJACqLKH/wxCzBNdYs0IQX/nIztYWeT5IX6
q4IKMWa9jnsMDeyPOTsC/0rzduj6jO/KzVs/nSsAZBxI7wz12tjhsYtl5p5UuRQkBdbsx5iXqf1e
o4IP9/fxbCwrtWWTEsHOY2aaLfP7ZnGkY4ImSWAdMQyO5bh6g0Kf4udyigCqdJdlHCLh1/5WkS+K
xvooKyT9/pcEjuWUfeaDE3e+bVGaxp+iup6c4v8sWYFvbt6chyldNviUkgnArB8aKo5FeNoVsECp
v3+j7yTq/X7nT7cFjutfVWAvZvNH+XgN8b3ES0GyZDYSzGhiEuTr2kX+0T+Xd5pcGKow1OshTeGl
cFjErEI7dH20Teu/yI0siGsyzYH+CED+VD6l55ygYIWDSmeaXOYxi5acfmdtuv1lsrhi4wW41jXK
mUuTWAoSeoWVJU+bLcMIjU7I77a1IkkHB0avrJ+i+qxdTp8iQ+A1cWouI68oPk+YwSfWpA/9fvkT
yXq+7ebS5P82Yb5f8B+wuZ3pjA/QpMbBN3ih5vtAejx9Jcx2og/RaAqSZDkwxjmGij61iLGOlmr5
oTz9GV0hNkoqIGsWdU7cwnBX64Mhjkyc9UGzR28w0FXSmRdE/0I7VYVEZOaYfTaIudiONv2SEUTo
C0oI7x1O8N6YdZdJEGOpRJjnSTAYO7McLEE4ODsyzyyBe9ijyLL0Ye4F4jWuAaMzcl+mN1WDqwVo
TatO8R/Us7Vor5mIaZ6rPNFUPXho/2QMBXBI9j9elnAfLI6C67ZV1p0CKQwRlawnM9whNbz2z6ym
onr0RyKI3e7+ZtbPC6LQVQ2wWYJPPDjFb/1qBI+A2GzBy5l4wmdtVDXXyZYKA9KLO/6+q9hU6IsM
Tg+so2XA/ZouKJ9PoHn/qSyjIaedUHrrxDm89LD6ShLprH45VY0/vTYzkCA7+0sYp5odcKW6sTLq
VRc0mMz2/q9DoqwmL1LRemMRmuQHIXduAVNlSXOPUGK0c4SaJ+iHS0ZmeHiwzEqeh3uc0y4gNB/Z
R0x9j+sY8f1Dz0WCoxgLPfOdm2KkETS+vaUcZ67vcY2QgN5Whu1/Dxm9U19vyDycbUqQAZ8d2CPJ
AA8LflYhnW8MahmBjxskHIQzO2Z9S1ll1z88caKdKuP694PEuo/8qQVuqXrDdd8/RXnc8J3wflyY
XnsBJ7yHs9uBOz2vZowCXx1PLALandVN3sk6/xoLzgCD6ZmnO0YM/KRIdpxR5r1BRqJfVmgNH0YF
5Mk5/NTWlqLK63ZaZhlIbwX2cBfSJ7l3hdI1wec93SDoNqUNDieIqQjoltFSeubI44UgjanWXyhA
UuXy+XBl/zkD4F3EHHOYfVath0SdpQcHbV6Hhj4O4gqjBo7EEVwk5Hdx3QAPZf+/d6tvcAQwGRFf
glkqCfv+NX5f+TRmc/ea8WojJtnvGTF0vmrcR8f9xG+V9aPAEKRyYTWqaJhq6iD8ytwbzCcWcT3H
DAcPVMKUeRvoT0iox7WXMDxrkqi5Tyiqal6vzTbr7nLlbBBJN9BWmHIylt7lr4mlm+bndnrtrQ+a
2/10Nf7rSnc+GdMomXBvOHSoEichP3VuIyyW3/hye0IofEDSCkOnrq3Uzbiu17Ua6Ncfp0wPmQ8s
sgSnXUGE3ztwII9pui7Xw57gr4yeLKN7OvElFfM35vPpCpRGZrRoBTVh6Eesw+4tZibgKNY1HAYs
VlD1CMEubCVq9ZTT39AzCihNSs09JXI3pD7ziqNgTUEH1hyINzwMOdOwXPY6JNpQTrm0stmPSAu1
KGcZvI5hlAKs2XdjnhhIpYpow6eI4bSqVEobQ8UYSYz2SZCFZxpcchx6ug2hK0yVBaxClWX2AYCC
c8r6wbT8fnI0tKQ6NphgzW+9hDmz31w7SiztXwC66elGXQl7mb1eYA0PHME9qLNl7cPptPFUBSuX
Y5Yu2TPyL2ZyL3bpSij8B9ClLX52sPuSVLif1NPcHYQFuJ0S5QaSPpNhIoeJWFl/rB87p5BKLxAm
OBPqs1FEqg2OoefECvVehvOb/x6Op7qwZnfqhvuTHwJKjh4UwKPUqw5s4ZJvoXc2NGBGrCZP+WK5
+S05AYUD7HIyQPBYlMyPj8jNVgKrUPdaA6eOuWL9Zl6erGTlcY78bfoiyay6Aa8Vdpf4tp6aNZ4k
+HseQmufwi+kPvkv+bsQfUXue7u+E41Voa/00/bQnLIu2z/9oBJSRozqA4eVpst54mNvyiQrE8WD
v6Hq/DV3yUnaRVypMLW8SUSTi5VrhV7FaxOCp5yB3G+qn+uW4QBY7J91WZMvQNm3REveeMRSmk5C
mqYHMmnbDBCFetYod57BW3UmNARukyGY2luzvo08pOJi/UfqwNp+9hb33WwDT1M75bk+YaMZ4KoD
iSS+uZD/41e67pKouIVy3L/+XI5M4ekPxVav7E1/epyRpDQRK0Z207WZbN1+nS9ZXtnXIxw3/2vQ
DyQcbjeEljzwvDqnVaRwHca8g179pY96KUCPhnKKs8TwLWLUYabwKQoZ3QQ0+yLOzaSLq628fE3Y
gFysKp30TWgaex+0ijwG0KlawFFv8/Zwn9klmpMOm4P/y0UKaOMnqb+9krIEAoXxZrM5cgoFM2Tc
pj7VIcYXQJ3xe10ZIENZclNwg/NYHV2fDGnxojPJ3cLeQd3McZjB9ZDsXYs2tcBnw4VMUjCEhsqf
1SfLgMaEU0jzZEP7MMMbHMvIiqdeEUarGUGq4Pu7NKAZmb7F6MsuReqHRITCEVx7MdBYMTx9vGB5
Hz4RlBHAPzyBC5lMv67AAXe0OQVwe4Atq5ElkadeEq86d4Y+0w6pTtqnWeH5/zBpg5EGIeVPvwxG
hBLgSsxdU2hgDMTTgzGSvuF1iTeCuwGmgmShLZm/psRQVmuHuz6ZRZP0VqnnsZtGvZkktg6L6i6M
BMkrW3R6Fvv59/4BJJ3jSdK1MoOXbKxi/UfQdiYuiGTsGFNFSRtLOCmBVyUIrPd0AAnxK6V06vnl
iDFS+g8V+FlcL6IbncG6WV//BiiKhu5Vr63Oz9x8Dc2/t7mPzmU12UE07G2MSv204dMGIFQ9/1KA
fCmegwmHF90pC6STiiAua6l+V3iofRpf0f0ycjVbfrPUce8caAaqUyXza/zheXuF8UkCQodkB25b
h/96uj2nVSi7wgvM3R0koCnbvbh/uxVrdqrLvJihGJNrMpjuNiFd08THnOu5bG345Dn35uSuZ57F
5drcBVOa3xVKj+ORNK8y/GQwDqV/76za4iNq2t5h/TNBTysKl8mXXvrCIoec8KZDH/ML2toGZBMw
ixTm+GW00sha3XhmqYZK8RhOBAQaNrvh4iRbqx2iEnmd6uCxldluPV8FZ3S/1QNTsAf03sato+Ka
6gP/UzJGGkLHwaW14S+vDl3gTSF1t673JvgCw5rAxoGprEMIRl47Tk+3zBKrm7OabAbWwUnHWNIl
zY6OO7MUc7YU7uONRuLo6RkmZWC/+mItwjf3b38ygdUcyQFwzezMDqHul1Ob+v6WN2z1mHy/JaMo
7VHuB/YeuWbxvQTEU5nURjOlVMKWMbP/YmvTdprr/6xH6px1QXPVjGi9VYMCA2tbZD03YugAxcMF
VMEyVPi3iPEgAtF085/H3IkFbWoarDot0u+Hn7DorHqg/srFiMkis8jAdvmdo4zZbeiRVR9Y+m5X
YvQu2rh7SzqowqPMoVMTvJjUUIThU3QSujpPHqhWpQAke6o8cn0WYiGPYSv4lAMMW3yPpLV4e07j
9kFvufnlakh3x14yvabSlkD38KPbJbGavo86tt2LDr83L4YwtxfzgWe0tNVnjvl5KjlLCOhSaoiP
FTSsqlzoqZj9ZYZ/SoBRajZ2VqwTETPuGAolFnE2dLbMxZtjRB0grsbYeCWhobqwOtt8zwgRidlA
UxEuAwCn34/HP3N0XVU76JdOUTLqSkGUzZsA856kdTgimKihah7jYVWmErTT77KpOCBe5g5oSxb9
Rf8sARGLIecD8AhD+YnKTt/goHeEzn0LMOJbYW90KtEV0KJG458/BDhFk4BtOwn2OzX8eAmuwzDy
Bf82mqSytX9OkIO3g9RBypxjgJdm1F1GN0qPMJK8tshKjwKfjcwePZVXoEjLjJFYBPDDWNLDasd7
hXV+bfdN1eYpHhWm4HBrQStHZkw81d+bzLH+O9yU84Bge5M6GiHuwvbnEoABw3bOPKMlm92ziVXa
KnxC7vWDbkc2vb0clKZLYXGaAYXgtJh65QQaudgQKmF42zU3VIcyMlmAyDvEWCo5HQNboSvUeMNT
RiEazYJUzorPtmIgfSPoK3mGA+2Ohf0DaphqKAQjPWbYdAUAGMEM43K4/I5YBHD9jHYw2uAaGNVY
jmQUetvDU72PjvivJQaqBZjWhlk9P05Yr0UJypYqxILuApD3oDfhgyh1/oIAEEIkFUcnNECISwOq
MAbiVOhCnt6U414qwgb79ZoEsutgZHMrGs1PURj7qIzT+iNU4Y2aledf8Q00M8/zswm9ouXl0lAA
OX6LmFxGsDX4mOhsNmDu2D3s4yOKe2ymzLs8OazZpB4kTz8lPPwDRwdn/0Y3wBf9ym1BFzHwJPTj
Tp9ZpNZ9CimNzdjS/GVwb8Pfl8E5cvXsyhGar4o49cpqSmP4zOgG5a6Tj+j98aruS1J4YLXUPyAD
GbiX3dchC9FjDobX5oIaJ5BWAq42Y63kpvV/dsvxDSG+rLTUTZJJxH5+Ao0uQEJ4wXe2ismDf+W/
ciNjg4MSxNiX09/fYnmQqCRZS+azq7Jk/gO8jCZ1LTur5dDEPhCbhIIYTTHU2vmaXJ0vLPStFJ3i
wgitarw2NaOfuBSeJuHduN9t0TJ4rPPD+gH47heI52vannFuUjTeq8hBZ44hSAQP3iNyzJoNG3/B
SR1wBWlZ2JVt5GYBzRVAITFtfBZ6EmwnUN4CbU0tTxycRVXCaTOjrX3O1/HPMloUmjyEyV9sreZc
SgBBZ1cDjYukLSJT04EsfrKbzDlqsDMwQ4skHGonQ/oIYhx8wZSBXy7wD40JYxjSmplLK5qdhcm7
fvuCh4a2xXpTefWLfW+BEEsxc1ipemBJ3tQ7YBj8bjWIfA7t6wFhfeibTSETk9N66S78V3oEvCes
Fo6Xo/YI5Y5QS4FsWefmu5VoGnyGM43khBLoASqRg0O3JHcIAhmvzr1nGYDc9m7LhPzVczPuyLta
tmvwAh01KX4mwUoVmGwQ71JI5VfwUW5HKmUSp97M3TfxPZ2z6LMP1rIL939kCKgMIpLAkJjMpF1u
YeW9lqeQcX4A1BfU8WfgsCCnca07fPLGoTPFdSxPKLbr+KtQjL7HBWrsbH7P+fJiK92pmM9VDvFW
JYpeTBGraG/CVAE44iI+EIYL3N9QyVLpJt75zhG045z6rRGagYBC0PXNZ/KNbZmd7KxG7JhX0JZu
luBTQtq3Dfk8y2UbMTsAXCPfq6T6OfMRELPFLfHnEREHWbnFid8TMr0kgMN0NNzWe9jQuyXWxcNX
JDT8vF956+lAFjSGvx6jyPRGm5287T5UqCTcLXkCBF8FbIBuQbeOsAmJYUyTLCVKG0bvkNGpHuut
YQwFhuV42AtD2x6+N1WDwLMjsq2/vvb24dL4M7wNQhPwRY50oTCf56JTm27+eP+49+sbq9RylHXM
zOdI930g2VLIHE2+j/OY8sIXdmQXfIOCIgGoqbbRJtsbYu4gzZHa9So3J38sfSAaU2rm1DjV6O+O
lILfK/64zgGUYxUodKdec4oTmX+gp805zfsghtAN6GUyee4amp1maPDylaADXkyA/9jumRb1HYrO
a2zgIv0/rXiWwaMEH9OauHlzPjFP9pmNzaWS3npwE4yeqvKz8J4kmu7zKdQQA/v31/fXoO3KAHs3
jYjRML4i+MSz+TLsm7aMj1I0Jp9mhVR4Ctxkd6SnRk1xsylk2tLto90UObaa3XefONCDYp+taqVI
ILRHqo3dcNNuZk3gtyMbOuLnGs3Fa15AtYU+DBga1RjzcBkqGu+mjuuc1j1ymPR2YhB0kN2Ak1DC
SeZwyU5z4UQQ78HAUhIzWkKyqWwWqv9aJ6/9RHVulENpkWsENwSjbk7zmN2/fitC3HzpnkAGJGSa
JrPNLreUOOoX4ZgFQp4mZnbQMGjEmHG6Ev8NBdlhT+tPQBhd5WQgi43GzYs/BWjeNe2dwgB5MHxw
EABrsBkwsK3BekVxuh2cV58dHEsZ6sxpZu5dzQsBcNsQcQCF93w/+m6kIUI1cJk59cHk6iAAiuKF
fd6hTX3vyOjejeih/ZaKcXXdTR6EOyY7YUHc2R5yTntW4XID545sZDsobXYYEIQRFHwVujq1RH5e
0sTYLJMkLZNk//x9qwA5eAHmgzwtj9Pn6oMONtJ/j0s/6MX6RU8uzWgS73f0lz1QZLcJWTOnM5ei
fSff7jH2x+4WlWWI21p/47G5kjKLcKvC4YtZvy+dNT12m9QrUsjAKumsCUzYsG6Tx/gmVuPjlNaI
NithzVfaZ6Dhv8PdHquiWYHxYYC5aLmgzOnb4eoB8o1HC85ruP7jhVoUP0GcY1TmxPWAI+g7ojAx
ckzEBPAL0xheggMgqDLVP5Oq/ot4ARqERY46PJpuKKVIvSsN3OYrRQ/aUvKA6zPyRaMz31hjjtYE
i/JNt/mOdxYbXoq5hY6SPoEOlpxZG4/boaQpRwFSZpzycFbwEAYcH9dzT7hVhf0pYkXIov+4cmIx
xPJs/3+aD31rk44CXVkj5qW3Glef833JBJs0n1k9u1vbMx4Co4gHFrBAV/4iJnmcPUO7NhJhsWl8
Lm0Si1XXNXiyHQLNTVe0RyYgsXrYfZKxCVJhd+tTqL0qIFRwTsNSznJCMxItnJEt7uDJxw6Cb8I9
0zvKZCs6drunUNWaxnMhQMkbbToEWNjgdYlSeIo2GuSOW1JNKX5BXDi2R+XqhY1Xw0gvBXvyNJGp
5NT8ESARgvzOnLDcTCPgl9qbz+WYiMPuJekGpsqCU5vzm1js9VLdvQxqXSrh50GYbBIbgHZD9nWP
F484KiQ6NsG3NpTR1x2f1kVQJLfcG+mWiCUtgBC3VkygkOxpPCozXfvVqAsDUwpm8flOJYGXP/lE
UBTljpgTUl5UXOuQtikm5Pt0cGEo4wlDucNHsw4U/gxcZYWFlt5OWn/EFBsoCvjmqyS+Sz8oVbK8
HnGPOpUqMIBFaeaqyIghiabYNFvdj5ENUXcezcssL1eFH39XSqu94B9cN/irjXPeSXhXhq/n6Lrd
+xcQ1LObW/si1uC+gYgH2BREebAHN5ED76XCG6vrQhkH+uTBbS8ydC+pO8wAaXT1tczGSpuX2x2i
Ga9jN6SSBXi55v14+/M/WZyKJnIkBMOm8eV0BSN9UVJOIFmgr7L0MaxHc6nirZ6pmwu0P4Y7W3oA
v1HJmiekZNxHL5nttEq08dVgAvvBVdX9fcf8NPXO7QfS3j9vFAyM5faDuGcJ7UZFKHgwCvkSrLBV
plI71+9FKSF7U9UAeJEc3Q4+8hjI7ziNGYgsle2y/ccF7iYQ+7NlUpVkDhbINv1Ign2xKak3J5Xe
GRcvzhGbxyCtRo7z/Z3SO3O+FZiPB6Vtrf+UO/nNm05Pw7ExvDsAjBVGO8Uzc1v5pkDNOCX7gcwR
PAc0VCW6N2pDF0C0a/T3Du2S7eGoGpoFdELeN0DQ14VMqiowqYkh+BMYsBmri5SHrjbVac0ZpLsp
l+697HRScAcluTRzpY2W9WaJfuNj7PVBAdQJqx1MRfrSF/ciKodmlsMtbBOaqjs8rGs7JFhX1dRW
tCJ24G9zqbcaiET1/xQn15supbyd/FykgLD2A5VjMhJjvv/S/GCsUX/S2pZago2hoqxtEYChV5F8
NcZrSp052ndm0rJT1CGLSoYCH9zdltiJ1kS9wFXKjhyAfPnt6xcGFXiv0IydN1Jwcc3WEqkmRs6I
gSp2dSw35URugSk5WEtlfFGGREJO4Zyam6VaMxiy9w089qwqavhi+UWf0r467LWxJ7uH2y0A/SNG
FywXbDhP7P4YkWMSpPIj2Oynmv/ONp425w7cO6+/nzFnQRlMcQcQWUpF/8Ck8LzOWSnCrNI9oTgO
PqNC1c6DKLs1d8LGbA/+PxBCZlXRhexzksTu5jhBUooJzd3xCQYu4RLATx+sSv7ixzVDXNnQb07j
6cTunndvngDI6P6yHERZFJvTdp9/OR984YQ31rn7lqNKXMvqaGZTmtPytGY4O4sxUtEiGSITZn+F
CDV7qbfZUJPEWpX7Mr7DoeNvgqHTY5blSY1F2xe4s2FHxKBZCgX1UEHoX4RxCo2KHng42EG2+rpc
3BP7+mRw/G3NcSof9zSFCNi/IiK9Dvbf55e8gLHZRfR0Us4jRpbv3a5QngeBK5dZnnHPMNK99KQq
0/EnAyIAmhkKdXAJp8Ky1SrRijV+2r/8kzpwnI7v4yLRanNDXbayDObmVHDjpQoA5XoEYBjfZlXK
FYSZ6uTsvpFV6s1FvRq95FvZl2cv4pSleNm4RsBXajZnyG0BOsIiqb8Iay3bx6VPFP/1DPVf0POt
ludCnHTPM1IfkKYMbZzJqOhrc8XcHa39fOG8d7wHJeKTgYRAD06Qo5DN/I1ztSChHo2sxoCbLdN9
T4rI33YzDmn8xtWa+daPy9n9ko/JdDgxQGnku35D4JfWi1dWwwCYITx74vyXx2EwAiRBHXhnQyT2
XMhU6gVDxOcgq25WFc7n64VwB/L0oOz1/EM/eojTkT//r47DZ3SCRxb5NpqCSl0dZ0kp5zG/0T+0
Nd1OmXHaZ9Yg+69sW2hyAP8oScsoysfMkof/hf7sk0gmgTGIXWqtyMWJbubBUbH3N1OPvZdvHEqV
Q2NcQZ8+9QjuvWVc9S5L6QHzGWF2mRtrM/LbQvzAe/ANdt9Pj7Y6v81QZ1wanC9xCset3CSFZ1Jq
4f/PxuLCKynlW1hfXnLaVifEPD2hfAwxRQqvn9NMTJVyDDTXMGGGaY3tbIGKHVxbABmcyaWUW8cI
htd20fg7B6A8S+P4hROmFMW+O5WhdKNPEEK0/CRBdTSMoY80yWM0AJSSc7zl+T4AG9x9fk/E4yAK
XGLt02YSnYXY9vxOAovEipkUpjyhL1fO6NlX+1nYRxYaAYd3n6x3JanQnXapPMB7m5jNRp3MyL2p
OBK9s40ov+HAlqCsNXTBn3z3qp4HaGhNW0O6ptz7q0LOTxMyslbW00j+5VDzgcpHz4/9U3t+IVWi
TEnyoqHLEau993Ho2RCeVpVySf6w9F3SGeSleETwSKiZghz6jdXYFhPe56V9jmimg6jasA+wmWA/
N0tdGNzKosGunbS111EVSxZHyflvyNGLmPhjd3ctlIpT6BZBHp/jD21f6uT8+Yo91gFKUKZH0B3p
EOFxXzq91DG5ixV3LrjL0YuWQPwBlrNvriA5e+enkSXfFbnfg5BJ8y+RNzv1D1stpVey00nmGfov
XgMzue3ioOYO7t/CGsW8JvMSlpxk5s4AjxNG9fOF/bVSq1/3v4+2zN9r34DCph3ISqXGMZpuP+xV
NtK/Qsju7UmdDCUz4K4OBPAPoWf8fPpnNicf9rVK8bxbANyzWLLZ9pdjsCfBzaBc09wT7Gjx1yoK
nzs4/AIpfVnxd0nXhoshuejcgsY/Zdv5GflOIZrD++dIgft464N1/SKTP1TnmNZIMdsu+QBiYEDy
PejpYsuW5o+5DsSdQ5jZ2/OD7NLz3t2nG3lm2FQ4Q9h+2VmL0LNT9+/zUXJ0PC1ZcgdM6s2KsIIX
mm8lTRLq5BPgRuyjCM+MefJi0tVppwyk6PQKdXMOd5EzhNAopXpfIeU0woeWd+kACA3d+pqv5WyW
C1tZOjp/76AKxOjMMLURbkRaR/yCZEVYyWe7slKPZwq6u8GkFaClTOf2PbJqYq7SWl5NW0QLr2FO
M20hKyE2x60NC0rxgprhFWKI+NztlRgSkkuMvg1MoRw1ytfW78+bAjFiMWEu5+B+i2zXJcztqWja
bNQfCn8zqliO4bceAQJY0FCjxxslBITQbakoJshCQLkITU4pDJvfDKHpgmY1Vzz+u/2l/UlrVkkE
wgCLxfNZSa8UhUHnIRSYiXgjbnT8QVEP6ArMOjQD+/CTO4vJGUEzqdmHc1078i/fVUfd6OeHWfh7
ZBJm9sjvGRdWE2XmE3F0zQ2vkjnHhpxxGHv4aANE4RGC9JiklJ4FnupyISIsO0syHj/kIhzFLC8x
cCiTa3MQZhlq7Hbs5ZTIiRdEcgumFgtGJdBk3cPjzFwzhh2gYxc04yC/qpxwm1ry46YlpxteDEqY
0PJRQhrNJaQEnfNv4tEIBFgAaAmZGHq7luawi7G0pqfJbroovL81beysnhLZ9fSlHz5BiujH9p2A
aOL8VlhORZkKEYCeb2lUsc3LBJLUHvaVKw5RTWd/Z+NiLK/jipCLlbyYq2PBKXlg60ijzGHwEgFV
xIfd4Ad7wc/h0gICNKmSea8FQnunM4Y9MCT41FGXRbqy2M28fAjNsv0G8/VKAUovODTDo6JXS+e2
XjALk75mzFAUDA4juX+Gte1yt9KZZt5e2QcP+95KNS80luK1sftQoWleZ1WdLs3Ygu0t2+J3/jnX
4rD32uhoz+4JRrfHFvRFR7RgO9dYLTIptiT+2bYCwQsMRbUR9ECUlu2CtOIWEOYBeBD9zx1iR4f4
LqnMB8qsLi72W4CLnVRwJh54dcYODFjJ0zl0Sj2kOc1h8bY6KZbp3J/ylTpRUPRR+j+D/DzNNYPz
aVUKD/REg7mGGmA2jltEhA6s9uq5QpliiAsC13nuSzUS3lEXM3KKTqiAzQbHuvMfBbjZeVbZS50R
4G+/RmNaz5rRX7ddMZmhhQFXvdBAEm9aTZdHDuAnlh4bYVBYLu9qavyW5CPgVbwDPXMEw2qFUlz1
ROnDZRe1giQ4r4YvoRooyWfcN5F2e7gpkI4ZyCVHNIrFP4cw56ZTx6Ix6a8i1nlwo6ZNleH2aqRK
5nkm5ny9EGf7/EsyO5qG6OD3euobmJSQur7/vuPlvjAxB3ChRP5iQcNXyg3t4kfO1cj/UpBGQ/MW
SnsEImpW7dskRQ0KMxJRB8AEjNlRSPcVN5CrF8WfTZGxH0OMGHTmG9B95R1DZuMQ+j1t7iVzIYlD
0IP+Nzo0ZlQJ7zRx2M4+xNKVBn5NDBV86VYek32gM+c6TvURIhvqVvXDKr2sJsGecyzXyYVsNKtY
Un6oyLl3iHjGlm3iqBOCw+V7eIit7kdCTz5YBtS74/2SwsKSJDdwfHQ0Evj8n55OMmH0BNKvSIPh
KWM+Qmc8jSI5qrN97jGuI0euoj7Q8VqBQkJ7bemZSjrtwMojyhVyf+nlQCMROZhoOwQimQrIrXPZ
bYs9Gh27rChqV8HaIivN5D/BwkC8C/FHxC/cmEAWjP7ho+0sNT+05LwJUECdwZQsXAwan7NPK19f
JGzSXMLeNAe8u/37GOl1dAZAkjZExOTkLSob77pe+cQpQtHxNwZckyk2MgYbkg0jSHGp4ZBy728b
XQT/XzHv8PlNd/CWPzh2gapHAN8LeIV0ok93vjcwCTbuEq2/NH+uDtsIIfT5j6POZLjbVQkzxn6k
RR7CaapTBBxONry4yCeyOGYNe/2W0pKaDthN8USQuynJzFrxQVFAUUf0MY7FhlvOKup6HeSU1YZZ
uf/+ROXYtraJPuNvNeDpWoOXuasJuO+ISojreIUM4Sf22OvXlzoZDCR8euXPyI9Lx0om3jDf4nfl
JKuvX2vl5EEt/7OBrA3qqhQffwgXiobodfxceZZ2v0dWoNb3mxAeVXJpvHpUpocgrbKFHRA1cK3J
X0paZPTlKZYaSHmxwJnGNKbLnIN1/9TdboQtMgoMug3QNRkoImw7R6siwq8Kbla4owNKzSVKihml
3B0FZjw6ObVlqtQINVj+ShrbXZp8GZ2xP8kLUoP+5w8O0IGXrSn1sjrHPoqvYZy/ori4AOS3knsg
tmPTM8H3hPvzBb8j97SNEEX7G1LSqF2AFWAlkT+J1pYdD/e2tNpL7Y3ue/HwBPwhOcHDbwwopxRo
HAZ0qJXupFd/XZTjCfFKEn37ydFzEoHitr0la4xSOmMAu/EbK+yrdwtyLTMZulWO624XoHBDa+46
n56vG5zlis2/m33FCqvvwlQCEmrrpduHfsVQKLYuU4QUb5Dca2Mf2wdeLL8yAv2RG6IEIYVtWaow
+0LWpJy7uik3g5TryTwYKkZ8PXZi1PmsWbVY1enJvGpFdb8Z1F0H4q/PX+MEnNyi/fgDNm7vf8gy
hgYTAEAlOkLRMBf0Q2jS2R8rhdGHQFFtllilfOpsVMNliAVNBn5XPyN7+A/GGXpR7zHr7ChkLFlC
wEyhadyt1sI9SHpT7KsYQ+/YQn9plrBMZkrSoruFV4k1YTF051a8ZiUdF0YscG+khQPjOT2TT0Xg
KdqOSietoGJvcAE21eJf4/CgCk0tCJpDGsL993/qQsmzgWENXW3kLMJjeHpNEUAErC9Ut13ZcCtv
eNec49YK6hEpw/ozNxsVdQmuUBUgsBp1DtBaTQ3fd3Sl7iz4a8Py7FVU5PLQO6G9DUOdUoyzbgbE
tWhhajicql6IQV3h+CJ8a9lQ2O+SKK7+LN5XUM2azi4rxAucO1Qxr6mGbeu87oIwu+2ks1pBbVuG
0wpwj9Q8YUXow+oI69rtOVjeEuBO2NtEsJSlnmOYTBs2gViikXAnjI+jCbQQyqGDZuuPN+6bqJDk
kKZUWtmTV7WPeSOPbhdL76TaZ1+WxcScf+Jamrf+R0t+wW4iL2+ktd/NYbGYZgxURWK7UVQNH6Wk
ijQ4kf0muyLWZYsSsyFUu54N8MDWD5+QWKuJ9q4ejvfSnqdr8VPpXazhcmwJzQaM6skhhz8gcccp
ajNOFpWr5Uvsx5WOEk2+QujhwQCqQgDElo5AL4boZ9pQDA9i8TS5TK0iaTzKtsSrRi74T2kjZW6G
JSHZPYaM6sMo+n9AFowgaLyrFOUyQHrhj17+4/4x/ZcvYZbD0jhZu8Rxg0bxyAoJLDq7zw0eNt0G
a2W3346b24149S8AzKtJH/6vvmP/Dvbg9IuwU7M8KhjhmVCbOjW0+1p1mMiSWnnMm32tam9lglDB
Co8oa4KmeiP33MTf/QYlAgNhInE4v9kjTP7U54c3AZQIBBrMx/+NYXTa+7BuuXNcUPq6eW15nowZ
/0t/1mpzVzZnUkju4PnhrYo7j5/88aucNKnRR9p77aDAoQk6XpDBwl6pBKx0yaahuzAGYQ2Khcyh
Vnp7um+7YJV+iS9X29rQ+hia8PdbTwAfM/4+Hx6ZjyFDJZbqsEknV7NSL9G7nQoeXQC7ByYR1hJ/
5Qwq85QWnmRLFa8Wll0WVkFbI5VsyWV5dBbETn/VUvvntRnwfPuBsuifHSKjCsU4D0M7r8vNWjYQ
oC0gPKsQD5QUGwmtwzS9ai1RpcKZnlv59+l+PIrLtzuteHbz1HE5v6U+8/yBJhE8YmQHwj/Rr0Km
RDu39HAoxTyT/FtECuNkITSK5MbD+X/f1zzFFUu6C37ztNJR6wYSGGjyz2j4G/hOgxoMGE9GgjSn
RbH9iI+BryS+WoO9XeTsmM/XJsg6dGcQvbxiZqArnspduQ87SuusciRl3f7GJuFfedaQg2K3uxH1
1hD7GkG0jrW4OS61RYnWbKXSshMJAe2lveLXgZCqozga6MpkKvo17OkRg7jlZYl5fPnZmVwV2OM+
jySui69w13LsgB+XchDQGKZiXseZVFAVX4P1bAH0h3VEZDY4wCAhNt/IYHRaS008qTmwucTC2d6k
R33PZ5YKSn20cRlBTCUfs8u4Tnn9RNa5b3NJHCrHbm7r01JsaVXbv1KbeSI3EZeIBRBDB5y6v+Ux
0sZY85wcCJIKB5xOKGS5hkEFJkg2ydw9yKgjleGolGvuEJurfFTK4BAbvcNhPRNQYFpj4cIEEiDj
AFLk583AOwZwtA3nPkBgU2tMbYN2zWfpmBEXAyS8/1sGJZG7i8StORqk+NMSZAoUvTUwovex3vNs
R8Zvg4cnuqrAJv3/KNosX1lPWC7VMldsAtLs2RGjTVwBYbdGrLPPQhrGjvXdFYQkXFe62YzsWfl2
aXYDX4BnM2cL/Vq6cfWRxRwg4TuaL9hoXauBLaR7MROfdDcLf+vCB92qrc8IfEVX0XPEzoX2RqHB
Eh55rZAvi8PkPH4ImHjaAVu+KoD9YU1dKjSGGyaWmgxIIRdrn+i685Y4EMa2AV72uTTxFaCDNZFc
dkSix3Vw/iVXLzg6POvvvHtipsPTFLb7anOp/xYkmB4H9uUP9XzwLNupsm2vLVf/joJ3W3Du6hsm
vEUnweE03FMPqyY7F/dpMslNWMOP5459dhfhb9xuv2UQLPPqvr6KJmT9vjIHnQ+Jv+egfYt7M0aB
SDsdmU/B+u9DrMW8L7dGpL7tpDbWdhKH06mtRREOJYP31ZsjJRFO1vN+MTOfWVYc2Dkd/hMnhgXD
lp/CxGrMsb1+LfR0ffJesTzKkv8zmEuLCwE35NihcneAA1uYgZKjvY2aD+ZQWxK5B5GPnj0T2Upg
Qhd2U21dPxs+rwEWjTvGnd39FM/R7nq7xAbKD6tvjS8KwjF1rMD/qyaudQwmv7l1h4WoDfSXZeHE
R2Y0RO93XUV52MucJFzyyE+6N5x4Fj5m1y+vw+ehEluGvo3JKCtHYN1Z0hhXFStvuWszHP8h4h8j
seOYzibrrFfTIL8oHOmiyjHtXNH3W6+gLXiMvfJ/3HJTxea4mssRdr1FWOBtKOWVvc9h6SvuPtgG
lWkhaiexdY79jo/3Qk7dSGVEqgV8Qn0/1eSoqO87I5JRiARU1RJn0CpwYaKeOrqk0DjBrRQQ9NqU
zMia43Fn+sFOH+rRifsePGcptjkLhrqW6v0l+gZebW6QKMmyik7Xl2LRRRS20Uxqd84/oSWTxBxn
eHwicmibleUg2bn2a7nzWmynOu8uGRAtqRnbICk+ZLiF1eXo/o+RQC26tpYaP6Pz5DruxBC0Qzaw
Lb4grMCwEsNSG69GMkPKCMOiGo6L2PX0YdG7JtNyFDkGN3JGoSLLXFtV7m+SGzih0KQcCatDHPtM
7ggWMxP4b4NIk2LzTB/hh4U8ItHms0t6sJY0S1NWtJkAP7b4DuPhipRaYQQeqwWiRu2SFW7+HTIn
02CJzkNIOocbhw2GVMwjrC0fyyK0dk4nY20g4RJLfmRyphjU/R2ooNCNHdtSOcI21aQzYItM+cWj
qjShCHlp4NnY3UnRkD1K+57e3jE8rMDep+sQfTrtfPKVq4IL/zBsl1Z1VJ6WVTsD3MZDCf0V0pvZ
8Vsyr7vaeUtouWVJuVm1eu89dPCsG4MdMziYl0GqBLPIuPGGH1dvW1V95J0/VJDZV4/TRx0CYJdh
7+t1Y8d6/yJ7mvAuLWo25eJEX4D2IDl1/MeVUzF59NIGiwuyJmIC/RubZ21KizU1vHWzk4ZuoaHq
qWcqQJxNO7WoqSfJnh6TjetEzKgvS5AxrQImJV6/qmPG7RTSZXpcsaTl7fqdo3edbrgOGYMChFLh
1V5hGrdUseFXLpzhC2fB+EI2/1T21dK6VL1QbiV063A0FJFKU19MID4CGSzgnXODn23yZXGvBegV
vVSvhhK9Wm/jR9LrglCwIF35Ype5HvvhoIMHOVQucYGJJyEduLj5gSKo8XO01u7UDFXWomArCtSd
7TYKQ8BnTWpf0xn1jZRCb2lSCKOz9x57lZaGaJWeoMfYt+Ln1PZ31NkledGqJFpl6+YO3CX8FoIk
XKraWeFK4BAJpMgkmd24+dwWxTN2KCQzdSVe0GOzDgaaXv2zYxjU5l1RfjyPsDTzt0wLlv3zKwd0
qoQn1P1r3dpu1uEsfKCsKawKlIT8w47tUV6+J7AnfMFbVrqdKPxc2MY4IoKyzzOaTjSc27BpzSmB
ZERcbpNCN5Hjw+pG5wBMcSnUs1OdGzt7NbQL4lVG0AUuSAq6MLU5cYWvW5L5oz9MTXTSPsOKcdlc
DPW5O0vk6L2/q4PPT3wI8uwB+XGUpi8g9To3FnyH/lsKEJGFGo4d2GsTTneMC/j9xpZjttz5Bvvg
JWKbE4QDICtZj3WBdhKLKb9xQkFfhr2bhiPRRmalXc95J0FrPt5GMIQ60nRJerZCWbWe0qlmebFP
mJp6BjU7lDvggA5Pe8VI7aooYugMFUS6XRBhtTpV13aTolxyXs433IiB/HBho1t0IXy4S/rSM40V
f/Re+Kt3oL9WVWxocUwk0mAMfnnPT+Lskkm4dDhrzRHi4P+KfysrzGsrKIZctZPnRP7ivgQzUaY4
R/xce3+KX6VsGaW1IganSsOs4pcDk171n5Tu/4GePJadqw4db2mNIcSkw/0F1S8IMwOncOmHgogJ
UozZIzLin7BUfgCdobQZShSelpQPXbApNlPmSNMCP8gb+4Vgpl1weUpd+cPqle8jcd1SytwCAQec
IdP0mafzGD+9gmUyid6CEQ65H6CJK9I5Hfy8dIgYd5mDUPm4M0VlmoO8T42xmOJDLv18sSIY18R4
oS7LX09FD/Jr+qwnwjyZI0gkb95cwrdRRKL9i/8DQnPHoR4wvBXBaunYnbPmxleQQKC4BDxtKBKk
pOaklcGha7n4LNVCLzE5lyjdXHjE+X8BP4H+LrVc10exnTWH1VqmiwpKPI4RihxhSkxiz8MM9VC3
cvITr+03L8Ds/4Tf/S+MQMkU2Ph9/j+oblLHcXIKJ2dTzqFWFYkBeKdjHIotLWIhP9xSvhoIvXai
8wGi3W+9uk4mr04tKZ6ERu0mdUsp6Y0LH7hOfdj7FMEMIu3VXedekNjj9unO9Wmirhawa6+SbsGM
NpgB3zZPgfUlnpT5Ndh2IrHdZoabCU7AUZRSWDtkmHPv5sd/ny9QGxl8PWZ+PmdwrVE73brXodve
UFFBWzhh6FmbZBP4KvgJadI3lal4iQUeEDiQsPIBAXoGYP97iIq1Vaq9QknwUUsoLLqAi8ba+zh8
hT6XWKokaZ714+R6RPj+6gifJDkkbGapootwyVIDww2fOiw6BWTD+mPJL9o7upFBBSBSzP8SD7N1
1EUD1OYj56Gl7dIrxwz7ekI3Vfk2e51Brk5niLOijDO1xhmatvW7QkG4hCq2UTtScxvTTvojZ8nF
0G/6yZWdWd2vvK+EkQC1h/aoAyj1jzS0rkA/8xWYwdDrFAMvw2m+35FKZwROIfXHuUrmEB0HCI1A
L8CMrgN88/pafOdxwCtn1kX5lRI3UytI/EDNWHg7UeObgCQCdXsaXB6bbyanfZr3LtE78vq8/3Qb
3IhKJZjzMKoFkGo5HRA01JfQ5ftQ1zRQLh0+W6P4vnbDRA9E8qF6bk/nGbPc1diAUN8s+XF5fTy6
YhIQNwuCio5hyVaBhZbwhyQVaiwAA8t/DQWwa4t1HisKR3yJQkc1VLI367aRsiHdIrFnkNaSW4i2
LKj36242jpyJ4U+i9lPGk18zpmXr5XBzB7hZfGBKuPYbH5rbO0IJhi7zZVIqa4DzrhQj6suQ79UR
mt9rsB04Z2f7x1QSDCUPpTR56a5EPeSfsLSWAWN7TClB53s0xdxl/2tojrHDVJsfPqAFDDNQc0oa
BRvSfY1W4Pdal7W2YIHLwX1jI+KXzPP9gIXBDofD4SxN54zGZ/WurnMO4muNjxHvsCYrsFqjV3Zh
60Y48oAB22mFo9ffNGHYB2O9CZhgf2buGhzDi+h+KQWrnkrPtGtfdA37V8OQqY8vZmOR4vROIuH4
V8VlfqWH+0k8Vr/a83Ccx+HaQ7cikZNUlxw3lxFjE+JIPW8wyhxg5g/Py5vXOu3nli2kqSsJtLZV
WwwZfotQKlbOrkDcpH5FOJDK+rtDe/8yvJccYbUtxPu4zwN6ZVuRpyxD6RDN6ZKbkJ3GBvW67/xE
L3Q+MXNaPcnt/BWfJ6Hcg9uVdgIEIYjbEsz6patiy9W18dJaANAdhLduwM5Labmv960XZq5PFqjF
bfKAruhnlBscJ2W1so41EaxtZ+Q8UAIVD4Ee4rEa6kccsmIgxqxhrB0RFpzuMXjPX9aluqH+w05i
esu7SnqRCqMbFUpg2Of/YeY8tudS38S9yfa7jkD4rG/okTf8OW3W/XqvwFzrVvOC80rJCvHeT/mx
i03q9oU1b7w9/fOHL9trgBCfew0IO1XVO13Otu3Gj3STF5rvnDsdTICVAfZ1Q0xJqZF++yOpnAKS
hfhpL/ingNLG/O4iVnu6eL7Hu6bvuBt8H4Auj3UuujwBX7gp8OunwDGFw2/4k1a/HhMah0+7NTPd
NTiuRg8qWP8xUhHOChl4aUx6uP9Kvaf6qnVm4fsFx/Y50TgYcZ+O1tecxKS35Jn0c4zOkOTMbzs+
i4RVM1dVqeTP4Kzz3WhWlSX5MhrtPnU6dmh94bG75Mw7IM52p5MCS402+HW8CtiS/yZ7JXvZJowg
zqWsjIf4+1TgehslOsnipTLmeCSqMPqqqVqUUyd1KHe6uqqAV7noWUO531glm5rIvk6a8k2W7FZ+
KMDxQ1UCV7k4UAecM6RM2TqbHZXaEYKcIWeyURjb6QXKvweWe+ztMiNEuPiYx9p0In1pOf4uXWja
ja2pPgmSnaHl32RphRQ1PwRKlYfNN1iuqiEj9acnW3IBpWCpB5khr8flVNKxuYIX6HO47WYWHI0i
/75EZDZpG7FEDXPcYebfySPFzpwLWjgSVCHCM5YIHUdW+GJ4UioK5FwbbK/qBvhEqpBrscqq+8V2
zQCDDhhhJ/jeBhDuPwFzm7knH56JC8iuG/iLwit5kcjrf90uPJyCZ/UApVtgUkB0PqJjubcT5bAQ
GWWJZ5TsNXHeoCiDIca21JmIJ+d8ROUGxgLvbDzyafT37sDbgpMG2g9aPIznldPFwDqK0hntI2O6
FPH67UjLTC5u2vBSnTWKffByLZaTLAi0NJaSA8vV8LGrQOd0MwxNlALBNFCZiQkIBXErDNJ0MuRB
KFePA+EiumdFt7+r0wTPUDq/3acW6sNKVT8Ms3caJxW0/8annPUn+cnquyQqQFhrpe7Cq7heVR+R
LdsxiAw7ziIOv1CBXAJSHx8iUvDmfukcah6lrkTUa+g07JAH/PArJBj3vICImfKIUmthAo0r+N/a
2lG3gFqVinmRPLodr58zfII/aA78yCqCqhqEwBzeHSiaKkM42RAo9eZ6ZI0LZOkekwOYBj97nQai
807fbm5EWkeBxr4F7eacd/hcoW0EXAyvP/NQYeNFRXOqa4EqwuDaOBaBk4E+YkM4v0y1x1GLXXoB
G9h2yVDDV2+QIs/1rURYHJ/17VBUTf51bC1RcMlLhQtFMuowKf7ceTbDkbpk2jfwv4+3NWsQSExY
gpfRpuAc72lwODa40JCQAogMTBZJTkN8+ItbKrvv6FOiDYWL/PybYsdpLE8AkCBBFweeu5CgugkE
1RyjEWcPRSUp0C6pw+rhAinhmH4VSQK48V16HFZBJj0sXcHD2K9jgX97A1vyuBbaDSDVf/of3ko7
UfyVaS5LDS/siJOclLWPup9P5OMovQ4Tt2gLigkhmAqzoUqtuS8OzpF6QkkKs2UBgKPEI0c/Z0Zw
UygcuCF2oX8zVxhPdispOg5H0B86MkBSESyx1mPuI771/A8p1hFhfuJlGD5bh2s9qli39XxEi6+w
wIVyZ4CtmrifqZgbIp672ScCDRWsujGP0nK3C61MPMKcbDx4nq3IuUWEUXcS0DWq/hAyL3v7Nx52
srJCHk4Gl1WF9fg0L9FdJGjeYahuOsGRti6cAHGeEygzNvlDFmtHk8yOaKvGpT2mehjmYQV4x9kV
Pa3piiXLLVBtzY2izJ5h7UiAaga4+B+9MNXEfKEmcMXVVeXxSMH69b2wsb4q0XjuUSBMsUvO+r2Z
bvbvcKrElToPkCTYLhD1dfio5iBm7yY39MjJ3KAXEF3u4AhJs2lJddxyJP9kmPUcyctrhV12d5hH
vRnPuv81AvsvEbhQakc7/G6VraxD2HksUHToWDtqs6V+RM70AyFaQLoBKtChetja0B3g20DHUUOe
0B3LaL8CRZ13hiFhc90y7Tyf41cVjJ9yUaaWV76WpMVidWUnT2FNttuwbRHiPfg9e8dnq0lNheJW
Gm1JCPjKuieULbFtKnTRcYYPM0e2rUHAsYp/4dF5wJGc9ckweQPCszMVFujk3e2Jc/C5jQTmHp/L
fNl1+uNZvPNyCB7YI7LxZHqV0U/F/t3dVqAW3OfLpqXXF2Ilz+1dm8Do4IhptnchTC2ykYkPmnP4
hdZmPVTcKbtBEbYKU0JYPCtU9dTVQEHI0guy4EqQVAb2BeTsJwtrsGWrqGJRl3wiJ/Hk6ghgsOVf
238rhFlqXFt7JxUGnJe2zIKtD9qJ37v2eaVfDwEvwSXUQ2ttea7cpibwWV5Lw1X4RscSvEtxpn1l
OLsR8eLO1dhw929CzSbLKPDTmY9HjEKVxddT+MFM1NqaGpAeNhZabuniN3l6n6dmhlNuxahegVnM
vN0T0x57D9VWc8BrSzSJT78rjb40arEYkvuEOyEeAeg4rW89vEKqltpM9aYpx55vDgAhKkyV2HPr
OEtZ7ydf8jAWZENF1PjBGgKEVj9xPIhCtPtKEz2qK0R7JdsbT2eWpSJTSunRD8LwdNsBFuaXSaSx
9JEFqshpv9/9J62XjSwenAL/8H7jszLKTaB1hUwpnebbqyjDzV3xNLPLL1bBu3j2IKU9vUpGXVo+
e/Z67KshOusLSyEjXc4KOaV0U8xIaP4+Zu9C71hPRiMys2voTRi15pzVuxJN+oiNP/4gPNBsFhfa
6oelvNB8SzEdVvQB+/2wtfYLirogSGI49XwQSypI4GIQYoO/HPB2UdGaiIfNhtFfQ/jYRTse8Vb2
F4Yvvnd2UCwf6VPsmM2DK9wlBoJWUFzVYiKYrXfv+d/MRdIiAtKaUrCImfhazOd7UHG+AQhJb1cp
9yvkm9Bs+cvDcH3UalvOoJL0gtcZkKkVzaq7JAJBuAy/3iHxbFfV48RHFYV7wyOzVfSWreFV4cu9
nAlHkejhK+bqaO/3DoRADLervfwwG1wZxgpaf3/ip+rdDgNLhHObLLXRZJBu9lde6Y87q6dhvo9z
dVe4MBONJKglOEZty/e1eNiGKG42GAI319ELlpRfu3ZdZEkN6eBQgdDh9TQ7UrJlJV2UvmGGg6Id
iNQWxWrmkggj007UwDYqFb54m1BLee4TPZNuRkihdcd2HwYBNb+rcdwMuvemgh1LFdy2ogFsWqpH
6ibv+pBIo9VQILEMBUJcOlta7OeWL+nQhiXMvhHeOZKFXSl8GC5g8lNO7MxTgZ1apUeAke46PWQj
FPfDbqGkW2JRaUQTB9vNIg/qz/awxxF/5WiPVKknPA7pA66zIz3jc/bkPtGR8am0gKjtaw7X/8uz
eA3J+3eA6BS2ybvuWUZHoN8ONomatZqgfpSPbihiQOFFvvg3e5VOB5OcdFiHNVT40tLchQe2eftA
P9vp1uCMrTQG8IQ4vCaS68J3vUPcxmIeuwtB3jMNlNWr+hPOVBXJlt0Z2W9tnqDFyQsa+fhEySX5
F9xYisO+nzYkJZTzgT2ODAd31HeoAo+2yNnjS4GYVNH3VAoGpxz3MY/0aFtsRpThRwUsHSw1I/2H
uNGfr9u1xnwLpKtRWE+cssT/3Me0Irjcjck7eYD+q69yIXqKSOL1yZ7b6+0otdmsO9blpT7EQG86
2buq/lCBcg+16GI6SrMc/G0NcVzUJHuJr/09w+tUvyjpMOlcTovbaqDIfzTY/a5sBvRWiyRmEx2l
XXKiODIpuQSMZk5ZZI1srvbXjxFXLxKfz9IKFXJXzOA1ROYUBdkho3pMyi3e0Gmq1MMtGvGbSXCg
8LEVfWPFqsF4hKUYMVuCWOY5sWbayTXduceLShqumra/7879cASBHQdUeZzhBdD8dokFwGATVw2a
cDyA32m5Br/tYCuum5ncSrAIljPhN8JQyAUUIEIlbFtrPZ0q9wlZ2Wl0hLdXdDCajB+ikYw3x6/Q
5YFHo1oeOSiBQuGBOJAolejkCzXiFscrOjNiTF+2lc4M5NsBq6d9R9j6x2BF2AJEuahu/TKuoVt+
xC2dQhkjiVm3epCPmUz3tyMOL/fgl1h6lsleXK5h7pl0dZ5nqthGRXl/bUAW8u7MI0R82LCKa/oC
0VC0P3cfGqYXr5MaLT3L54qkOn6kA4w6kl8xKdquiJOorAEeLRZggixNmXbNHGes83F8IndmOMKS
fNagPzS+Qm8ScF+aHTqop6hxAMuuBnNaEsM9cM9BsAJozFj6MwncLCJTe13PiuWJkAlXW83yqdeQ
L/rtcVd2Ul2kZFoTsN7U4/1x86TQRlDSi1hArg8wW5GcsWSEApV2RK9ngVshM+toH6ZtvmhpwcFD
CPD0N37qrelp11Dg5O+hQZbclf1IPiWY9rPdMtHgYIXmUQtNT9qtvvL3EYYiT7a6e0ZdSEsSb3Gj
iQCWAqQ4/u08sn0jFR7VOMhj9zyQ2L34r1RQYYuiLuuNsVqOJmxvhw4rNNnyHgauBcmM+G9kdDKU
FDaWrn02V5fLBn4sl0yHhA5ULijRiPGVwHD6TxfrtRCSFDFojhitCrdn+5cM7xv5SB9wH1U9Mb5n
HuXJkc/Ets3VhfEN6IdEsyzOcIenFhIau+rNykkZg56h7qbs5jaafHl8Orj6sZAOGZW/vkIQq/A8
uBZhbKCSrZp4L+EFfGp/412Ot1yjDkbDm0iSimR6x/3c5h04WXfIHnCX0t8TMC/bgIuX6gZ0Nuee
m1s8th4yUCbwqZuzBV6q5hk7eYL7k7eWstUm9Cp4xeBvm7tZCJipDNRbUCDhvk6NcVYn5FGnhhal
g9fFSMxPvYPUEpiBQpw9dIQIVkPMj/Un9PSODhWCthBFackLamsEr7pfC0adMkUbBiej3bsXuHcI
HEKliuNjrBbI7+LFEiopT0WwBXPKPpZ9w/WTSEfgB7N7rza6GnNTDbwC7SjD7RvzJ+5kDw2rVJ9W
MtDKCuTxTjsx7L9JZrd3EYO0oC8lKpYIjI1zq7FE/msLACwAUr2gXM12QHoKlq+MLC8kVnN3jC6P
MEQeQBDUYseoxlKTikd5qzI5MXKEo4O44dR8wqTrhoTPKRosWf+SerZEv3NcXPnS4c3BZKvFTuFi
xhxJ8N7nBOeRX8OgMf1EtfW3AJ4V4wVHL3e0OLBD1Pc1jkx3wtWsMyOI3/Z1aZiO6ikPEXVKH4dv
GAszuEC+QrzOex0w6BG7SLA/2kVzoWaBx6lAIJ3ekLOCslPf6tZJa2hWQvqM6vP9V7UyXluBieVH
Kq7nwB8sHfFRJpjVM0A4oPUnOy9L59OEvf2uEAzwjOYWCZKOfkATDzq2ZB5/Vkvoh7Yx4JiZZPGv
7Eu/fz2u48yV2WUPChVbS3zHdaLi4geM+yxSbYzVgoLgySvw2eV/Ekcs6cd/rI3g4Te3JIyFQt/I
58RAgAup1fr+GP8RL59/ac/ftZ6UbHKWRnA77HrY5+/OwGEunpIQS3hJfP6DsIk6z5LIneNSWGmR
SmTW0VFtiSAlNDLECX5hKP4KzOH4TFfT8omXs9maQlE/T9lICWHi7XISYCxEZ+htIW4NN5O319zQ
/1NIvKLZZJt2VR4x6+4MNnne0RYeRgOm1HYpfuedhGVvPRFZUornS0tzrIux/BzJxV9TggXvyY39
R7Ts9weSA5qJvUgkR5qTOdcLFJr6yJmjhza4587W2Tppu5Zg5euivR7MXHPffHd8QJKkhX6ssgfr
Qk3zGp11SUPeIsW4lwpQWjLHGaqVQ+mu5NOgONBNKJgtrW+O0RY8XGypTyo0eUG0bpF737fCFIL9
0Ma6dbg0EhHjpCai+JLbzusMHTHn8sNLg1avZp50v8JEqTnWCaX7dGoGY3giOVT2I7exFAsakPSc
HDe+VmZcB6rz/9kf7LeEzPPf4m/6KCDvhB8KBRSu/NL2v1N6e55FdkgRJtShSbcTKFgqwb5jrT+G
lXZkqvV3yewUtLzoLZ6oV2/9FB8qX4WAllQEqs1pKECWcQKP5tn/95hGJy6G7Nvw3EZrdxgZVIbM
vajLBWn4Sbp//U4+XcUidNy8pdDhgSvzhGTLfk6h/ZLQV3csIKDhhV8Z8iRxQmRYKDHIXIWonkJn
1b8BiFbDjh6jvAZ91vS6rtsa/NNQk/e5JzD3jvk8HIvAzN6gxLrU6iAmk/9SU2mhmjNZxELbzkSt
RMhXcfqqD5EequBcbcYI/mKzo6wTtyBnQ1WIsqSA7gPHKi9fadTZJDbTs68EsVK0GF4kC3JitmKF
rLU8cMS0mpqNKbixmP7uaNMLVx0pdXA7s0+GqcoaeNZQ+lSDcsB3OF09VVsqrC34diuWWKaMELCs
0JNlvU4AOtTe7/Ynj2dKzzv6sAAV3ImDjE/haTEs1VEX6TFIMXVIsnmeOUuPimx6fLX6D9r69ek0
uXg7O3mt1c7E/9UZrm0W4uzcbikGAxp4KZRrs8rgZNOzuhXc9EjnE3VeP+S7jOwmZNGLBgixaGrU
QpWluExQOlfAiBKGSg0I3jB5yGLXWyrvMxrVfNZRDgXcc51+RTla3WZeghh3sSMEteFcB3wL+2gm
pdhY3KJZg3cNTszphO39GUDIL2onf/V5r1EeBoH6R012pWMOoiRMWrtXzWx1cet4fTQCA8J9Z6lk
NQxpc72E8KrFuxz8IiMtm1wkXQJxRqQViipmmpWM34ttCI8xJY7n00/R5rSIPK6oGqUsSSb4O7r6
cCAelPA/81Pf4mPN/V7TOo1+aqQbaP6+qqQK4kNibI6wHaZ7mmVoPlxtQTuscSapJGLDy9W+c8EK
y1u0FlKt9kmaohFAxOi7jhp01JyAA1qRElxh+HtRPJw6wGWIvHoYopQYmHenYz40UCBL4WvKOB1L
J0neVS2nEZRGV9iZpzk/vT70PmtAxEuQ+TNxtpz/LQ+Im7uf/JBOIGggeKqGL5qGSaU/sFS6Aox/
FG30qORVbCbPws+fN2hXRR18hPypUnB9erpms7FAi1qpcgpvtPstHEg/D4GrwcUn/yzUn/Wjf+zM
1/MlUsgJ68ZFgYfvB8WnIJwrZ1Ckxlppq0uJlLtL2fLC93ceJ+kFgYDcDHYHpICMkyAKWq9HtWBo
yiHAUB0g/1kyr+srXSfFGU8iYxHhTttYEOn84LcWcd9RZTqZz9b/5ppz14rIeNVXUk7kNiCJB2eh
me3RKngVzCmMV/dD7qW+yNBFmHrqZpjoIfbRC/SSNHgYenbnRsfHjJWfvyFBuH24UurNa+n3lwuz
Sbo5vSY4nU0bntCx3Dt0JSxTuM4j0hwQSmxqd9ikDQUDbtnIfmwEtvpaV9kIrDYNotr904dXeAoq
8ef7AsA6M+xFJO60MNo1aSFE39SC/xB/Tf3J1KaCO8DZ1sYjUjRaueonRIuFcJfGOyaXsBKRSDJJ
OrYWn06vS/+D0RbpydZvmsklezkhIb6KNUGKvFm3ypt75qQhosVLSnqfje33ndrtf2Lt++EKjPXV
jwwTQ24NKYWeamVNr5Yt3K7AYcL+1KuQKTNmpQ8erpmuaAcjgyJTuzaJJzOSHi91oZf5EzYaIb9I
qj4v2g03EEayvnC3yfQlbmF+5aCOH7/pxX7OgSW92VFlhsZxkDR8gCx57Gvdd3WXTGKCzpqn3ctn
Z2FddwgPIHBn90wjc38WgsiUCZLe0MfUCAjZB7NW5DVdDSaTAKDX/n7AWm1xpFeLFuc6PLDP5/Bn
jIg5fHAisY8D4Jybm3yexcT3xoEkRrC3ERiwD4KmexYop0MUwJgk8MFdarJQ7z70U2wALb4WAciy
qUoEQJkwl38uVbgJYHa8wVTMIm+RjQVs5ph9TvI/ABO2L3GGBCgU1pqGrWUwAPAfW8o4PIYgXGob
1oyqRpFd1xA5HOTh7N8ZosyueXef986tE0AEMQspQ+XDcksh20I89j/TJ9vKSwSrocJ5kJnqjWw9
8BHfcwGGkBPBgxNgv9rV1Q11xsvLPTExPGef1A+OAfOylNKSQbCvVS0QK0et55y/937AoY20tc6v
qMsslX/0DahaPaw1L24+JFhIAp9rtfy3vUyk3r5xMDEkhOXZMGKcboeYPMHuMXwH47Vn/j37vxfp
iI5/L++GRICE/o9RuioNilkWtzl/Q4x9bB8kCbTx0F5bYDnkfH2nDjFxv6EWuO0ItM3PZwWJ8Gbb
9XRJH55RETN5xa9XSw2HlI+qlozOAg5dsnzxORe8SOvBFS0nPumikgqOfZwSEdV+/302oVO8O1tN
aKtQCeiab3SKkcQFBVbinJNg9Nu3YYhyuVyPD5FrU1ufOcJgRiK9LjUvcLKLbqBPjKw6/2DjdNk7
MwvasQCVOtUpjpKXVhNA8mErHTLxdakCCg1zIL8awAk45elBQAoydaBpVDx50GLm6MFQqJomChwg
xin8izFp/RAOss1waJTWvsP6+k7gUXnjHWqNytqC9TTZ4y8dCyJh9HxOkXYq1OUc709+t7vdgRkL
GoN41Yr+BK/5lfNxX3xOEbPr1xOHScn/mIDuqUAqOmpCzwgjYxo4l0w1wsyfCRnsWv6CM/v6hcPY
2Yd0X2S9HH8RRpbAFqn3lL87M0l9INvZeFRvllG6/X9SYHxNu1d4S8TKH9AATPUo8O0gNWtSavG3
vGW2HveHVD8YEdi1DqFifBMHL+7fkndumUCC1SaP0jD68W4leDDg2xjHkMSP4MyjSRKtg2Vz2LJR
p8oC5sOxj7arhx7QJq4MzQD0+Yu7YP50FmhKp8NOtQGUrTioygx9TE3g3icxdGM3yJ2AVdbQ8wTN
A5fv4X87r2ifwrCckRXDhL03gHs+tQFuV2u6K08KmnQEek+1W4gtytepW7Cian9aXN9lGfVCGIQT
x4FgibQ3uNKCNlsK1pURpAHIdRV3IWKKK5KSqkSA2nzYFKb4kAzUuSk8vJPHLYQeFTPzs1wztFU4
uSxwxfdjwBy9ovOAgQZyYJuMz/XjaypexZvWuECIeqchCzu9h/dSRKrIh1xXiAaamzXKlCGOJtxj
+DoYcDfxhZ+7WKCdmOoTMgtWHx4HC0IOgWWy4W4mLQgRQ6HCeklurxHmH5biZ5oHUT8qcCd9aWGC
bLIUIlVIYwVLN7dpJ01n0ZYUgP8ESkRCfx/Efcvp1IFLH7VTTXkWngyBF2an77091mYVQjf7EvPO
UINz2wjMrKcy4XT9a+MiqPOquz1Oqf04+Ig3D2bT5nX1NZrvll3zZucDiT45HLnw6joQc7GhPA+Q
WwBEUHaMStmf/hx5fjW553CW7vIMVqgooRjXjp3vhosYhU944J+hGk8fgjPGJt2wO0rZBCukHfoe
Avl3L/7IyhebIa/03JaKT9cClpqXWBAl2T6I8uZpP11q3gqo+CM2l3K6l7thN1J/KZ92LE8bzePC
sGFBW7Sh+uZ7JnjYN99TaBYpFDIG1rCfmuubV6q0SfzTleMkER/75Bru7GTsGb1vgt97BxtX8TYl
B0J/eoerpqj7AkmpwSk3ZbzSYrN3KyOwo4CIlg0ZkKCJ6OV3tT5FAoh5gI1thU7su7ki5nvPq8ME
ZO5xaInUyqvPlbf9WzDZT40CI2s+z9aaZT4M/hQLZyriPzs3tc7HzJbzLaM/sgoj3guFtNeJpOWc
NyNEQU/YHjQsUew86kkqxW49qWqfhhXklhnlQ7JQNfh5FsNrA3qahCXjWMBVscrFcvOfLdJ+Xxxj
MJ8G++ILHiOI8m/TqLAJmofG0mH1BKwX+JdifUH08qNuVESswbMKd3gIdXYIwNJd8kS3v0de86wr
xKDsjMt+TUOFlmiAz4+cNqQE646Rdn3oqXLgziglMKkmpSgtOZF6MudLBDSzT45eIzUps2sGCShM
T2dNvMXfSXbULlpd/Lhar2U/dHmi53h37iY2cAkmaxpZESPCYqHagbgNHvbnPjhJHdSWoYiYxTEt
lv6+JViI8e6X2xcz0hCj1vfCXkx7wJ21feUB5X8xnRqFG1/v2NenQcEtA3xB44i+oa7o0msrovx4
HG355i4vm8AZPEb81/OPE5LnAXHOVDj2myyeAGe5S7g+YWjHEbEpgq/ySEgbtLxJfnzkdXTcMzMP
AIlU02WTBKbXxzHb4DBqk0c9kBgrTrpJtPPbEa1VJeB7ITUUTVbgDjuuaXf+rgwSBTHBbMl2v/gA
fHGt2YjOJeNlV/X2CC4LRP6os/sFT+JoK5ts+WWhik9qVti2UdQyY86W84vOd3+5zMuySMDLdFQA
IhIB4Bm2guqdASIprPtYC6/ftx0LhZZIhU7XlNddAtCzVh1Y9U6OXH8UGzw1Eg564srO6i3x+8PU
9KxEWxbW/4WJhcKbiQXyCkPu5ebL1Et3mgsX4clQGQjaGKC625SVurGchr6RI/H6uC1X+N7wPkim
xPK+Yh3gmT2EQgg0eEYAGHFenZa4SRX1oKRQ7cy/coU/lUAW/N4BYg75U2mir5tnm9O9R7bQ/hVB
cbf0ewQgEb6he6jx+gs/DFdWIoEeyg6W7MBOglFLhcm2mJ15zCPySkX/GE8oevfPWvvAJ17QFi8H
UDb5JNmJ1h2fUjr3rIyCpIWsHcZU8AmxkriduGjVzbUM2sq0GbaMz8o1eUWxVefSVcuCvmbEh9H/
M7kXbPNT39nQgJjIKgVNwBt81Oy8A9Lkl6SSAxENSeDidtBJyJiYtV+wu2/m29EKO2Roq0E91yX4
sIlOh2uFaijHIs2siynIKF6FKa9wRhRGzeOTG1q/SkRzaLJ1edh0sfR6B8NXNcRFA334KINYH98B
8xQh4jTxYDE7O67ftlmJyt+IiR4O0NEtWTJNWTx7+tLySFzRtuRfzBpYy9HRMxFCeGB3PfYpBfME
fRGyJR5AiKu63Wza64kUfvT//D63g0yFB2bCP/01sLR0Y7I9/5+WheFzXhmXsxOtCgTT5INECiJQ
3e+WaNtHW7zU3k7dRec9GwWcJ5WPs2LsZbjwkG88qOC9mQ+4qR5JNnawWHauVSZPWivdN311SjrB
IYZJCAsiV7SVrrjT97FHDRyJp9x1PH7SmYvUqyXx69Ttn59YF2Mq6nPKS3ej5GYquqwTMmWQ/AVI
KLcMN5D/FnL7eG1ViEXE0KGnlcVfiWAaJWNdG3HENmn22aWgXEYSrrzDr2CLMyzuajEDLBFpkWQi
5py8HFbcKp66b+cBO67RUXLNZpjb7YKCcHvkekpqUlieKgY1p25UktA+xxIqmi+TNmladu36lq+s
0Krlkg2yRKxp6HVv2rjNrJfwE2+dHfMfJJPpj4TAj/0OdOS8bxWHeUpR22PClgHRIjBQX+XQlRYI
kAagMFQ6tR1cX/ombmxGX9OpbCEL7IVzhw9NzgUvkfz6Vlgj2fyYMze1CTk6egEF+9UpyUM8YNb7
FzAlNqUkztpCKwWonOGrl4D+pFxgfekScOZE7yb8bvjEPFCZ36xzg5ZXFUrRpenIWvlrS04Vg2Fn
0bICPp4ByvUek2aWPyN2lpHtRGcspoNmYY3XgTdHv7SxN4SSrpV94YNkHNAktlUvKZuX23s4aa2M
GqJO1DfTOOvXbJ3PAKreu++qLFc7qw1a/ULkO/UVW9NYTdLCLEKyXw/fkkiRZdIa3nB1zJrTiq8d
bbDz+JYkcxZCQwSZWSr/aoIddjTkys9DVvpMabs5qo6GbTgFSgZi58OqWfBXgcAlAMX5hExH5yIl
e4WcVLrhooe4XdqnCHUvS34u0Bdw7tShvRS0Yosam6SHu1EVqH4JC6xCpOBsWungoOnDfokb3nG7
2O1MS62xSbJt6SaCMMp51vaME88dulPDnUucIlzSZsOVl6EbcxaIyjlkNmORdeCgKGa3rTVx1tt2
BMZK0bklfjtUjtFab2Kk6e/p7psVsgCd+G2tf53DwTqK/TBemHi6YD0tMqJSCq6us/MIYwU7/ZsE
AJFonY27sDhlR/pg7Agl+jbx4HPSELKjpAAGWQ83o32QS3YX+jpEgmtW+ClQLQXfZgdgEv/lZwhO
J9u67HzJ6iItIanDO6I8hb61D49Ng9IJDW2hhjI1a9RWaA1+dunJxCuV9LxSCZXO4eLEwVZb8YxU
I+8VmGaHFxWAGI1fgcuxPkdrCo5XpBJRi6BQNhR14szekGL+0NXyHB+xm6bW205IkmEnwffxnjc/
a3B2RtRPNJVHz9J64EoKJDckhjPzOmS5oRYvhj0yYiGjAeYPhFZ8m9zi6EazForpqraxJF7qXfJA
L9WnKbivNu4o0yodi7JZgh16vZfvdTWZ5RMPfCJaab/MjQ13evgHqaLRBX1uu3xNPyd0RObxXZ51
8k1p84ZSptol+koL3nJtSQ0a2pkl3whfLyjdYeBkNykgaVXWKZ1hdxZYZNURVdMymt2J9p/cTBBD
IaAyPw5tDUYcl1yDwrCpbFrTS0NJN0oqL7JjP0we+nBLL5YBJVrjT0mEOsN439QTXLykqwenTNJ/
KkCt4XKr6AzVtJirGTXca9cX4r+HFFEmUnmhhR5N+3gIMmHBgIrZq5CixMlVT9kCXvlVCoNQcPIe
MYc1sJg8qFOJ9HtooNmZ3gG0u64sTYr4JllddM0Y/N9Lonmbx0L+F12rH6h1yMqXJBk5GVVn7g2A
wpET4zCmteeHi6PR+zIxhK6y/P9nM0kK1xRN6agBU6weSCPeztYuoL6Atj3ZOFggbJDZl9TzbqvM
xv14FKL/TD9ppGpYyXxk3jVpNcK67S/Z4HwqIohxaUtwgk+lAucPsHB4AYbAxn5YJqa7CbiCzEQE
ftsNiZdeyeEWSRtnln3ZWAS8wUYq6y1ikcBGymufRXLEtnymfpk32CC+7W5gLmL6zSoPIwkuktw+
TIz/XEOKnPOUL95PAaGz+43qS0RAy4Q19secp/U9ieEBnshZe0UV1zHlwCZlXVPe3b064PJzuxfw
WVRyeV+YqDP4Ypdg1BEFxISGcf+0JHuxYxxOMBcP5Zr8gO25wZ2Ki8HgO9G6F+hgEFXZxu6XCVmm
I+S3mn+ywwcWsZ3yD72D198NyTBLo6uBbr4surdGvvX4tbREAQn/TvrLuykzXbhKyIPFU45IJkhC
ibg/ikbKeXlw22Pr3dGLw2CQQ+3OeKNLCqPT/MOvxMl5altwLJxu1g9kKAkc8zB9f9ZcOpE1Fa2I
Z6YyTxrsSQakaOvDAqfJ4aPK1I7CEh1qYctudgjfJ8HEDQaf9xscHCi5VK3vQmqWbMVFoF2B+qE7
lGq7T9L6XJNk812mAHG83b6K64QlmkfBflr+vTxrrY3sieHowjuppmFFPDBCp4t5RyKBJjmO0IcE
lsTTd9hHQLGdJBuMjoVzsElS3nsXtweEyLFC3yWdV+Mvia9M07Sgwf64HkYVlpwas/iwcUs7A9Qt
K0eiCExXGHe0n9aH9AM8jGPXrd/MQxGypfHEtajUeK1yXUXS+syxUFRsFYyfgkPKQkA56oCswClO
PO6GYDLd11lo0sk5KdtYqfYYM5HdfvWhG9sHm73VXKIcq/PrLT6CUbVoJNoiMiWRIPIodjCMiyDP
p8Jyvans4qgk4EDQkMWHv8Brb6bMkv4K2AMy+7H1edh24+GzpNuUCSskJnuLorlMCab4jt0LWPQU
+bXtSd85yKboORwCtwdHLEKnvoN6XqXAsj/PQ++zMxQfZad9NQTgzVvOrIEiRn1FnzB9tkeAmc9V
i49knJR8TIkSH90yviPIB7A8YDmBhABqtu+KhfcKG0wGkl9eRuXO+277Q25Edf4RZpxzmVuBK9ue
dc73Xy8EbpAoVDUn15TJRuDjOMrzv8dccIaFrIlwzr0Svnp5K7KFsRhKcYNagSK262sNUjF1IRpB
4qVUHxdQbHS5wHIlaFzI3+mEYesWJJ5iPr8HrFa3OWoA/BH1s92b9JdEs/V78eI/DLexkOBz62hE
kis4PBcdm+Tw79hM+73y+lZEYr9ldCnTWeJ/DR/fOeWU9TdULCa+xIoXkBS7irKgnR7mnSFOJjN7
Lx/saK8oERQtplodrrU9a4ltQbdhAQogU9O/5AGY/7RLYH1K7aKQauQJ7R/2pBn17JG9ockFJMKS
STYT0jq+JV0G92BTg+BM6CTtvZrsr7S+s7qzQSlIYxWLnb//x2f3zQB2FZPtLJgTkWU06BigfNMc
zt25mgiGeoD5foK/K/XvO1vEk4VLJveOuFWIxSIExDQSCI3y8TRIujXyNIhZDYLzkoHkO8tLOf1F
DNcOPpZV6SyhuMoIGXGql7alc9Dm3i+phe7xKkKQUFJXzKQzWv865r8oTQxvVe5t02YoC+HzOVI+
EIDPR5GeV4AI6KJCW5ROAQzzov5EWeI15OME/gQFX5wISu3D5hHlg+fALs10qhKINRmfiwZQNick
jyrkoH6ieW+ktvf7Q4oiO5ilfybk4yrW0It8vpKhD9MZbUckNMomLdq+dWxYvN+U7kVWNWAuNMEI
PxUeLG7b0U0+ezx2OCN2Hao13Cw8vlsuzv2m6g+S8+IuSKwIclkXfHBAxefIbIwcv8faOFNQ5XQH
Z0LEjk+24JXwgdTnseujjyqXqO1ryLooC56qH5xlYI3PU72yX5gpmq+GKZjgKLGKwdwj/X8X8EvW
3y6BiyQvs+/bJ/1WJTvimpiz3hN/NQgh5J5Tz21hADwMy0erW8JSFyOjR0iTg9mexqO9LtT5vxK4
iFvTYuYY/jDPZc7Sx7+SM0IRKM8UGEXUaEoKl/iD0hLvITyu3qjC2EzBDusQE6Oaser6XHenB3ye
H4wf9VvRSY0b5wtTvPRqUJZD8WdK5yee+FpToYEWASuBt6GlHtezHo3zEGwTzBJWxPgNdzGIdDpr
diVUCKNQ6AFrk6eaKXrejzs6S94kk8ExjaSNwGr66vUwb9auxAFFSKsebyEkdqZEb0sXDmNeSkX/
RfsVVpqWzAGs/5QN/U8Z3ND//dFrGZWBvolQRGUDSnD2cH/Y6qWkhS4ElTJPhbpk3zeh+T5Apb0i
vHI1diYhU43rdLkrx2n3FBTgs5aq43lasauiUJu9H9TfLqoRSeiTwukIrK1O3y1z+GWM0Q8ybN35
ZxXW7YIlM6xib2a9uxl0NHu8oZ77Nq29C0kxSfILX5v5KyP5V9IS340cv6Yrh1YsUbX3qyMisnpP
nsXD/VJQPApwOu2a56zzwbuuc4fJWrirZU7dS+x2BtYJ3sRk72w4xt/Q6wb4at5OFKM3zwlBl3q9
bVeANnm9u8cMMMmlSin9SR6zG9uXcw+o54ogdVrheBuIMqDVcdmENunna4A6cNfPru7pkJh5Qs2f
8OQUXQGKPT1ty/GWX5Zxa4R9KEahvtqafBX0oPO/35OvUpPRJjDXGedpQflIajMXZtsekk110YCn
z3+du1UQiGNxilUO9+kAyzoS2lUZZrJyWo6l1Vc5K1i17LZ8hwjNkjwrjFiAkKLI11Of8b8m6AuR
kpe3/KImAEinKbrT9BbrMZ+zihJqNItNUTZCJstKiJLYFK3ZM0qpWXe0vb3yeltV7oOtXJQdmcjL
QtbTb1ZVIXNCzDq/xFcUC4Q8mozoU4aiWje1yerYh8Cxu9NPh+XrsYnj0rMtjzDXk+p/w1rahXxC
JuKXEz9zX0JlmXox3jWU6bcB47qVnxx39GcTDtLRo8PxtKxeqbwWduKCUa0pFU6Of/LhoFo9GID5
XzcHb6GY151XH+XfheL8lOf3LUnwhEOlIZ5rOyVcyAWEg/axf+y/eJr/tAVQGh4q4LKQTKEQ8Eer
pczDXJLBE9J+TeHfsNxxVTYzLk90jq/FVL+CKraIxe65jsQCdS7fL28aQAutCGn11n4OXOSSd2OQ
zmugq8TGO0g2h+VGiPz+KBVhF0mlKDLmt7QMJD9A6h6DBArwm8OiqA0084NciLxmoqchv+GAW59Y
0eON66J4BIdeyNNYYqxTgExDlDpgZpR/KlXMtN0U5NOTCoweLJ+cM3PeNZuEZHRcFq+1QlrjeBWn
2EGfKyHAYmcg9KtWk0XlcVBst5zGTtTA4AK0OV3m7cK0djHjwd8Ud+DGwSj+z7xw5Bcah7Nr+PBQ
UMGnRLlP+cN/FjT04LKBq2i2Rk/SPwvcjRiBgTFEkZAr5Ae1gszhwn93va0UWRIY9BZB7zAR0mbb
LHeFWna//hUzdyXE2ctAkwXmXi+OJonWNd9vNn8yEfoF3fNTOCzgIc+/IMhd0B4CaoG/ao2ZHXiI
3RvUqusj+Ioa9t8oIBiAHrthZswaKy6zxtFVZdSunWzaGs/Cz380drfUC0SrtqQYLPni/WUNZ3mE
w8e2boQcG/BfR0lc1OPckUfwhNojvyJHN1vYPuUgJLQ6peLs9uilxAtkDbSQGRW4h6fquTVbh5Mu
2yz89yht8/xN5lM1bdpH5uFPNbJEq3CCrBBctBC0lWMki1z3NQZzDiy17zCHo0wDeZt30HSiEcT5
eV7RDHK+Sgmid23dblqcxdIjcFqvNs0+B3aB5Zftn5ZpfNmGh7859XCk0EgBo3I1WYIMN8efM/u4
bx6z77qpaxuAnBarhBrDgyMTlTcO9uyX0x0EBIg4o92QhGXXAmfOg8pOcu9O5XAM001iQC2Tcvez
7bA+bNLYb0WVsFEIIisSOLib1ibUm3i4rUM29dj+tgDLjXw5cLuQRht5O4EA7avbjWUGhB+L581f
fQW8kOq23vF0KjYLf3nkVqcvnhV9efMJKoUOzIqX8LrksuU41X7HtOGVeRWEgvG9xPzgEiOcfbz6
dxLiajNHvEySiKKfRAGAXs2b4ht9PFsbiBjAeCJLY0SD73BZ/5zlmL3HXYKZBCLxgbdb8BAQAL1L
7ulIpm6CJ8D6Kos2pwYDFHQddEIIqVStdKnEPK21hwREw7gWaNlMTf9Kl319bA/mzQwtz9FnDGsu
Gp1GqqseeSP3OIp83qfP33O7mof4BQiNpc8Tuj27qpNxKqC166q11k7MZxedCzPuwF3ceGm4s0D4
d+UdG/dWDFtnmgovsIGOi9b2O2r3+U+5vpZ+7WLxovQAPgry1WlVmDc0V3ifdOVVj8WN64B/wKRK
LlWcY1bmK3GZzLLh8YzJzC3hI5F8neuj8QlnimPjE6D4M1rOUcs9omAejTnCCKb9PsuCkKOoWrt2
qHGX95f2BbLGAr47pBt7D+cuopi+S7OJFMCrzvYmkz1gUY6XH2QfgYBupCdZEzf9HTy98sRRKFDy
dSr+Nu9Mev54VKeUqN09WpsX92/+B7gunOz4DGF9C2Q/SJ4OdPLlE2xPVrns5CoNCkeyoJ0XDAdX
bIlD8cQIxHCCZk4pB+eO6R09S6PsP87sWuccHWicqwQvuZbBzUUwZnbHSEEkVBGENPW4L7s3CIIR
VJZKtF0T+TUFhANMaqNsaC4ELB3duDnO+OF27I3DpbzULgFDJYMbGLXf8eJp8Yc3Qp1rygeguis8
JRJP5A0YwbTJnqcvfV+PG9KqyWVQuMrWaDumMS8/6hBuL0KL678v6SlR/4xqPtstQ8NA3K2mlsWR
IcDA1FlfgR4ehXPvJG6uRGGZCX6MtoiUlO47p9NrjnO/yFhJN0T+cSsSaSxISqTuT/2G7XI8WtTI
vZj7bLp7gSda3JIABCgm22tCmLalensSpVEYsQmeRg2H4H3f6WeK7v1LoG6px9AEuSwFeOISdeot
lrG4AMdRzLvE/xQhoPEYdruKkbmHAYiLSgJDq2dpTVn5z7zBJZ+7NYMQ4wlXJC4WUg8D/vzwsvtX
hFQddKO1awEgdSBAbVaC36RcYRHB5lHiqdKYfNa5AqDnoRNoWUrqUJL9NKtoGu21qJjz2lAjMbkw
Hz1PJOEsgwukdegoiArtTwnU++ZerjWRY2DOE3BWwIdg1jOS4z/TcRD2MiB2FJi/LZ9Dgkq+Absg
z/zDdZVEUWM/GHFccoMzurQQXRFAwQlp8FEUby0wImKwEIgNhAVfFOWfxADzaGOtGEUUrojFJmE0
YZYUNXpM5+vOzTTyMPVNRlUJCoJW5R6uRSti9aohHYhAaKmMJbJ+Sq9IHoy1vXDtDt4vOaNCwKvs
T4Vr1Z+mL4xUqx7RcgfxbyxvVAIhQeKwOPNOJojOA5l3XKVHfj3LvoHxuXpork1+pF9lChTuYpJm
deAG/XQi6Angv0UrxmwnRsQ84ZryW7kyB1EvdP0jCvY393HtS5GOnVgn0Cd3DYQQwnRQmeWzFnfb
s61zsy9jMKj7BChEHNhoPg7hKNGodBcZRhIK57lXYUSi9uw1UBF7iNsE6UWRdQM1iREnWysCs4z4
rkd8qxfsEw7Ad08tUTmJWXYykitdqEMtjGFZiVBfYAQxOPcmDQplo1yB36ULXa4ERwAUbGrwMwO2
nHe2YTILs05sVun03xarlEu0lfxjaS99u4h87BmWog0RSWwU8rjrnHoC7itGpuphVO/xH0YS6Wws
RMJVJXJn+Ahmgjkivxykdykm9FBr6c6O/pxVYPcxMAswuGLGugX1fuNZLFM0LlGzIlsj5DmOeZE1
345Hce580d9aJJ/u4ANbJoqhxP4oRXWG8KALql6kJUdToJSE3AEUkQtQqkvPaOHNK270tiIHb3BT
EzKLlI2cRUs3XxfxD5uFLWGR6N4SyLfhQjBSOqvxORGM/4tPNqzx8gLNW12lTidXBoPXNMcEpXGH
szzrqtOYNeZwQmijP+IejRnJ+TyqbX7RFrO+J/tiAdzeN1rOE91S2mCAHnbdGlrxx71oRo4h34jd
efiiAtcsF+irylqYMkJCORimCniRCsuFAWmzYlGtBX2oVEa+G47zoD4KJsBGLvJINoUw6aKBzWFK
4x46bvZ24Z4OeOVeiCIuCT6MmkiPSEtQQtZnPdyGlH3hNVsRcNLiUmlkQSyqup77vvDPzJ53qWs6
OOHsbmiWLAncf38lLpklDdlALS66cA1uMdhWM3RZGp3dcDLj15XpCDgw4/oBSry4T/R4Cnwss8Ov
AHJ0dQeXeZiXWQzD5qDNaF6hswTMJ4PdKH//DVsfdQk+5R+9LjBrK4O5ZXjVbRJ6TwuoIvMPh0j1
nbCOLJFlynvC0SNWB6mnxXFXt58ZGZ08/6zjCcz4oUmq8rjGKvMWc1FGuE+XpKoXdofAvVurk3Sw
PmyucevDK2tFy59h12B2uyRJQadb3TEHttUEPndH/t/qWToVsRdp6rym+tuF1kBhkSGIdKzLiiz7
XmgyzD6Y1FzNoSVzn+b5qYUbRf6j556KZUlNKL4Vh0DhB7S/6hccALokZMlfFfNGY6FA/uIeKm2K
7L5D1HxChaC9kiAD8q3yLmEGiELKGT0HyOrMUKwaEfqFJW7SBRbRUiJ/bO8SEFm4nu6Ky46hKpcF
W9ZyIX+/zjRIHUb1gKZtsJwMiei3YdxO2rHax78gYtZGXvGsrEaL6kGS5G8ppE+DyrJlc6JdQuaZ
6237zZffksSORKYpkmVu3ymQ9gHNrUEJ+sUbfJjSnCytTFD9/ZGZjyTcF6gxnoz+NM6M8+ACsMWY
ik9DtG8NEczWopqRCgJKQMYy7W740IsEv5LsqPeam8iXIdmw4/xP93R4kXXyIjmnWgiOuWXUTKX1
nC60l+F7jYQMRLWSUfAjPvxkZXUMTpcjmEhwVoaBD5bx0YlC8nK4ILams/wVyiSTORBkV52DnIT2
idaF7JLsCDW0msc8Pf0KA6LDzgMeBAMDnLCHSIIfOnGv9CnhEQ5a3iEj3Zy5lA1Y5JvHrg8VhHp5
atxmqZdxB/bVPfHPjUqtGzkAtoZ/osNtSAqj85pVAUkmBDLAR3LSj4u7QgnNixiyLPXVT8cLV1vZ
O0jT0Rd63ElBr2OOQ6wI4opXuMDufE2ByGWFcAln27OgKNBGykAVW+6q+2hnPkEQJGTIBn3gpzsA
V5eMpUdyWpBP844dSrWSv+xQG5QtHhdNyDRrzCih8HIIcKu0J5OCN2w6nT6Rp/1+ax9L+Jvk8RE9
Fjk/iZWe6AK3qhrNJkbibR4CREuaNujmAlY9Pmg+x8QJTR/U55QFafJ68wtOEMtSB1PhIKLuCCpg
5QRlIqLupHEXREM4BqmFf5JoSeCjprabWdPZoNFgBxYqvoIV1OkUXL0QjL4CpWvqvHu1wAjg6LXw
zPRiKKP0sUPcYh/fhJz9Df14ptK4df/7oXv+/eDaGpE+LOymbjsK7HY1/lWzcmUmvrVL1QFKJOFQ
BX4TlYFAcnILZ68FnNF06d/yM+WHMl0KrXfw5bj7XL1MthJS0YqhZikO44xWSQwl5cZ7Bx6cYQge
YqYUxBqz6SvgoD5RjnIhQbDO6xluXzTInlG3aP9twfPVM5LMy9mcYgXTI7GSH+VX/vNucRdezHjK
FrvZj14uA0VusVFlL8eRyilRuzFWU6zDv4EWPlga3AWs4tQ4vfiJvf8GENoBOQlIxDfQsCdo3ATa
6KgykBkoHHSfyqIW//7ixPcfbRpngV+DI8yxAdgsg1luwJB0l+Z5VXFGwOEji9qxpdwZprpTFMA6
U+HlRASMJ/F5CKgTHD6hcCH7siIJjLEz6DpyuW+evOl+Vqef7r2VPjCIloxowDf/KpQLl5xe1WDV
AyH6TcSo8xQpXXDCFoyuq2hJiOHELqlPnyHGNSJpAT4UHP/WOgjmzFUcOMVJQ+ORaBL6QFQUHVDd
/ZWJzUZ1V3MT/2VZdA3yyO3r1PBSZjRe/wkZ+VzeucQYblG+CJ6vQFMD9ImR6ThSQfPtCNTNAIhz
fiVPfLEABLUNIOhwHJVr9fyrkwi0N6PI/4hYxFemPpgQYGlCCGv6bJ7EMS1m1YL7C0pNAnx1JmqS
ZLEpOk+zOxv9yTbZp280lD1bO02TqzBheKrqxTlmhjZdXIctkNUAkw+PWAdQp6ZjW2ba8v1ReB90
7h1tLn1jYcyhY93L7Kb79NZPRCs3/qLitMO83OZl/wsix9A8vQRM+sjDe8nDD7dG849gXJL/Rjj2
MUH3gj7GB0J1vLP5ff+7tjGNRiNDaj6KhpsKd+HRybQEHypJ3uLHUQmphQk32b2ciVGqtVgDGaP9
G7KxIRZXekceklwsSuiEpdxNNkDlm0jjOVtVFHpzX00lZhm08xcWsctQJMbWlSdW4isKr4TjJXv+
HzpD02lfNB+H2X3mxb+QkF2kk4XD+m99jNC0mqRkrD8FuFQvy9S7ywQG3q6myhhaIOPCorvPi2ss
C2sdfIMhhvnCho5/OCKoPqWOA+XzA4utouEzJMh0RgOrTabZbFJgdTb2IXxGsfmCmCRpfSImnyVF
Ks7b9GoXIe+NgmBy74t25wOfrTVowRkYzNOSnhwq55o1xavIDG9fHSQ0UPrtJgWeEUPvGsamqSdO
B2S1STWBA1y94IbiNCEelgX8udR+qc51/BbT+SpgXZCqUx5gaOkE9j+t6lIWBuNdK8OkvTe25mls
j2IIWG5sbtsB1hWoR8Aqy3zvmQjl4SOR7h7Fn8AewuKsu99vKcXMIssvEyoSvr36DjPpG2aKTFBE
snEa1pgD48qm6qe16BNRIGSqDcUNJmqL/OPmFNsyxG7Ly8S7ogszBoGHZmFSkS4hTZfX8Qj9+UrK
sMTqHQRfrqe0Jq2D5Vy66uIdhP7Gxw2skyKwS3AdnVuD/XAHC0j1MokjSDQMqRczJLoRKxWurBC2
CWWTRvzvaImxXivmUr/noU9mm+yKl+wSLFGo1vXXvJF2BiLKvOgO9si8JUGt9WZ1YLNAIfOK1QqS
H1uR5Vgnf79wkg1tFQ64SEUj42k9g5ECnhQQp6EDSohrIfsiIu4GMJCWLhmZEwneJnDU9klclZO7
9XeC5fpl3DW3IkOaPgQRgYqiMGqOz1gI4LoqlO1+QuQDxbchB3bBrn0+Y+BXCKNiQ8Ucxdi3vmCf
DgiZsLaKrnI79P6U/dLYWWTkm7jNuxLChF9chJlLb+GaJPXWDuLU+cU/b102hwjYI8hyT09hrV+x
F/ZR8HcmJHvp5c2V9tl6P7OrH9TwjfBxa9m4SC4SyZcEfPizu4hwxTPfepzHFm/TtMG6TYGtsd62
cPpdA4RC/d8s792ZZRyvS2y2xS3mNIqnw3qqBR9zWFwtYUPMWExavcld8dVPmHzRx0BhizUA9LvJ
EMF7v0lRu0AeeIYZ/MXTE0uILZ1/eGSyxIZAfflA12laik0x6MuaDVusQojgxwoSkwTQ8uyC1k97
+aNeuKOf22w3MOojWdVlVLTuKjJwudRCiFMvf4+KV/iARb8V8od2EvAkO/Xj8XxPQ57gae16eIq0
lB5CfkhWUHPmFIxzvRFNQC0zWY23GUhAWXck1Qc/lvap+SAtydUO5zYjzPyCTQJIDPKNu/vo94bx
VJJ6lGUwBUbFhJb899mboSf0tEVYHQwkNO4FGig1qCQ3YnAvMBe6FywOUBCTz2ivLpgeQZuatMOf
eHxI5qiZ4/LXxUf3h7LS+Gvy8KugtWbvYu/puzfKMXuS+NjZapctSFfqVINBzaweWlTlft2DWfQZ
9wWOIwgtc1KFG1xxl9JY8CY2zK6cYtZ9IofjYMEe6tprdjGKReXFQtV7mMfN9VKRk8Kog71216n6
Uqqm+/QQF0LlNkiHJPQMffa8jvEjJ/c6F1rK/YT9cFBE4TwnoW1kGtBdTk/odtK5k0M/fgtczlKt
cG9p3k4p0UIVejoD4c8YGoKMWBGlfARtXhE4U0BlOA+mLuYRhuuB3WLB7Qub6gcQVlQv6iEb8Qgr
v3Luj0UDHOfkta/axjmgpBwO4gKuNW7ZmVd6Pm1bkZb8qEV8RQ5E/cunCDV5m0MWQQBacmgt6wXV
y06YZ6Zmk1hCyzBpr0Ru1dbQLkF0VT4s4rrF6UE4JQnCnn4DPLmZfrbtGzp7YbM2TKly5IgvJHWc
fjQLuiYeGEnCxupA/SvP4d7chJM33PMgzbshc9oyQ5SRWPQ+Rhu8PWjAn45iOd4Izbv5fWZ5VvsX
AWWpV4MPincmLuiIZ9LrW8X6/0y0XEJ2mPsawLRNUP5hsJAilOnyxMOgvJCusOpnv6EIuX8P+MIm
dZ/eF/v4BwXb0xB3ZDd43/c+zvFF2FcUpxh6xleuZ5acQTcexj+/AwZSiISryAy1Vwdd15d/Ld2v
rAaKcK2F0YhsUuw/6iSgYhfZiVpYLNjCnrFwMU5hnswwUQBQWdKaV5ka+QDjpoJbjSuEdjZaOrNR
7g5+ta1FaqtNm1L3zyYrtL0daAAgC2Ow65y57cdfBtTv7WfYuPwzbsmOI9fwJdzsvtTe36njuMUW
zCVf8QWkXKKfB0eWCGeZ4RAsj/5FYI+fT6i7eA0XP9fFYjh4cP9q0WCtciqoHpaFyMxM6ei+cQ9m
AHdqKMdJNCpnQDsXs/K1HRPbajOfusSGjJpuqhMVTkZIYyrgrgLlpreleA8vbVNKy2/UyL4HG5ah
YTbbi3/KhUhAcU7uEvtj3HdZNhdIR+GMEbivKqgRcreGk8dLxm1k5DvUiwN3KvVwHmQ9y5rW04Hj
4VDnqPv4Rt38yQziLDHboz5+1Fcx1neVyUOgr2TBf0eo9pYhY4lOUjANKF23ECAfAsmNNIJJ+zNn
C//7uLj906IKU1IvJvo8Ctxlan/pIcNyDxsduLerk6jdR3LUq8SKkoehfHyoNi9bhZ5ktC61KEqq
9QziMVklZowr3MbuXK8U7U7uZvmNYj8LioPMfmfndGsAdmTwGDj6m/8szwQp+rzJG7zYfOQ9sonR
Tast/WiwsM26Xg6dhHw/kDNW8XaXgmb+xf9pMlCNi6QdcariJ1z0+7UmF8FDd5WihuK3+1ofa6rR
ZCRplnXraXXSziBP11T1dnk5lQZYlVnga2hNDRBWmbLkMe+1MrQ+BlHS3bfENRxXPKUSIO9ehvzK
Bmz6AwPXKDHsTUPWRLK1uPxIQAwVYkrzuSI890jZlObOd7mpaiFFByu2vdUTwxB3hE1vfC0FmZT1
EcslASjP11917h4eqUfova+4yAJP52wLSVxkjVN2Wr42VUL0yQ24Cq1wlxVAc+oA2WoA+hLNnIst
lwojlc9ZHpN6FmC4xlydhT6eNJAetc5be6h3vhzcawr1TCzMQ5FTVHbOvu0urC1I3Wzl1VGP/du0
XK6IIkNiOjlbsq+KRe+6vxCNnKkFDdMwXPGe1wcOQ2EDJrjElx77+98+E5H2QKFNhDeMy7CXzMWD
f5tbZsZ8FI6ednMFZkjTd+o3AvkVZwjc3hIcDgR7hZzq/FoDDqf/yANoTQ489IAszPPaR9Z044FI
QI12EgWlR8+AegarmQPaRTah2iGeH5NRBAyUwN7Uj+jyDb6MPAgoDhHuTvhfDatjYUtzCZtyzB+D
WcHBwgZ9ASFgfFsvL422R9gWbAXlyfCcPeURfdHq3svIMXEE3NyP1ifeIaoaVYS6t1YM+8D2f8EO
phbBSuU0Im8LuXp71dOXl4B6RWuYCe5RWc1qEhE7Tzm16ncpWNARLQIQPgiB12jokH+v/CLsoLrt
D1ajpJwFO3dmqNXppAVojPssliLFw0dcCrS1lksZXgkgRwoTVPRlpQbkf2BBpArJLyyW6qyjCJsT
3/Dnv/l1pNKyuHtzB/w02RtiAVAk8VQV8fEUzgjikRim43hPTRDg8MoHFSnFy0Z1eBsxBscAW1no
Q5Z4kyAd1ImB5PWPdDoPf+qoGbzxUyF7j5HzjmuErntwwuBjR7M9UtUsjaZPlsy4DKH/S3rhE8VH
gJWmeQ4Z0NJuuvPFEgiYlif/y74SxMSqmlRVzfRjhr1MwKm8f0NOb82E/sfe05ExsFydpkxEizLi
9UV9y5O8+NclI9Kv0rDNfDLYsU4lxKatZCMLWPbRdCi7BQJIubeheRg39bhNCQ1msUPa3YN5D1jY
IzlWicdRZnDcb7EjmFpPufTAO8bRidEK6DjpTe3bFCU+9Qh9wRys+NaL0tqutMbR/Yt1ZM5PVoeF
yy3YKkI/zc+i15UM59FiKV26PQODQEZvvC5oBjc+9oiTS1SQ5sE0I6QvuLzo3zodyKi3WTLFdsAv
RKcRknWCSDbqF6PlYHvR+JdyhVXoDa7RXOgWk8gjw6CihKUcXyEkX172wsIHrscdHbo59Sak+tGZ
d83BXf1ddO1rrliwjNYc6IitiGEGovb1YT9DpZRq4wHfWdm+ZbAOXH+M0v8vSOwqf41IKVgYYhRR
CgB8Lp4+mBQQLo1VsMBwyUARpsGd2ba91EHTbnpJ4VWbVxwMFAsX9XEbFOv7flsSyXA8+QdxpJMF
NR9PbXj5cdP+xYbmgAg5ZQRORh057SGX0TngBTJGvJRc0ZQgInSXY/tC5nwJ2kLaSuKsUJFqNZOz
9oM7pccwwmVdsSrJPCBpkFC6rqiFJ77lMwIHSRFvJyXPIbhbBf+hrvpu0yrodzPEidxff9M4ZfMQ
d/lm8epQIxyxI/QECf5FHseMmpfwqo/yivL51ckuRg189GMJntqgQCiQH2XakESLcCx13kOhQsKs
JnHlLTbncOVPR6cMwTDXtsn6Np75C8PKSEyPttZSHSAmuCIHMO9okqpfXl3b9gzzpHeE1+sNo/pl
s+R+/SJgQ04SW1tZJU3MHS8uGlRji0SgMOSXh89gt1ENO0KBMYNJqduxostdA49sjFv2ABDN6Kvf
NQ80P4fw32oeZ71FBVsB2GR3pKbJBkbZaTfsSiHi/6B+0r58e/2sQHMae3L497Zxv7cJ+XUyO3C+
F0XIlyJo0yPcr8JQWLzoPyqlCwfgetSbWSIbYuyp5Xher6AYayOaDulJ91RaVYOJjdtt8PlzvMKW
6rtEBctp4UJ+lEhe25gdTFwID/e1Kze4fM7DWFoCsWkfXiCW19TgKkKycDeu9BxuEO9XkuXMvU65
Dmf1QysNPqOfj0/1u07CJmZ6vIGkYO+oGEvjCDcKmXNI/RSt9x84HfLm9MqAZe7P/cZLPdAyKAE6
NmbZavYIADkcpRhixGUjATzASOF3U1/ffpGDdGuxU0LYZuvdYl1vojfux6b/otm2fuagm2+r609S
eRPECeuPcSZ3/O0+Auvtwh3v7TdUdoOA1c4Il9DetamTWIph7qDapr0UjRPmKdPQjFw3q+ELdq8X
jq6ZGvgy1fDNdwglbdTZC6ZsTeJjxeWaP9c1M4eJ3ZI7BuO80GIP2TSAyNx5KPSBjoHOous0YxDS
fpUU9JmK4ahsuAVr5Zv9R16/INV5YLiEVwp0HAZZ7OB7Wqe+U1+yOjAdYyMzydORM6Z5R0kHjnOs
9549q8IieOXN3qGE7EYh8ikNuufAH3U7QmiNGmr4qWIz2QNfv/xeIW1fNfd0BnQzIESGw38HMRuZ
BgCMvZrD6nrpJYIBOovkHRr8DfU2AP6bASV36jo1z1wxxBMH1DxlK0ezmGEGNrHBcDebAlvsDNHh
2+yoNlq5C1AwGh8Y649BnZviMN+2ueuRNB+WZvT9fF5ueigi/9lWU6M+aa+yZyQwk1qriySoSXl/
M9L5kZ3yihuKH1sM8o8089kg+Q5lXYpSKoskV7oLDInOjaQ4Heu3XQ7bW3VemIc8owm5asxdbYJX
gr8/IldyE69rNytfHFGf9kvcCPBzIv5oL5l5MRD3J8IuHHTroqgotYQ6peo+UV1Kd3gq0mSYThrw
KndDYYwHclCwKFsQJ/FE6kDinkOG8WCBWSFnIJRW9M2JFCqx6DcwV+tQV30PtmjtjKMfVDY/UbbD
MpKEPoB8rVjKg+kNs4teG3IztNskX4c01wgqG6b5HDPSB+A2AAJp43/brzIknFkBivq+WHTEwAOL
XI93CI02GyQjJ2J8EVCgDCD4+A4aNjui54J0LeU2T4R3wcmqtCpsJRLwJwjZfh3MB+U6MBv6jlcI
m8ZfT1z6BzJPc5ZfSmTApdVf1ZnYqm46DTOZZZPxcMxqpE547lrgYZZiVuPruARwCNVGaF7kSjqi
/bppIV2yoO5nGH7c830Ao5gbslTWKxEjRUB0KgbfXqFD2wVVWi0NyQXZKm8GqvuyM+DX9DGLsobm
Fg6RKnGbVbJqpGnbdAgttgNEgjxy9eND0Oeeo8WcwTB3G1KxgI5uFrlGwJSl7wruH+vmhHdFs3R9
khDGaTpBzV90rutuwVARpstiTzSWrugpjLxW5hgZMFlGJQVw+e1pfZmTW7arsh806lp6FSQ0zTYy
4cAeE0fiw58Voc0JmC68swKSr9PeL86RHmo0fKRr/YcOJiyqm3oTRy8irWZy7V3SLEqpKExTcP+U
1/KTZAV5S6mSr234P518ZxS9/H32kRJyWFupFvUzASzOQCTPMy9zdViMwX0IaFwgwmLDXRijgYlb
DyKbWo7wiwvV2RCs2IYA7AAinDgjiJQx1qO9vFidc84tJRU5S2kCcQQw98dzFGUpu5IOsYUx6TMt
UVZgjvPF0J6/85uP7GnWEqbrpz+Z/5pzN5F57ozeO4N4nAkAmOhrcSiUc9n1J0zl88gLcP09CtOp
bGUaGjgKG41Makrs/nnP4q3xyhDLdsqF4aNIa9Hg/4kSJrqWRqNADTjUUwJcDeL+wqdI1Vtv9Swz
zKqckXWqhF9jiFHrGta9OGQ3csajQ3jv/AGtZeEgrZnHVJxnbw7hPrkj/XeXpBU8ShoTScsluLTI
+nQDdU2HR++vOIOyOLBsZZDYqqEaBAhyGO3BhRFD5gtFlsnGFpkch80VO3XyWkeoMT0Nem/Kou3a
qgM9aFamVey5EEaLCcjZGrRusHpQzTysNPj4gtMtwR/yYn77ZARqyPVqsOsb1AAVSlZxxq18pMbx
2NHfDTQHWrlWNQLDgjH3ZdezSrWdKiBEMPFGthD82ZVC+1GxpV06rX9dHwA/tTc0ugE5uv74HTcm
lw+h18nWrfbjljzMBP+SHaobo2B+lRhHj0ka5TIrCujpLcIMqm8BTDYnfW5ntudaH0miCPwHYW43
RPQ1XGliN7akoaw2STqgm3aBoy8wVMwbrUP8vKkdICTDymYoqxCrG03/pHV3BkEos1TElqhOAoa6
vyCknrJPlG6RUU1g8ogvheSgnNtfrTQVkW7ZccBXgHLS1wba706wvuoOzV44ypQ86f9vDRNwogHg
YbCgkHUxY6E6Jp7599T1g06/C1R/jJ7fs4NLP11Mji6HWw5tzhzs5izx+ZeRTcYNUDsrTMo2GrEe
Xl+6jUYqJZRQ5X88XpdMxJlNWQhWfs5RMIs84UO3Kd36HJguZzQTchv2uEbugrzaAgZlWkaQhMJ5
/LgXhKIrX8iCzOdU/7ll0NR3PxgQ17UM49NSXUn7v0z+YQeyBk4RnHy420XHwb8LinLOg7GLPHRv
K5bzdTWzzle/BBsvkVMZ7BJk4YLkDDhfD5uBsrN21ELxd9LtOzUP8K5dRUWeOpH5FHLnnXCn4JNm
5BzMClA5VGasC6K7vfCMTtJNO6Lr39MIIOdCA/WfHAyRHCWDhItCdew1S6u7f0NdxctCNzI71C8z
WB/GZWVCbRXftgfNyaVlR+VnRMp3SC7xNG6cYHvq2N4EUS+cipVQHR8+d8CVy7K09TPs5KitugIP
Gp1uv04NWMewcju1UbCvCF7MvjiSbuV8xu0RCEETq+RgP878g9n+KlEmS4dLzA4WDLIj43CRcDQw
952F0ret7Oa1/Pda1pXspcoPyLLCfzvUTv9pjlXf9diFTAKOUSOZ6m5d3RQGKFN/IVAFTjb3b3aC
06fmlHMvL/TrMDsVZ6bIMy0Z/VgX3sb74A7Kdo7yq2g50iuQSE55YiEFprz+6lIHZJogd6iyeMDW
pJx9NKLXW1kiqDpP1QAoGRrtnVh0IKak/7jEjXo6Fab/V85ZWuvVnqP54fLSRhFWrWHwj7le5r6E
Q9DJOaqn2slotoNcG2VCFJVDvsxCEjjT+vWGWQ5INLWkN4Mm4eXKDRXn0Y7DzW//7PjPg5o58vwW
4Zk56Eo3ucrUTLhTfngKkfoUHQdqMPDMNiBdBSt6oBoxUKlLzaON9X3v6LSlMlRfwPQtskjxLqHn
diYu+vO5UqUvJPFE96j4JGGz9iHFjotVpU+kofNXuV6By6jV6hCTOxM6uF43pmYrPFRfNcrZE6L+
Agni5sii0eSeK27FeRNUWkAnMl/4TN75p76kw5lTEXfX07UfiNW3rab0FyLdcBHzQ7DATcMhA3bH
po92lw8Uv/mOqOGBUad0QMI02rN1md2Kf+47h1HAPFnLx3/roQcW0pLZ1ipeVEkJI25y7X8FhlTh
yOSDXVjsFQ0rrN0oTNK4OKCHqmWGYGpopiV6DgiyGNsnHUtTXVQEP9cZypYs0tY4YHNJX3ZRGaGG
ufxCP/YSBigX+d+a4IG8lggSimVl2kqlR0TeDOrioeG468FRj9yhovIrCyTeknRj6gKMrw4cyXJj
ZIIpMUic7sh5lRwHPHan2cZ6JF0UnlY9tbjtTTA97TxaFjtAecMz8LV01xfPra0oyEJnH/4hSlt9
e3YTqqVD5vNPikztWmQCq7UDlybVv9CdOJ6yLPGTW4KDZoYt0o5CxgFktOvgQLR06AvhkZ0adO0C
543v5tZjvd4vuVnlX3F1Zz7yBAZe0Flvio8REEwEVG8b2Vdk97/lmXgxl0MbOLe06xy/Df5vsaH0
nYUqVjiDCdCgtNMDblX5cxbvA4Q1LDWkrDWDYk0E9qt76xqisBxKpAz+J1/Al1H3pkeafGq7wc/n
z04B8aCyqNTtF6bVDDFiKuxHHzbsrBbM3HipUCv3frYMgINVqUC2ZuC8kkVe7/I0a45CwVbA26YZ
VRH4+fVHPKWqjcNJzavvGuGArF6z4BrL00S0ppp6vVBHVM34NUgqdCtb2a9wdRlANyE/ipEE4iQy
REnB62Lq7nP8Nez05cRnCOdKXOTjyaRRESyYgXQ5eGJwtUVE1/fEy1yRa4TboFg4sSNAz29co/cG
TGsJGbQsgwcn1+tXibyFsVhmNr+HO3BLtXcV725Xgb9cJ/IkoGYMke9cxj+pqfIpNMOyC1uDwggb
YlFNo7Uzvgof3D3nK111otnZ/fPxlBwfQH2EEFmlZid9Nl79KGbMyOVHJKhNUiZGS9Ib3EgVa9+Z
vULQWKY373VoOD2VksxQ4rEFQy0ThnSHmy0Y3gl0aUpcrvYnwGcrjcDGG1/Z3DMfUOCyAErJHYFe
FSsBtoWy6ldhqPNeJHXDVKkWcLdPSi/LJ33tJT5bUN0Ovd/ICiba9kYGsR5RPamCXX327i5nMqXy
jUh+POTitP7cBTgAe5tRbrg5joLCrTBG3VSUST3FUYtqjDgTMK1sefmy3A+us7zI514obhWQKPdH
BGghyJjS58oP8PIE9loR8kzSQTuX0bHBmTX7aKTzNUhyE2xD3kzODbEZuM4rWwY5uL0bu9sFt2NK
Zyohe3YOV/BDC23+hNCSTrSx2VRjVx00Sf3M0f0ZMdU2T0wOIEZ3ibv8YZ8WkYkRsFcnFaugxn0B
yNRuBUg/iHW90SKdQkTbl6dn5DuIrBocsZJB/6INo1iH+GzhSvGqIss4mYMxPlL1DlVpC9OAYQyx
ABBGcg8J3EVUTa4v5r9VnbKb/WW8j07vBKfdazCdPer+RtyFOU/qRgnJccCxZfkrVrFDWCo+IKFp
p1gVc3eErYgTpe2ChRGe0bXKW9JCmVOYndMnHlNo/w0c5UWXAVISdzv6Kx3hb+JgaOwp8e350b+Y
DvwGHap4QGYhqbsqboy2d0FLJBvf/9hKMgUya3Na/WT6b0I1/a001rNfovjsT9M3IpnA+jv45ijb
FUGXkdmrMOQtS4eFB8FtsLN8NknYYMgDlzUoRv90o3jQqjTVtU9GB8KmXKEZve/1nc9EfdUguV1F
oAHJm/ITx0/I/cAtVwLJpbhhe1vfO/M7cvsmCA6JWrWLuqoh/Wrdi/ln5d59Alpoxy5Nw6UfZTCR
DZmNaFUOLmpHkj8Q37sAuga3L3o9mQZ57ZXULFq5JgtsUeHa2N0IVwZfWBYj73BZ1w2YB0UzyL1E
TrN7rnoRyRMztW/NF4XcMwzsyIGxOyFEAqcDXW/el2jO2XhJPbLOoyQoNKC0jRGegMhc0G8WxjAO
gBU8aVfUUB7KwUu7Q6W1ZBTV/GU6XD5X2k2Oymna5tfSfD+XRKWk83zh5WXupCy8SPfxXPXCUQLd
nYKT2effNuF5lPR7XnOpKKV6NDLFr3JVsMFCtOOy80RYyVM8dCi/EXkrWhQYWqnED3sibWyVzL6W
Sl27jh8vkrHSONVoSgMKemPVsKSwscIxfZYwue0gAReJs5rw6G+x8yQqgJi8bmAg41tlp8T1K065
CTXDptWtiqYaya0kO5QLbxYHvM47ftcpgWSGHo1u1mj320q6Ajg1dyuFiaUjIcwfWY4uqdgJt7WH
VinvO1TS8JvPCH57THfzf6qtZYxtSRQYRe7llS6YADUEng1AgvJWgnmgW+loZE4oDwiG7QS3n2L4
dH4eKS+zpnwzan6z8hb4JYDHSxAbWZSZFw4CEVn259/4GkTfR0YPTWmVsEnARoGYO+248oruZLEC
ONGUAmN/ujMhJ53kMA8v4YLCXPsOI2zdFc9Z6kd0zsjrfhwy1B3SjPo+2hR0TlW71LASD8x91ozU
IEhQywFeYYOKC1nKael3aIfWzgx6He6a/5DBPLQ0uzdxQryvjnICog7A6OMgCGR9yUMdQ+IPwlK8
C2nPTXyX4irDqozHdPKmYjDoOeYD+7a/ueJgMHbFPua+y8LTFpLjEN15i6bJSt13X38BrIrlmlq1
XaxFkPKBlEmC+Jy+I4TUqqDpaol1QdwsY4CUjUXQWxyao8mS1Towz1kmE2Py3tkUT+s75+jZlYrT
SUtBnSpyhm6tV0Yx0zYbzDy1zh0+zJPmM+rYTAhoTe3hNLMshXL0qVhLitwCLdljxeDHF2n5Ze4s
KzEwEoDu6ykINxpqtyo3PYVT1J2+HODdlkca9Y93Oo7p3YYEZXMfd9j1fsFtvPye5Ajqow62GDdz
Igrh0QHsYLqi7YciZkQu0xzqkhNpR/lz9axF8j9rRtP+8PUGF1Mt9cIfZ+UPVRTK7tTfq8WyrFCT
u6i2hB+wPpEFDhwwsJmYOully/uItRHLoyxCDZYfT3O+f44SoHTH07Td+mXtQ/UXqMaO+cH+P9VY
iD64pqAXYSKC2e3V5L80a7+yFnLBysl+GJ6Z+4LUABpahpsY/OlZMNl3Nt101BRTKMJCy5uffgHi
lbdeM2tt83TDAVhqrbhiimZJM4u/Zv5q09cp3Hkkapc4OhKnF3RApD7SMUYOZZ6ggYYmjGkyhVfw
Raed33NJZgr4aKoQxZYoZKTWNx05UxMD/ZaWubZZbzSLsmG2U2Mqdc9Ht8eoc8EQzyS7d0/FtF/j
r4/1HmmIFBTeCt8e2F0jtI1NhC9O+b2cC7gUhCdzp9FJNgcIXBAS0P+NxHA48MLDiqXwoGGYAfRG
isOamNrzCJlhbgc9Fa2fOV1DM5ktgZYwQmK9FRlTO39IAEvLx9ULdBvtAXgpSg3V1kLTBJkGXBA8
/FcKQ7J3Vf6qAK6mGSsrtpeptCFtNwX9PsTsSz0ahg3MbJjJ05FuuJiPCGQynA2FmFwQaapSfSLH
fgbHImK9dEuDIvrn6RpPz0Z+eUWHTYWSHSPSdrqiPmI5RBsKXIPSkLrPkslwNqwy3ZTtsemSDN1a
SPZR4gpskH2dD3jAF7kpHK79slK8Y2rAOuxaI81JnDqdSEqu0Xbg6uddY8s8GpIjKC7j37BBliEG
rcX0iDq5GQJU0Iq4bRTJ16LYIZetW4zrcRwxfTzFbq8A9J6WehVu6yRRA+O+bcCFWLwYrYd+yHVD
8SrsZul0lxFenQlY/eUacrAn56xD97W++MSDNGOGze9Vz3rLyA/VXKFHAWVQWn7844q1j4ubbQbL
zyEFVtSe4hRS4cuWA7TZk+mEpofkg3lEaBmLnSFgDT//ZDOsnts0UnpehuOlXbcQLUkmUPoubW19
ClZbJ8OdHvZaFGGBCdCBvy4bK1LPiUL1vmoy0t0JRTltk2d199bwRhCMCE/32rK4jGNz6JrL6FzS
65NX2cqCS6/u0fwt1Xxmn40PYpds7+kbvC8afQcuoIy0gfMNqE+M7AY7ywd+kIZp9wXF+KOR9L7b
1OXL20fIjozL2tyimAHsC0L5+6vu6zlhFCU5FI1QI9vqtom3Z0+SZTEdtO3X+BqtyN7E0Z5HfhZY
uMab22+c68ehPxB6gbI9bG2c6LRtXSig5zOzcxEwysQwueIwZWzOpLE6aurNTtLmhnRd0WFPm3fw
6Q/NT9/ke9buZe/GupXK7Iu5TjZAjZA+xmZwteG+kIMVEpNaxZAfs4T4bmwYLAaAnxIgDQggT/jC
bTYjsiCzpw6XPKPby1Ny67GZVeNKjiA+pGgqgMemdjbSGeiJ2YOCwDAToi/Ldg4RSuW9C+ynPClN
ye/3UJmFG2KiO/ywFqu+seHTAG+ln/lbjm+V7w9pZnGav9zael5uJWdxpvlNRAa6/bu2BjqjfDdG
CrCAVIiyP6ODc7923X5eThuOyn6oZkGrGcTMuPlhf6OWIAkLw2A6onJ8V1qXlI7cXlGjSIrr8yvs
IDB73xVzT65au90EPf82fPuG0oWOWIAvjksHqjJXbAjOpBNcMV0uhHM+c0AiQJV37S+8Z9izbNwF
MgpFsTijHQFcX6eo6HdTIkQSAnRNvXKEGz14lDdu3DAOmxyrXeou0rtJehEDoQ+R2W1WsevLqEkT
joMi5U/ELsUYOIJOH13T3ePTJmFakmaV7eie6ZLzFJ9z20wFPpShKyOwMrNnBA9Bzw9LZVaO1Aoe
ssly+j5fxwunEW7yGzgIF9VbL8XBGUJYT/0vXG/o9E39ChnQD7DiYjmhjhq1Lui2dHFoTWlV2D6k
5CmZ4KZ3sz8Ghmnc7mRjm4S8b9pWt4p5FrEHH5ogOVtt860HT4iV5BTSLPX6mlu2hDV84kDM8NCA
ddTkTpTFS6GkDZJ6Bi+PyqykQ0X+7fEaiD2TWKVHHiTzaOixs/Igu97ZJFTiV/jjopE8XWClhQeR
Pcn1RSbRaqykUpZQ3+5sfR9UP9yrx0WR577lKWfZSrmjOPN+15wCWGH7uZGCg0dVswLjvfjCINUq
v4yDPev5W6F0qcZRgJUABOJ7RPDjhabvd+76Vat1HsOlZeOMuTqa54BOMZ0Yrt5CbJoi0fDQU9fr
HRk1Mt+yqlTEQjIhKN5gVZrJ9tybEpX1BArfTxRQdpJ93TElFe7zyisaM2QN1a2fkulRIvn2+YTB
g69qGL5VM8QOjO8LlZqqFEBoj44kBo6dYA4PxhK36d8Ibud4PQJum7jHN4VqD7bEwxfBFbZQf/sw
2CJDC6G95GZz6dwfp9XqkPHklVk1hkM28MF1HHd+lZtKmbL4P1v0KASTpzcb5Kx7x/P1OY2SaZ0z
iXEfv8NTR+OjNhd85Q5SrwA4FRQD5NDxvPQy3x0L9jw8uMh6OZ/Ty3Wob47GcEiE0ZqnQRX6dPdT
vkOQSzVycAUpmtjGSem1yGZIXQtZEFBaRC36F78rbXGMauXkV+FWJkY7sUn4AcQMDlOn3ARpzFjD
M6hjvggRHeDw8nt7gIOHXLtuNwS5vgc6z4zcSBMU7UWqDdt8Uw0eSy91uLy2mNHTSFTmwJbMvtJn
LeMV/Ame29EeNnID3RzPrDQiljrSYksrVtIQ35BCdMWM6Br5HABzlg+wkSXor8xoCxsDomXvXrVX
wtXqdIIBzFnwTiuRO9J7Ce24b3qnsO8XfTCWTbXc//EOiihZCux0i2dgkl6agv21fIcTXWY2hDb1
7LTT7sFQIzA1bDnf8n5kaPOPWM69ryclnvCBjDwxu6F0zuF0bOmWGRsBRk8pysbCD+Z/aEnrpzXL
R6h1Rr8BFI2yb2x3dksQImYRFiVNe3AmcnAZeWGrjLqyuTzC2llY78NBWl3JBSW2LoipZPau7v+9
YI2+g7OMMKNynuzCRTKbZVtd8mZyj5uo1J5wfu8kqY5ujg9NI51Rgx2gv55dSFPS4Q/rN2D5akto
S4+5Ore7NA17XT5k9S0A/PLrS6fpGSLw42GhaEAPBMlr9l/8ZezegHwTPuIz+z2zoQkd4sXa/zoZ
h2Udb9y1SAv4H+oQVVoNUq+RolD/JlKOjPU7fSjxZwBwnHKQc4P4v8IzUXmXwg8OkBg0Z+YknkSI
Http+m0FM0sZ56ZlGfMKGcxoOQB/PbF9WCz2cfMWvf4Lxdc5myM5OjKP4n1ycONB9+NUFk6SM+q5
O598UAeH0PiXR72NBFQ9BE6Ys+7FQxequf52nLLjlShcJDNwqOQZY34fVVrcig7cHpAg+sMQk0FZ
rHW75QgMKvtMpn+MLgY30hWU/PP44l9j7VKs2aVlp0OhYu5GrtcSS2F/QL5np9iFUzy2xCXpQcdT
SiT9A/hVOcN0AP24rWllJTL1qu7w+8ArOnGFK1l7XeZt8z0D8oUBP0Y7b1GWvCN9+PS8lB21bO7X
JVSt9TFO+IO1uigTge93i5CG/so9sjN13tt61iwZHJjxtHpKMIzfWD+QYieE61JkjroPLar0kU6j
KTHEr3yKufElTl/iIBb0q/cjpaww1S61mLbTAHNrXuQy60KA17Jpv2miZCcptw+65iy8NtgaymvI
iiLylX5E6zSlTCqeNG6kxEP49co2B+5QvlZKgWeR6psmkg4ATptMNqUYJbo+PgSGrSVI9v+hVsUt
2t6smW4H9a9OfXNR52LU7BCwU+ZahjKQJt0s5d0SXunpi1R5VzaIUbseLZOb05BN5SbS4TJIYtC+
IAJg5YNyRXPX7MasRXJl6P1uMjQ2GllFeOqu1rYpdFe3vDISJ7QwvKc88yMr+MKmaNoEAYbzv0oG
BBAJf3Q/c8YrAVd2p4ZCMTouN5J10IR4Hea2OTIumnnshr/2i23TOIqThW5ALvZn3/FUlAq1B6g4
JTpcZHUMB+PMNpx+A8yZrq0ia/UssucKL0ZAuCYUd0mLxptbKSPiTW5E/l8j8TgZ4F52nC/C2eAJ
F7uuH8mkhBB2mKOHTAT7ktPZtb2l95Jo7GfYLSNJozRwTbS7O/MC6XAEuKVrsoxzYp+GrCq+iaaL
aqBM4+u7HZ+JTbB0ns0yV1ZTvCvn8XYHs/J/a2L/2jNou0MmAR/7T/kIITFm1JZS2pM4mSfVPXR6
vWk3QfF4EbR8Yvh3iFcVFTHSikMLxcLtNJJBqNSsECV+IksumaEocac5qsB8vWtjoLdtGqVmFOnN
Gma1aa3rfvZLGdQUE3KFxbfVSabF9Dnl2KUsnqzyKtA9mCXN2c2JQPiRtcyeUVnrynIq71FY1Yug
l2r0+hgTMvaOYPWW13iFQ4Vc15NQ+RpFjiAimuXROk2eI4wm7ML+tKPVKi+OK6emya17WIdbANZN
eVIWbhTvsJbiYloVwoiIAEcTFEg8zSvDKk0z5bSr2svbq9Otk/o5uB2jKEtU8Ld3tnYU5qkM2okt
yM1UqMkp/mkiKUeYGYuH/c8eu8M78SWOPb9uBV2anq1S3PdLw5WRK+VQpTkiKVISs2UFYtW25NNx
1wEjyiJLJ6WYCMzMUUYJF1lgd+v5kTfmrPM7QS7QDMKnOUDTuJuLygauSTm/inSLoCyYSX9QKaJ/
ETzE9m1+osvDpcwyTvVVJJTbFGUeFSSKd9zNep+cfwJcsr9F5QHgX4VM4r2cPCx7tXdt8oeyDlhZ
1VB4PzfhMM27ukuFy+7w8wU7gkHIjzakEg/X+QoDN/x9zu1Od1SMhUPIOpXgFb9WKZwFAzAzdh84
3sR3udSuygsN3w0IYaDMMvWseO2ViEIhpTdYF7+BkCuSbZYzcXeo7jXlNdGK1MYKZ6oXeC+0qcJI
UnMf6cm4qaQT9PSzQAiREvmwAqEsPkys9/XqBd+oku5pOVouoV7tKHAE0cjSnQN/PJwIUtJZ5yOU
DFHA+TseB/tj89hXgxAzF0kzelV/KdAtpxsPEBsAlN7CnzG8v68wWquzSs2pTF75dsOPJ2+vB/UX
nXMZ++JPiwtkk4I+LdBRlJS/QzzuEBA1rC46PGxA/f8wTZC/TxidW3cJTAU+6QD7q3iHNWgblh2Q
PAIMmuCn3m/HAuL6jlXZCODfJV4g10C7xUOFOqTOPJ1kkYVeNokPqZ0Ck1N7KoQ9JjHU8uDOi/8A
Jv+4P08OlEBmZ9wmzzmm2893wBCX2yNByS904a4oPeua1pMmk/ZvJO0ysyE/0jlWmOVKb+gA4y56
jiwF4afQqOzfbX+X379lL7lcoyKl7IFxAJGn+7yBbIXFvUuJtk0kj55H3ouqLJ6CAnQP8mUoK7iA
9zCfv9we1HG6AsrwKUZ9AcUmG4W455YroHG+zpWfRJANl09sAIOWRGJh4uSPwjPEDiIcyWRrQicl
hS3PCLmbYnh3w0lzHdAZWfV9F9xLVfgbdOeo2q3qtN1HugpixaUd8D0/Ra+M96YEULoAOnYp17oF
VrFeYC/PEGNANr5Nv55w0Bh2EUbdOtKZIV2CwScg2G+Ug24HguCKq7gei49y/AKR2hHGTnOMpdS9
95GJEOVUsus0r7GBDlfSnfKav8+/jxhQciVPMy+U96lK12kbFTEkvYmFC8SrreIhCSfGi/XwpaIF
/ODJwJ/dJ65SEGVxLbulWhUG5PZ5SvZWPIZZz+Tbj8B2gc+0OfmBq8sHTADH8IanqUGUJ3JOJWPL
1Z9umASJl7scTmfl/rf+YapMxuJaFz5bLcXsUFGxSm0U6nIlHxJVazMCad82MXqKgh7KiW7aEBv/
qTkVCqvAjULFgXRovLMmMfZ4U0KpYQvVjfWfe2kG4+MDgCzmBIrZrayUEmYD1SAf5VVvnS+vEpNn
QdChmPFGzP+vA1KtomkAEzfB4F4HBrYdBUOwBH3mp9fWprAxAcG+v9T1OKXzxoa2LiFxLB8cSyr+
3iPj2DlHXbMPQDFm5tFdTRCEF126nMS/O1q+TNZjwefLXaKa3l95bnrcoMbX8mmHf/dzB/p4r75d
nKz8juTmohwaP1CPKjmhTrEW05MtTWNlLNG0mjchgGsGbVbbg3j4fljiUfo4rQiUsH2Xkc+XSbRu
yJGQH5soKfeSJeMgmGK6FXQoHGSR1AI+R+5KGtLIesPXpEIEsvbFGwORRtCKOPcAiAs7GMmhFivG
b+Nafvm37PyTmFWGMePQNa9VBkzOc5LGyYMjsg40Docjo181L7sFN+MjZ6b6CCBPPbcSbYjruD4Q
JJFOgM6AnzDPJlQnjJ5JuwQlZS5x2bkJ2QEYzbhgI/0m3F9A/AOuD54tPC6kxaYduxdzLeTYNxPT
HyTspKUTg/FzdlnXCA8/l56q9jXnGHejkAh8XJ84wdU1NZ2Y1e8VEo+oMlAvAYIC5KzahX1nqXPJ
elGOVxrNMWIkv2i19EJKhB5Wu2disypDBpdQXvW7d0Is/VmfDKwDmIsuhei3iZXe1VSsEfz77t2H
c++Qdo2ugvZJPGjAYN/PB9n8dGIfqskg1yVYFMFyt8ozMtc2tS/HBPbYRuRnPWhD8rLb8f0AtLCc
G7C+30iVH0K508YW2cocbWHKpxrrh2XWDUUhjJSGBoBMz20CpHUNW3zbXF1W9fC6rcgUDPBx1LHz
6GSZISSIci92do+fkHEbTY9Hlk9cOH++D4ZNDaA4yllzM9fBcNywFzItdrUH4HWOUbB7W/gguw5a
zRZhB/6fY2oxXUh8jy19dgICsRzJKK2aHBs/k3gxsoVPqiQOmwhEplVYHhfwwxU8FEuryP5nJE1F
gXe51wzWilPX5nQ4b2sqj7CvcuhrZfDIaBSZc+EqGn6WUIP69OULmA6SJg4zxuV0mxWj+sqhoWEM
EGiDOS32MQ6VvU3+RxxH0N7muwkm7UpjXgyaOQH/E6HYdxhs6dXC4oEXNdAnmEme+QKrTbFMrLjD
soEz98cBBy+O9TZ6+JCiPCPDCeXNY8BgUJZj+GR5diruXRmhNhVtKPD+pzJaM9LiMo4ZJSvTbTLE
/UOdjJR83c41EVZpWFw3eqGkbWfJSE/WMAWKp4EkFiWZYhFnn4/zsp34yvvWlEiSyvhsgAuh2pWC
dWV4xHaUYrGLT2u1Yf4hAlNVw/QZzsT4xbQXi08TsJU7bpUyzii8Yn19aJm8yKHE6MOnj4gnW0LM
Xg4wIU9AJ8By9iufHS1JAHBXVCdNuKapzPLvZgUG5rz8yB/GnHtPsOGCWwhUf2IcaZrh0uw8HSBt
6Djw+StB7O9io5ZjcQ7VosLXOF4pD2hiXqzTCZ341ulsjiIAWzxA6h4Ec75JPIpk6Q/b0nEb34gw
GpXLFjsLRvg7Nxk5Su/3n4ykfbGwMHooWfjvtwFeP9uWgqNg3j9Uf9/IczPJXoNI/rinNDoPs26q
KUPXv5juLSgt26dfrLdpIAIglWTJ2Hs8aeOvjj2xyeFiXgGedyIqhsD7JH0deTHQ7j5ds3vWjfnr
zEGHFXWEa5gpqn9DMBB1RgsbF5J5LvH/6D8eMm9K+NbPTu8HNWo1rZcp5BjWxiPBLRVDy0JY7BLt
GmtHk0qJDqbRykrpi8zNNC/hudxht1ur+Zp9MvjsIT/jlRUMtNVxjUQCQBIKaEHXCZJlcMzHbJwV
R+m1ZylWNpw9q549WQ0DN/0YX72B9M0v9oJF1Ey842cO+mkFC3TPry5qHM9IMB8Nfiv3uVefphTX
4Z2cAAsbGjHiXvUg15S2GZ2QlHkhu6daG5J97JeQ19jyqAOI+gI4hwrbX+ZNUKH0IA2zyNg9RSYu
/i+pv8hVWMjVSPJXCmpJHe/KKYlr3bjDT5qlkqsRsZ09xCQS+dEGoH3l2x+grJVn1524Ch+dtGvU
1DsDLd73gefzXxuXHgrwY7/UCGCLRMzRYpygG1QF4oO7I+xfSZzCyNLKYTBeRyKGvypt4s2SkzE3
2QaUpgZ05EAve32U6eLGcNaUghC5fgmWKgwn1a1waZHz/xNUiVNOL1epG9QsVcq4OJOF31xGaDyG
eypLIFfdJwEOeZTuSxN0XsKKDgW2Gx3YsS1nFEqNX4VPqPI81JGFWgFRPJfejVvTsl1h/NWvjLtF
3qWedoWVkiLa77mXEx7YIks22nCSRZM1yCq8S2S0uom0cy+2/g6AZJuRydG0nDOS8ukd8UCLWfza
+imwKQleqYUiYK/OkgHjATPOhsXFmr9tf70YDEC8SfRJW0OqO2Ny55hAQC6G8ovscfsTx1XcMy2K
5vWh+XPI+ZFE+j6GC8/MocP01ljk/iVyp0hA7GXFbOx5iJFcRctv6StCHl052KDjPg+sQZ7HdKEw
+B0JhNFaJn8zXya9Ke8DS9ipIaR3jvNNi0l55hRULPfHnGXdqAf8zLNcSjq8rlxKkFyvhA090IJp
7EZc2ncjHcTjlVeD6X+YlT+VI2rbFPGfmIm+JMh0tyuuv7UPRXg0RcgWIG+dCn+k64ZqyLIUNY8s
jYriIzFXsJgFoxmbXTIKrjz62s+7WdI4QeJHTKH+blmKUsxYWe2AqYsd/5zdT+Xrnl8YVoUeyedn
HUL23rLfxj9rODGy61Zgfo7CYEzG0wKLqdZ/XLkAds90yRPP95hp8SNDh0+a1RudBO3NexfKLHKE
/6qtcM3u+h70tIQcb8dL2Nr8ZQsGeIHp/SO1qFLjbaK3RSIVwfZsU5Z/YRm7pAAtCvZA+yyvMvUd
v+iuTne7DTc6eGW0KnVvNl7azGXg1lYqF+ie4JkoTz/a6Zb5vrKeB2pZll7pGmppezI8pc8mfcwK
GcdpSZvSViwYhRB8eSQEQVyFt4sMP0qu2Lx32PwyYuRc2y9aPmG8k11T1wJAFlXY3Fqb9CguITMQ
giNwZLANK/KaEiBcTgObWFOiCUFSqcoUqapaAPxzvaSGQ4PxtTkwLGKoU8f0K8M5P4eAasHhMbws
hCExWhoR0M2XOluuSJ3rUZNIlkngoXaDKmUzaMt6Y3cTYfAq9pMbY+7S/Dem7agR097nQKzF58ZJ
2EZ6jhsG1mcF6NXgFRVLD4LjLhsYqi2GWDvWLQbv7h9EBWx0PGeI6u+SLHVgcDMzalBRot8hHtF/
ZKS3QOjtCzkaX+bnKqa14IBKlwmdqV3lJFwYd90/UpK7Dtqpo6Lcu+IdUSaq5ubeDqBjOsrCDVY0
btU1IlCN8zPFSISvZrEH04lh0Ic0STao7K2iT21dl3fjK7ipTAgh9ILlHgYYMSlLrNaHIhNPRNgy
yto1T9861jCMBDbL/cdg4Nft1z5jRA0wkUeUgAgCdREReham/dsrnEyiODjAGnc73gJUlD1SmTIB
7zcay8vjIkNoqNc+K5OVfhD8MqSWeM9FJ3x2FTgdku1YyjVEvc5A6ytc4v1hsIp45fhy8q/1TJfh
wAvOAdaFDWS196qXtixXSDJShkZtzGb0YQfz0viAIztJ+GLau6EleeGHyXCKRrNZyDmllYimjSIe
FRIp955QKmeZohBirC7CAQQ3+dsPGJxc4kdCCET3561UjOqo01WScBv53FGFF6RUslDVZP1uFubP
H7l2Ij0DqUBb3GPW4C1HSzdgJ5qUcLpIfgRWvDYwN4yNdy24j2+ondd5Us+qfry6Mrh25AOPMKb4
vLhuI8UWtQC9r2KSvM+jlD4OvPoWK/5P5c0K7XbYjGKzDhY5cluRJ1VK4aC1ZPEN8zXoC0tRueHH
tTGJmHyZ0kJzSHIf8obXU/Xuq5aUvYK6uOaQIO6VuNlnF/4vClmv26+0y/GH5+jUf+2nprxviB48
WU4rPu8BxINmlOsl7FebQvJc09gcf7RqNgHbkW00R3xVKBRjLS62HWhD/lExpxilVVo35k3DzX4O
ARwNFm55rv21EWGws/tcMMythIdb6WbNkDkgGNYyTlihFQbCP7fcyqqi+ZCH/tF91im/neoTV2ge
i1omXb6+USzWc4gsXbDq1xayG4PznQxUfivZrmJW55aJIO96922norIYjsHs+BU1Pkm/elDixmle
Ehx97Upu1cXFlLbI0aaZYiRjVma+sf4GYxlSQciOvXPYU/6IClLgX8KeBgHb2qZ08QdOvLqMl/4k
anTYJLbidDe/5xYDzVQf1xD6ZQFqHHcVBSYMzTAHqEOuWGOyeM/k7Z9lBzDWwaCe7JVskARPrZby
dOS/2C9OO8D0CQZjrbPiLG+7RTRsldId/onE3B9gwHjBvlzYNh9dwj2mjX0M7GKkaQNrWHvJvDaG
76uGUte8keHfInDsUe41dGexGMBS8pbCu2lhdyDn5X4j9/wlWAqa2Q7uYklvq2tSlh9gUc8MxG+l
twoftYJAhp+VdmXtGL9Sl9QSeBYwaLVdjoGkigSXMEly2D1aa8cvYi9ATpuHT2kHCvxsODa0pQ3o
38z7e+ZA2uqDaDSwlUkstkSqemIQ7eNpCRk6Sb+sTaLiKFQwMUnIJ7vNLBwcKjySpZrh7r17EbZA
jqYaWeP+JZgJ8WnGQs/raK03weP7AQzIb0rFPhPSPRyIKJ4uTwuebo78Rt4WcEk3O7cqZgIynauH
ddnNkw8YFqcLa22pYWFR7dEH8OZFlJEWv6gKCVnJcerajT93Y/psLLI8s1hGEBL1d3a9DFhEt6mW
Rq38n5yfUN/ngtmRXLL1Hn9c6UfrEnUELtSandRFzGPV6W1D2ty96/dXBS7TefuH35Nyl1/yoFYe
rqrf1ud1g4OMrfSliM5oKSYrYXmUL5zq3T8iaJGEJhdfBiLPu0zKnN2Dd0fl97WesAUa/5Lps9Kk
h8Inv/DnR4+vRzgF5M3hmiiEjyw7JcO7X4BkVt+Y7wVhgqREO6dL5h3cEiR6zeWGF6AhlyAzHuFq
pPeULgyHTc/5zZZtMOxanh4/hvokHMiqh1u0NvvAib9JcO7BICjRCB1JwZBlFeMZqgoHRnfJZJee
2b+hdjRJiRbR/Pzg2dCifTVKXxdpFoFt5PBwUhkrsVqueEtJE8oriD6TTqUBfwZgQsGMOQZ8zZlj
ZiMKeClTKcZ62XmEfYYD8IL3gn7BdcaPJbrg1ZoHtXpvhMCKZBG5U+eG31m0bkCEGQhMtWoFWaSP
/zyyf24RFr2TeCBVIOb4STpn9j5CYpw181UdlQHIphVikZW9qE2QjO80FsyGmwJGNIKC14+bT+7O
A343oopD2kwTRIYWIUFb9CxsfhwtTrsFawt6Ow1HXNJH6NfqVezZokSIpCSsxASe5WRVA4vjNmxD
sD5sCbF1q7c3HvW9HfY9Igl/IqWhXiRrvAawXfPg1nEm1hwU8BpF6w8p6g6eGVaJHtIum7mJ5JnF
jJv86mxZJWRR/XJ6O/eA0w8ui5OjsrdX49H4564KVPEnziX0KU4hXCwqIMky/0FhGFME6yfCu1PV
wTCX/yK5meoa10FAaQn9b53xovItrZ18kdTtr9ERDGkZvjU80aJONr3ic1Ept2Bz35hkr9DtOClz
CqWfi2kDqppFsbeMpRkPbJZVLLwAqb9SD8ekOrB7/FiJngh+MfyMhqn3nOhit/k8rPKPZk2a+be0
ZzXPebIlOBlFnG87Xv+SqyH8aFBtoN4eU911cb/epnxoSe6nf4SyrZji+DT8eEWic0YsgghTdHGy
Dl9HverNlb95vxmLArqDB6lsWOhIcDeIAGT0vt7fu7XxKlHCDjK4lB31CbCGQchxyGmQAZ4DsZo2
isGBXYs7AGcJwVsjulYqhvLr8Ads2xn0zCSYDo+BGExquB64rUpalkk3d0rlrbOj6p3dsLoqAe9p
Df3849eKrW+mcKVOVuyCcxRUMG2J3MtfTHkrMmNagfhXvaJTWkDJtL3bFN6/Mke702DSfJVldRYA
Qz0WQ++yQssalVTL770U05pjQ0SGlRY4JknUVDw5rZWaT9O4l6c8lbtSYsNOCSyk/uzQswejrmpV
xrbZdylu61gXdDU4FDBRUAwOBFNK/6G0rBEmYWiDm14+btijimPelt2/bUy5CARs0qwfxt+77xTm
zUSEfqSaIkOIGzjGz1mohTn2tG3CigcMZFVB1xGHgNxkt0hDf8ypLSD4jgPxsjBQWqV5MnO43/br
6nVtYBjmPlVrgyNWJ2wEmnPRK6lqGcrZby7jni17c0TNGPkY0cff8CSFXWfs17mhufTGoFEnpJGE
Wa5ZMRkm9QsQ+VPPach72gBsOLVNJ4rX0ztyr9p6w9F/vONLT/uQ56BKwpiEul93ASEtPmY4fI1J
KpWHhzSnT/OnoVhBhsHfyKU1t+nr4TX4QmS7RzhRkULhx25+xE11bqIKq2DFjcpt8FRE6bXCfu47
EtKLJXXnHkw+/iLzpey//JYJwllNEVDHHUlsgT+f5N8J3TERQc1sGTtD6w+xn8X+omlCw2m2vQ/H
ZaFIJTcGhi1CX44N1ZvM+L+T9lkodEJdtrDzLLRN04Kw1vH2hrL7/sPG2bGLM36yxtKEvqljeV1Y
6XpCvENM7aChjEsm4Ot65Tk6l75jZMPRJ3ZukvJSXP0sH5NqH/Jkla0veMPKEDmZrFJElQRNT3K+
guIC6ZyhqoOuxDFbHYw4vpDBSbGD30C+sLfmbdkv2IxfzX7hg5WaiC+42zRUsNwM/nZTIY6rgNTl
OJBWNaTQNPaO9pinK+Z/mwWdQiYB2rFz21MZmAfXFJm9qDCwiOI7xshH7bPd9PATa/hwipcq8LiE
xJdPNmyJM5r8crwHy/XnkgmcVp2Fykh34nQW8Vb92nwHWQCWieaPUbMbXGnhfaMHB62v/NvRK8j3
iZWGc/EwcMLm/oQSXXexKlumgIDy73KGABAVAGxWb/stTSCMRz1BsQ+o9dporins/ZNUY4t/SYLF
VGvhOnDgADzrM2D5ICLSvjwgTBmQ9KJJZ3Qi5SK9KlQDZlqsvF700JkN8I2ZsClhA+M/L/OAXNVW
atRERXgB8OzyO1bQQRstz7qajFPzh8GEoTgMspYxVX86skesKc1N0Pw9nKP+f9HBip9B4SvL8imo
eUt+x0yMHqY4s8xHCnNWrWwsGbxQ+OFeNBzSylsPZJZfbWfGtggoXIPwmNeqXTzfZUiojZsGGIY8
M/fLAHlmIVmpmEzx7rQ/L047crULlbbFyUcHKP3Yk3ts5464iJIPiY9McOo3LpMq5Ws7T6r9Qbds
G3PLnucxJoCYBaGElFHFcC+QsoR1dYvsDj2HkL/uiEeb7I1T+CqC6IHI5GTV0JE7w+HzPngYr2y5
bpy6rGdo4daypRBev29Ry9aklE2p6NmQq0yy3kB3YiP0ynFsRzPrdqnKsjZmnG+uWVOMvoILURn7
iMmtYZtXUap1yxOtLkXyxGjXxM2e/rz5jvqt/0n5Qm7WSJX6h8Wz1GrUdgJOAupkkmKaxkeLMZmu
EY8zaVNyvPX8Q4Mq7qrnnNcq5NsGJT2leKnQZ/7HiqZ1IbgL91lCaFHPMDwgHvJUjmIswsSDlCNR
dYO/ohKnuFSEviy2CZc86cVkGWASshnTPcJNnP3khu7XstfZezhJjZsgeJIQgPjrRrIp09v0GaDO
hbNiLlPyagDWJfRTPkRgV+J/gMC4iaeyFNHZGASSMGnhibiJ2zOQl9yZ839q+z+rOlnRV4j8FaNB
txmOr2yMigENMU9jbKLG4Nzcd/zXd5WNxzBdhl4nqSnw/MhZZ4ly/zYNswoNTPOkOuUU4ttjUpJW
3aSnsSqZnc3zvsixOcIGat1JWnguCJ9nnDYrHb8m5GQWURaRfA6tTh2ufUS2Az1x778WftPj+nI3
suavcnieqdOOVuLAySoiKjhhpzgWal3EjHYXS3AqQVbh6A4wMHdO8kDzSjGkA3Ku61V4JSBMnHhM
fLGU+uJztGSbMY+1MXsCFE/VB76u81Cix0JJA3PoHEleyL+b7a3uwrQIeB1m1cEuqP1ISF1fWc42
W2KH5Kd312fS/azyU+5kfJMjl7fxjInv8Fv8LTDXnVc6M5gKzl9IG4FzbJ/BZzNZ29GHW19hsFUo
jVXF2WUVcfJjBI9ahYC9YToohPJ113vpBFundSnjAtYeHzhBDLCYJj6GR5wovYrgiMq51/WS68aM
io3GhoNjfRb8LSctBArSIaJIwVJPLEAHoeCjoxQGCeEiJUebR+mBPewWq+AaPN87FjJYQUjeMVPH
vgiUY3hmTOvLH963SnFm+U+U9ku1QdhkGwjJ5cIbYZfkVRPbwX+PMdUFS1rmL4JRkMYUcIJYE6s7
FM6bhPIkoNnmXoo5b7CxrvMTbhUJbh6W6er3ks6/r4K+RTq3vMbJ1vrd+0Vqt2h4/rm1Jdg19lSH
gSq3sOm+d8+YLbEZZfRoLE633EKnwM/GgTNu2IvTuRZUgDD6j7ypxZuUXMRjprENCXzGGjZ14+o6
/1R5yq47wk4bftjzyUKldOQdHs9r3WgSCkqPXUiuuS+YjZYmlybTQcYYPuQHaJ1sk2zWftrtn2kI
2l5NtxgGLVohxPJO2YXGE4l6mYRXoVZlGwGuUOeooWArSKoj9Uphl+viHju04ZvlV1ZOh4iK3ek8
DKqRURPtVVoq7jthSIjvXHKG91k2P2fGhHoM/DU6koXYd/rGgwlkoPQSC1sQob39EdWef2oHYJcl
fEvuK/3pxpX79bt7/xT3RzB/nssksUfxqEv0c+PBiU5cLOmDdHNWPiPvkvgCeLqJsa2Xs5FFxiDQ
99fxhGrhuKM0vGFRGOQJHVy4r7AejfeBtceNRrg2w/zlaZCXRMx9eWSfJk4IkaHvGFyH1t0J3J5r
x9pnkQzpNpB1m9+m4unKuMJ74GXc5plEyt2tS2+sRqsXL9Y1L5EDzhtN4jopvsLhdOhwo5qpOiEk
PJ3UMO4BjP+s7mRx9xQB0WcqlLErffKCrhqrboCEIMWbargeNNlOIvc002MeB4KcEA2Gyp62u3PQ
xA5uNuH1K6KZWtSPzJ42VnDc/gWQDHPfQ1ouwqIMbczN/twHF7hZTfryObeIrHM9OixE8JxX6PMV
alGfFoAil9t2mgjCa5ktHmWReiSOpiQwov1vn0Vt0yKGTGWb+3+bnUfpT7sKOntagdIm8rJ9OhmI
v6B5JNEkAVm+QKJ8SMjqLbw9ZFHPJxsXbDCNt4TafsqluUX4eby06i/FG/3tEGrAIXatpz1dLTjs
dt3fEpoaXIluX2rW0kLJp9QFDIN3N1uIUFh2B/uiV8RBVPSTvbrdQ87f1hMXwlO3CEz9Eq6wYXGm
qOrgH/DW/9bTahiLDJET2s/C6FmkBBQJQc3e1ZtnU6xzb2vSISsKKUTTddZf95l2J2ZYn2c6aMgh
wOyTy4mq2iyuTsRZozoMPIHZAyvHO3XTgrE779UXV+MmeWQDdkLcc+IE8its11tRPtYxIwTikaMT
9A+cuNFTOGrTGNz6QfNAcwVhU1tuzeQr8wDmhHSGbyp37OTFk7JHvRrQR3UGYln/33Ym/4AjWIwW
4/qP5y+zvtVnJYQVed7LGCNdz35XD1r/mVve3c3hAwt18XKX6v2/YklHcACUKLapT5sR82ctEsGh
2jdzoyOfhk5Ak3LniAKgKC7zR/wKTY/AahFWV9IU3TAEJFc9kDozjDD0S6Va63W1S4yz2Z7UK3Ef
yTW1ZBdTvh998IvkAuMeFXFmbogSsvPr16moW7rUDHmWsq/IXBVilvjMlCiZRkk9hSgGjb6cKWMu
F8BRlg1it5WV78s6KAX3n7uCypM4jJjqj5hQ5PTfPGqOCXhYRD5kZK2oOX1e9b/2hzXfK+oIHr0v
pWTGtl616yqBYIDJsmHRKT64X8YQ2veSPqZay8/GiZ1IgYCPwCWdZa2nO0RVwY81zkOWJdfQfd5N
t57r6uxSjtyP9Osddxw+4MRZKaR3jBKgpBVe5P5gyVy8RIosRug6CTcEXkqVbIsPi3/2yy7AcsEN
7Vt1fqXRu2eq4UkX8EnUNYIgRdWmAZ5C5iUD4Ix3hKoqg15Hqi+1M9GNtjI48JOabtsE5noQznqR
sJKiSI1/DiL8AdcYr+Yrs5pnwHUN0+tZpBt/Gl5THk6KC45czRkUuGrObY4Upiw5s6JHSrBqV2dG
lru8zhxZZf3iGEEFcQrWnlqTTQC3Kf8vq1c3XiRne2Vjbj5gQ581iY/UxVsjG8Mc9hOQNHaRa0KP
MPIEealoxlZ62Qyw+Za6R9YRImtkEK/yiBhgpOfaGQUqb0pmRFOykFsbwi1HuZJVeKThgNYdiKQO
arOnlYwtdTOmSHvoCAnc6aKhdsxPp7BNJVfOUrQOg5eJpt12suYEipKkpBlsII246tGfhknzQMd7
LdCfAMm6C8tDMEl4GUAz93gChJjMtMxABZ6FbdY+qbjsdJkvwoq5aH9BKPEvScTgjYcJXmlzTAjp
JLIk6UdR1wSowiSTV390qz3CevCOxC0dIjrbxlNWtejYCf8xcizYgvvCOcMDvPewbpZ9DCFF0XVu
S9SHfL1IpkjZuIQSXPla6sd9Lm8bi7sw0TL3uPPRBz0dnQeVtzUcySQR/shRiII98b6lhO+HMdHB
uL9DPdmRvbxYf8JDtW5v21ZxvSXqYzu2QjqnPzDHgq74nuDMqgIjjucUtxO1yCiMQ3b91LdlXRax
LDpKhqdLrr3p7QLycPuVLLB/QdYaWvvPjenwJgIlC+GjN69InLr+79NvqhkXU7BN2vVN4yKfWi2B
3Plri9bfJBI0+9SFYRY9P6FPM+08AW5xxnRegCSQ4wdXjOKhT8ZGsi9fSp3VGOpeiOjIrqkj2E3E
chAHqAjbAhx5qHqs+1wlMtmKVcRH9d5xEhqWmJwId8V7I6B3Gs3b7zrhDUdWgfZc3Z5xusV61svQ
W6YJ8MKCNso71J36Zqy4aKQ1gxNVlzpOUgHA5WVPKNyDQyDhsCfVMQs5tWvWt9n0iLZDWSpkNobS
yTmrSQJbzDRp2OP+nq7udBkHX5cvrl4Hh4fIhRQsy/Ytk1rWB4qDwvEKZlDoloDwOPBq1srvuO8/
25QjbljJO0Jgp+067xwmCyRaHU3lV6ZcQ+IQftWzoS1zADpRMkOMYowL87d19sYa8EEPhbgCYXBs
owXENDc7cXAf3nlV9urnzEHdWH06Q0UEPA9K5bFDdw3EYghCZStAiAi1BJK5aLeCtZrA7yvX9d6F
IabiYNiP7B1XogkoIqavC8TYcI/OdKE0tR6ooReoxOY3++xbgG3NH/jMK6BgU8OPdjnOwtH9PVEz
MK4ru9k9QGoSQXHuiW6TbmkSXdiH5YrJGGqg+cq0rzzRGjjN/1Sjf3IAxCl4nQu5DNVYliATihE8
y7ANZOrb+CHdssBnmEW3XIV2MnOPfhQBmVMZv3tmYVUbFOvJ5FY5cKtvCyrMwT/Xv9rWZLMJf9zG
OrZvojCIJLiNpeJucsOfEIV+iwKdOOa1X/Z476o97q7wgAOsRKdy2BFUt+JP1IxKksAPfo0kI4VU
O5h/KMmsDYC3bi4BDJxw8W9K8l3b68GhO/J8GkOgPfmuBHfH4G+CebSYPMbesA+V2ksgDWaDTbPH
4XrayEFXGPU1zIOAY72Hu+l45IBKJu3IL1B8AIICHVHwzfyhyoQmAz1QeYtTNibSMMSfmXhPeC3S
ujYc3pz+a5NWkEn1MPbfIzJNU9a0Cp15u/7IRYe07hmz3L1dWB5fglYjFBvX7Hfw4VTWMl4K6jEc
V+AKpt3iCOrel2QMK1fEbEx6YYUgVqvjjnV8ZLrJGUy6LW6m++/lOQe2Io0Bbk4iB5i/Voq42Lfb
ScWpaFGNn1Kcz0B6dX6QS4CzbzD+JOHWnLPX3vJqboh+I4yzD3MehPLLe0e9zAijKj4FLrSlVrMH
7MsLZwziVdj98DXyZYuB0APF5boZKX2FEac7MKI9eYeEtlLzmZ170xtIamRjekZtwhxqUJ/FgrBU
OfBDaHJp8VhQPDULkuzHOiJa/+M7F/Dr3Y+g29XuR+Inz1btajhQXzN+EtrQxHuqmoZdXWd9xz1R
DlWlCgbBKlU2BAvPQ7RurtE/A+J3GnoJPXvR6AehFqgWNS4dZcYJ/jUTAejpm5NJpJQdGeqQLZCG
nOPu+SqVTUyZP01KNEQmMC/T035U4dJDu4js772pwDGQevrjvJxJZyUss0+q+SOP2l1UF5BgiU5T
e5UYBm4TNFG0gucFRaZ4+atxriemnGhXFBjma+9kPjn0/TyvuE6bzl8Hnf/LcPMJuVI0JxsG8BmQ
6F39z60wyg+ovMnctK7hMBzOAZ/FNkS9mzfRAfNC3N/xYL66nXDL5sx2kSuM0VoMA95CCy9PecK7
dvQoc5hgLVmgD/iBdOxYBCTK+CrFQpSI53KVdGGlaxkqrBdjXWBNUihkjXghgi/n0g862SA4jGGS
lwnmmaMKNjuykXaNoNe6Hh3P8+pcJe1y7kKZJ/KgKCSG5/eD3uBNW/WNCWduMnFQeeiSf2aWiiZT
wV8/sEtIPyXD4WtPOWSUj3P3W8IWFyKMiwGX5lMkXsje38Zm8Hxk6axx01MidIAKrOAf5aU3v1e3
vRm2j7HgE06IjBTHZa1tDFDFjulM/rkFhPQBfVhtxrbVYWTouxeXu2az5SQKSdKIIz/YCLOTFTcb
bdVdEHQvaUnuiPo4sBVBG8KE31CQQ0JtgE1VIPTUG3QgcXoNbQMbBFmZL1U1osH0Vvb4tEEGxd1N
/5TZK8RNfZwW726dlWaQoGnoEt3O7ahOZeLW/dKJoz9DvuoUDzC7hh5dzirHNoKWYXk5WXqlFsaO
Rk8KqL1hLYZWgf/7j6u6NvVadGSiMrBucoC0Ujat0EQme1hMgCoNHU8Vl8MC/M8NrCeFMgFlaehK
N8jABq2fHjuX/chzkuU9K//7QfsWv3/pgdoseAUmQ/aQBQqu30O8phRk+IH28P/MuGuHoYl8j5xw
3vitzPtBAtUkhbIsorU2Ht5G2Pt+K+MW4Upn5c4CjneiWxBicManxeJNU7Iq35KLCE7OKE/q4VM4
kQgVgxjq1QzJqd5Xt6dBOZLilisYgqdC2RAqHRuFJaMt+lw9x0XiMlvHANMHq5OcUiKMh/eBxv+A
RmN3YWcZwdvpdnDqOwxp5WioqTBLOMEohO+UOn1w6kih3BAuOxxXw3jyqiEhRA5Q8dOruXCQsSNC
JA4h5FN/cylNlMtxDom6+wE+NBu8Esp2I3Tz3m2rfRkgGh0NGUPokkhACvJ3hPKLfJ7A5zgJOkoT
zdS7MxjnKeEwU8uKKs87UJE6JZOPAx5HcIGoBGtVAON7phvg0BQ8UmU2cVjYSAoqOpWHbF36rpPd
xcUZcKvVDvTBezWg/n+iN+D75oPgAQWlzdMzX+VVZGXHlsB66j3JxTshGSeZ6LZoSMYkps8dW6IW
GWTkntolIzjoGNsx1U6rVQXceRqEqkHv0mxGDy69Iy4lITzV2Jt8TnsSXq7Dstdx+f9s872Bngr6
zxVuVaYe6NtjTJpHR+ZQuBRrbYozCBjb33oshQMR8AXokske2xQwL0Rg7cFMOHo34xDtgVNs0lyn
SzkSVw6ees/eD0MQmMSyKLaE4l6FDCVO+8Q1rfbUf+vCEEzAREouRVhzRUvk3S1W5sKzjVZW1Mio
q1FlL97iUgl3w57kMk1E8OtFC/8Go45/dJxHDPyWuMvbIm8LxVvukm5c0Ehxr0eXfzCUVftGwd67
SVdEopi+PRwcS7HfOGbT16BApUdrwNSNYcI6eL/Qw04H7tWNUFgGUdN0kAWuoMExThG+jn2I4HhH
RZsVCdLhoR8iQ5TdNJfa5ftY3qoPHTXF+Dg5wZH9SUl3+HmiRGNwACoXoz25C/f9tuCRpBShvKGB
K1A0piNGbb1xr1IWgHG0ibZfEhzwZlb3g5kF7bmqUYfPlI77b9BIsnIpYdHx179MVLavD/pqPHzB
tgy37nUDXKCJnbPeTiGSTdovlHFU+zvxUup057NgoFAG5gTK2Up/V49frhvSrAAvSASLO0vrOt+w
Vo8Q/Ke86uvR/EDXMqr9bCBwHeu36F5cJGp8P3mVVMvADFs/g9cdwVwcNMExG6q3i8/UxN1xthob
rV8WibgCDJkN9KivPXDwhRQ3YScWOatZaLfBnHO63wjxuQVm2gZwAKOdbyjymK5o+g6Qycft/+4k
iUQ5Wb9yk2CayG4QRe9bTua3LdkQnSkBOpalYYHYtlvTIz7QhR/P8/kPXLP1GKKLfJrQ4jk7yiqM
XBwP8kjrf36tOg2M44BwiVm0VQUMhHZtTzI3rz0LrPCCCPohU3nVFMiLFIJs4VuVXSncl4IA1hYf
fNDRC/TUlSS7BX1RVLbCqQQSA6+HfpZQyavJhlmucyvsLh/IHTfbNYEQKYchvxllnpa/uzJnAJs0
KPw37Jql2jeljaLQdkqZR7z+3e9E373U1UgDy/hGL0Xsr17I16xw3ExZmXyrZNB0lQTGXncP2z3f
yMD1WhvBrWBvrQMEVCNpWFTFS4y7zI3FYJLhKMi4tObS14ZHkko/XjKI0TsxCcc5yVD5JaCLb2LT
qeaXEdHT8WF+OO/Ar0VdabIfMgGv+VzOlUakn/KnUR2rQt6opEeT5dGjvR3DuaZZCwtMnetNEKmw
3LYPw6UxAU6KmFS5b9btsl7/cZ0rafF/Gq0EnynIRkr4na9c6MWEQrqshC7Bfe5a5rCZWCTT0vMQ
1yr+bBN7sAc6qHXDx50L9pc/4U8Y/nsvXhCbv6rCT7eJZl04qMWzX5FvY6JyzPqPIzhvgvmw83U+
xMocdJkELtNoOe3taH5WtC016VwOuGO0oN0jeyNYVuRlnLR3tvOLZD7SIEizegBH5VCRxtMX48JP
b/U06LSX4Iw9PWm7FjpRIABm8hj5Awe8w+0uBhMy/zj2REtcIoOzUrRCI6f/ljmRAJXFKq2dD62s
/fvVVKD8HqcCeqMjyXSXJ0zpIMRG4LHKe44/lu2Hx+kuUxkOsoM8vmYiDvYJbJ2/OqsloHbJjETU
gGHz2SjiRrDmGJYVChX5X4V8JUV7/DcW6QbJxt4tFxw8lHXabKrCjSr7X3/odh7n4KXlcYXdx7k+
Y+/FQyM76xA1X901FUFqMMDN/Okmr7va0agASZ7nZSs6yDmi62eVQRjOPI/E40MkUhDnJT5McREp
zb2FGXCV9ZwOiDN/HbXynt4MzRSAd9tWyh9YbC6fEt/rtBCdpzBdN1ECmafHn4ZCQnbr9TU6FFU8
t92FUSQ/DQGmmlM5JA/zqYAmtWf0E+zhcbx5978680kvxB4kpzWcW4T3EwqldJUQ9Nc2Y9udUqLP
mEV+L8S07LzgKMAXTBO1R68QMUqi/b8AlUYgZsmlP5k9nF+Uybvj1yl5lB8bM/4yJ/yXpIg7pGID
VrlXVdLL8MR1DMnAFqimADEhKMG1nECG7l7r7fAu4tXttfCBK1GwrlYpaVs2JGApkmto97tAzaEv
JXed2mdQdhf38wx1alKWH0ikjVdFqfxvfb/Bb7LVcLOABDAIRHE6MJH/BPD2bwdH2aEXjW6186mz
qXLao81vTJ/31Wz55SgJ12rTBShUc/BlDZ7wTYItA4RY0whlEqoMJzVmH34zMcOkBxRQaOCKpC5r
RAcLkeBke873Oz1CtzDskwvonspNFrEZhAr3fChnGvmuj6xcaxF7iwpnl2yYqcSKhFls9v4q+VtC
+kHlf32t8m8ftpBEYScJoIiaR6UPlfUBSGkwnCBXZbxbJdnoyRo53/+T/lSZEDbdbQwfJZscb64m
NMObbNDQq5K5OulQTiGbi5OeygzdbXrrLU3PX6IaaFAZsHwezo6Qu6SYZo9TMB1fY/U10QGmV2P6
SB56/4Bt+az6t7ZaU4bplap+A073uLOwNznQUO4PUe0NHQ/trDgPPp9nXhk+uqZ7apYrsHOVyqje
i9We5za3lGPNQVYo2kWcYT5NTSZsTfTyj4rS01MMIa4mb+gBrMo0+MKE2fogbFlBW4vLo4IdhWDz
YZeiOhFq34pSbthmnJROseeeZsXSw+dMGJXhdiZnBUDN6VqvsM4JTqiKn+kgaaQDlsxuMH6rJYeb
D2yugpSkMxSx9/9PozAj60hR962742HMFrRUxgvQV1iQXxn/nM89f6xdv16dAirbOy8DDidm9+jj
DLhPmNEysZakoY35wAhd1SJQ6Yh5eqho5Bu2VA5wUaJQW6SFyOwqBexzq3U1nmUmlFh7CNObqpM7
5ULbuISumquFmCjL9ihVxnux3U3cgycxDRLHH2O2livffUvrQn6rhJBLygPDCl8+9gh23Qzv+vtr
jcX4GLKOVLAP2k152tgoV3MlkL98nH8V3QKJO4pU96dCfvqzDO5KZTsUzFoWrr17vIRcTxV4S17h
Qi94t+W7Ojc58z1msvdgQCjoweqlakyHK7jaO/VpzHoaaXfUbFQG20rnvqkBHeftIs2fT0+G29Cw
Vqys7GvsuBDhDopHX8T+vC3kKb5VD10OVAE1LjIIFgslK9I4l2+VQPsNlVpnkcryE5lSIMWUXTjc
MCvIFbPoywXDyVjw5cxxKcionSrY3Q6GR1qSK1JJUnbWm8p8Lc46DRkcUeD8MII9ZDji80LsyfO+
nbovwCpgOSRDW9l1U+BHKG0zTx3fNl3aUri1RPyRIY0fxCvtodKe53ROm+Nf2+7BaVjliSqe/QY+
1RAAAlQXBg1+jFnWbDZfNRYTG7bXAXV7q+q4VWuLdSMt2qfmE+VVAtuLFUKZ+IGjXimg/xKlV9pu
D2gqxz7WhWmmrp1fSL5I6V+h6mgAaML5CPCojatNPF3kJqNWyC+4zcx9g9iR5ZoEIeYAbRR0Z3GS
LkhHbkFG9EborMej88nBDtV+D3M5FL8WkH1P2WrEGJuuHnq3IUQH4ynwjEgkNaxJ4094lSpFH649
M4qxjWuU51Q4Co+8DMohWqFoO5C4nyCZ7WYChvV3iqiyleHiVrJ2JM9Ct0eL+tURIgeqYeY4mngL
ijfy9+l3bZhT5Cq8MYbLM1JjBRVK9jKoZvS8xvK3ZtbNz3bL+jbmC3zJnTP3xU3CfWS7r5l0ICkC
4tKMRGFho72AYp/i394REgYReQCNCcQhTQiJq0mntu0YW4AEW2SLQz90OKJZj1x4Vt68TXw8qzRk
UhbaMjRFV6XBKEfPc4hOyfBWwSecIH95DviYtyiTxMygaKEizzEVSN5EHR6Q6+eqClAmcJ0CWO4v
DMYT4Un1fgjO5K9ofsHxHtHVhLPO+j+xIkaGHgM5CJTPbVwtBoDib6uGSaSrIqMQgoigZn8QY70j
D3y+OeF4ITeZm0HdUE+n5TcKlPJ2sTUcvHYpact1GxkjJcNqJoyq5tXAJLnw6IxatbnaELj0C9VL
VXntnqK4WIACVgmKzjMhd/aho5hi1KoSSCjHNYNmvl1taeQmS5ewhncz16NDaJUXv4KbEyygMg1X
bblooQea2Givqu4WYDI7gHsoQCzBCOxBDmPB5EliVXqQzblkSvm5Xt9LEQXn7c0S43SaWU6zfIi+
tnb229Jn9gjawIzyaj84p1JEO8Z6zDy2ao3IlGKME5BlhymM+/hcO2MuiCvL7gRw+OI3k47QpOJx
oWCwvw2cSxwTfpKYkGnlCvc4PrmiSQrewVX8l/sRHQzsAjZ+ZZsK4fO8TgKu7RL6naRkmULrUK0X
PVFTpuTlSQnIguOSH0XnkHjQRBK6zQmjhtUuoBnK3ZZyrlfYMFU/GxcUOcI27DOU43lqVqXQcVSv
/QDOjFN45jW+v+saI0hwnzoN03Y92nacH6J3cN4RaqmmgPCTaY69hx4rebZMzCqtONXeezzPAVCp
3UOc3UsiYwkzIJcqf3ei8cj4FsSyOwc82hod3ZQ4J9XIeE2pwlsvPWUoRqmlAsPT0rvZdICNDJix
pIFdJPTha/m5DcqR2WjKxqLlLXjU5GRZy2TahrurP8qTzT3mkNKTtnJf1eRcVONlACL/9dSCU04d
3QELNEXwGlNTkS9WUI4hbML0uonZPXaF4DHA7kWGmGCEEVyVDsIIyeb4N1i0Qd/niuMYnynT470/
o5AQbmGexIpitTMc/CoNqeiQ9HdKYxcIIPcJdUiy8G0FdI0ddI5WuE6DSC8Xf6stMvEawwxdcxbc
2y+VNAvHt2y++pd5JENp11QGZRNkr2dffqjUhrQP3jqri3oVzTi2FehXHIsZ0rPoLYgtc6sd4YtW
vo8pTS5DC7lpUG1YsD5LiKWO2M4yFBelmf93ZV4YReE/C4ETn7lANy/EbrVqKS7iZuspJGJ03gi8
13ewlH4beMyrMcZBiiGv8jb/4LVTsO4lDVyFjZ8kTLgb4l0L3nafCcHB7UBQwtHEV8NtGYxP2U8G
sfs8ul7xCrz909GpXrna1euYCIPDnUfDtsxso+vgS5Q/8i5PBkiFRsdiPECwljjGb6MfeHQG1/N7
geEZGHBuvoSZBgqVeJxV7kkp91FS2kJPx4i5ls7MLL9tscRKJZ3cURvQw+RH3qtX9Rj34KdAK5fa
R89NnR4MvcAIXC5OidpxBCCLDIuDdIxZHp/k1C0YPb8QiuzqYvo+jWaIEoCci6U5kVyR/l57Jiqq
E5OSw1/I3s2L7lv0mgNwKXt9C+fdM8ZCRwj5FAIxOL1la0tSOpsfCsTzq/o2OmOmXggCat7XwSRk
vWzTO6qX0oN9LwxVeTHGPgaTtE22k9nzlLnhjyuVtFWvhJ6zo+WHuQuJMAaT8/8ZSsO26BOicJUk
zuEu8K5iaH87v0S4ZJU8sqTVMVzN/5T431LYMDsiY/OBEhcruJTkNJRNZlF1cLbfKf2aXcslRWcv
nA+Z0eTdEQcN4BvOsvFEYlLWIHolSQaXNXjuGZ32ztn/zZpdCjh6tcKgVYUV8lZXxbmKV09wpmo2
RsD0Jui/yL+tI7fhujDF0Bzp6yV8lYwAqBNaTt31kZ4Lanx7x4LwhPOIv/ZgBGeMh2Gnma3Z64Sd
PF9JLzQOHDHitnQemsDxUVhOjW12txcW+FhVeueDFyA2ZzI2ZUa8faZQoPouQvY5FI5hMoCIjYvf
nqexv9JhpFTJR6uIsJ0UOAGnDJdhh1HF3smHG6HNcNbkP6uRLmq9NDr0BNdGEveyBFn6mUYZIJG/
dxBY2NgyfUmyD6RsvwwOK5t1su8g23wSstEC30YeeQEmEF4hCvsyEYujb0N9KlnIu+1G2Z9R71i9
fZxq4vpkXZIwnrpjm2EJc1W2ZVGAPj/qJWHDyyyh9oha68Id3NOadijrf5WRRka9g0mksPhCIAJx
hrDzjqnE1w3obN+9bP5BZbf8JHGtbDs9ettrQWnHaXn3gTjTFnfw3Vf5EjSshTEpooB/25r0Q8U3
yhe9xIDqzlfG2+LjK6c7CyI+ZN2EKpKfczDGZLSS0mENaYGKxQ8a7k4vNm9yXUqPhJIjs3FZXkGU
8T09Pk/mKobpy6uAGyniQMEuyCreZ7DZv9KkIq6/35d56ZUxVKKxPgu/CAbfolhRGR77le4D5LCE
izvvLd5hfMvfjvIl0F7RcfmszHB3hJhKktW1gOCOLL2AY9LFFhyMpYRcWYtFeNKJvOdbQ5LnPwDa
nOcuXVj0s1+bTLaV3uqvTB9xBzLwJYlK3Zi9+H/yj+JUUA2EGiz0ziWQvoQKRHagfjugCi0R9gP1
9pIW1H8qWecxkQIr73Y3kI1dTVTAYmLSm7g9qyQEPxn8ar1yOXTmKh4HsXE1ldttrVW2ZNxKupDQ
5U3mtK/JtAPg6pjBlgDb2Y3GJ2LX7xg5lGCjTUFJMdKxdnLBMTA2UMqrWrBGslHg34ZWS9PAw5aA
HSiSnU/fVPS1ofOPk6+dhRtyETxqDIz4K+XMBkcsDijqneIt7q6q5rzjWMXWcygiyBnMPkl15kd2
ytuLzA6v9qrLMHTAlEo8CaIm05Q/FyUzi5QdKPfLHXZcwT4//J9Blay4EFKCnq6a5LapwK9NC/eH
rg9urUPkKCEZv2CggisMVr7w5A4uSpY8JMLNMa+kyGWSYqgNqfy/uQ1PzizGlI3Dyv3pupzjV6t5
5oKwATHSboCeSW5b2bTixrD+E8fmQLFFFrtjk6de1OZsmpK61tp8jEmP5ohtbbc5btRaB5cXEEya
gWiLc1hM0ZFZA3RDRQhSy7C0phZj6xbMsB5x+3fbW8XCkQppbD9q/uxzIIjKg9wvbR9Iola9JbQp
2+r7i7JIkY6ttJ8EvpZX/uxECD2sB8xUH6PVirjVHO8A3iFd9LJpzh3rnWvLV4dxvh+loOdM9NMo
kQs+0AsJZNipZX6/b8etHzAyhSnO25Vm7DD43TcuynO1EAsltPr/p127lyddq3ox/dh9QS4J2lKP
+HbvzrkBgzeABefq3SqkhhukyqpSlZGj93seWaLTdmTTQQ9/2mGeOlPQIFGOWQoChO2Rtkb2M+xG
szoQhmHDiqaH3y0dxP8qHLviwTSiu+zkXxSLbJFExEMvf31BM100ZVOIZIYAMHijODP1Aot8AJ2G
1Bp/77I3qhmDL02VDZoLhn7mfHQVIjLFb5nMnXswpx94QinyMcmd+53AG0TWPB+Tm7C0evRk4fZA
Baya/IMx314s4PA8PSTGbofxU4UfRckx9G/7fhJ9kusBYn8aNf9QeKEyN+ic/MVqq7pxGK6sIoqm
+sYAbPI/aeK7hlDe1mDBjDpmpeeRaPO9W8z1XyL/saJ0nf95iaTRhF26UpaTYGFxiO1EzdcA1RQF
TXF+8eR81VkLARmjaSvSot2NgpGHl4NkKid7b1PP5m9s2DlQPIVnd4fMrkWX8fVxYGgkZexYZtq5
QFQDozmmNaMCUZ1w+zTJ6SZRxhPfWP7b5UbbKWIcyB/W3N3yG0IIIBLN4Q14pdAdnKIK5G7w4r5s
cSpUyct+SASbcGbha9cbovVDOITY2S3/te0DcznO41xojWrb5MbqStiiI42NWbyNDpzXgk0fzdcJ
9sJWDqtDIBEbCDD+SoCvmWZo3R1mMvJz7zTD9Fsxe7J8y8yo8NZZZaVssi3HIrJbYNw2LFarAVSI
qNu6pp8Ivt1/BGKSTO1eTzVDbAg/kDcAX5ElSHLzEvo3iDiEZbf0AD3KbMwqenwCHvnuz2uM6ARK
Re4y9efrzbqHpmD50LRlFnPqwIT9rT9+FVLhQLnltrZpVxnPlZGJE//R6M9SNRCoy3rkI4hCpvow
Eo89ePEonfXy7dRwSB/LMlLWXzPwumoho9+UDpKOKpmHKFeVl4PP5tSZjMgwHKYwUPREMvQbXLQ6
H56HWZ2cm5Q+qFtH8mXszdDA4YPWvY0VfZRbHzKCPEjOU0wm0wpydjqIhXkduaplVLuayyFzwdX4
uGnJfRB+JR5pAaq6CXTtg0KQdSxmFr+VQre9KcLnRQA+dEYZdujpqHTb4fWV0z+y27YVxU+RABbi
mDueRWLSAchsrb9QLxZrrPYanhm31w+QeE6FF0LxzHzBFH/2ConLHSVPhRPYx0usE0DvY2NZt1z+
BGpFL2nB5gKxNSkOARkqygAE6D4FRAfjzE/HQ0845bURgJIE5umoTxPgyU3EiAyCNjuzdRTC3zBC
4ZzmbdP3giAymB+p75U/S8Cz10E8LSgllMVe1493mhIju6aMMOBAnm9uJ7wQAfjh92lcQ4KclpQB
7ekIe2XfdH1QP95hH1vPOYzU5SYDcxPIYTTRzVgsmLqPKxnxkeF/0qchiYryF5/0T4q8S6l504TU
mrKrwSuYLjnIEkghZkzcra9JN/XMgmCa8qHnWi+33XbNA0TfCHJl6eAxIIpt/cikqxUrmTYpdh6X
AKuMn4UwioDWFaQUS5G2rqZMdW59hgVRlWJpzwKZyIS/TZ+4OHapo/RUDlzfk36IpDMbz5SdnTQD
+pc1qOd0sI1l5wCagEeaR75ge6eNxP+go6zxntmoMIXQG2wVLkyPqLT/OUXq4kai6iSwkMzgCFAg
hMhcJEIolztWsi89SL0+RlovA2DJeET2L4IiV5kWfTM5Vq5bwcd7ebbUV6SRl1N0IMoHmfZNODyq
eNmmFHR7DXpmPc0w1P4K5yIcnvdlqTQ6VNYDHRddx3wMkFPJ9eZQtRp6zivAvdguhCFfFF+1x6iq
xMYdIbGWPdVqJSS3H553EMFv8qgBO6A2BVx3bW/vtUwWARi+7TRQcpP1Oe8/oacLVkWQYngm0vqC
/G17haX2asa01C4pmk4bTEBD2Tjp1VgPn7kqXj1hHJ4O/V8fOqkm6fwQ8lGi2OTTKoiwviCS3LWM
yHki7RHaPGIAs84mjMS6O5ihSWTmR23jQ+Or5U7prLlDhn9ChgyKAdAeGClaGJrf9KQJCo3yPAg/
m96rhR/Z/54TTBZykdYpje9sEutTWSe4MUCGhP2euTUJBmyJvIOtQBfFnv3D7efNecK3k3N5+tOt
S8JAf0moVylTzOOv5IRUoMmzRjkw6xg0XaqAo/jgv9ADHrRxL+N69YcJwARWvgsITMwFFO4lS8Dt
2M2IUSUrQOJuuPjNSOZI9xGNFaILoDJ7/6omLYwmhbb4XvEZWEmlPCxcJe6NUaKaFnHN3eEuZ/kB
RGHHbQ0+DlI7G/NBFxCH4dA7wYht2aXwpXT43nFwbX7C5hV7xe5GnGb6DlvSgFniqAO1ecJu2EDA
QbK4cqrvJu6/qwCs+kNNcls+VQJpwl4j29VQydnlXKXG8mnEElYnhju2ZGA/+LfyHD6Wxi0Ub3LT
+7+h3ikGeB2LOFHS5FBfhv9yAH1CZ9Kw4L/NA22wVjj+uj15vQ2IF7LKTyyzpbsiapENPQwF9Vy4
mHJgD8vUIyDnYYoy9n+0cM93hkl3CXGL9hPBXzaksIkq/+/CKWJ/UWdvYYRmSD6JzzBnokdQzSqr
ObMkdHnOj6eHYpt1rerAXNb0ZBSfzIfqxkSCct0ImYW6QqGEMYKBePJXAFbosnyLdWBCDxcBtfdx
QJtmUqHWwpRCe0yWV47f2uZpGKTpzAUIwdOn0lrcJfE4/Jwsw2s9mTOcWALoujuY0iVloi3wpO9M
jhjW6rC+GvqMQ/bSkUNwm/RJKNJXh8NDmwbxu3S9EEjdlT3RkRePnwH3IVIY6sU1pWwC8zG0R3k/
r5TgPkKC3GtdZIbytlcc8kqqOXql5KtZIr+TOHEs+5U1AIcKqhGCz+Adx/1ETD2zk81tZsYePeMJ
KLLTyM/l6L1qBnxFI6umYxuNqyKVeooxa3TSTDnp3ep/gLTff3M/CD2LmMOsZQZ+ZshWsXY+E6EA
tYxxZyP6qejnuvQ19LthRo8OAEJMqp8gsJcq9M2T3ts3+ZWxyjGWchd0P9yf5VqJU3rUrMKAqzPQ
3BBQu8BaWEnXTM5fOzIatau5AUdqZ9VuxUfuQMcTJ3LbkegHS2M1TUMrfwjWJLxELpFpf9tRA5XG
+YO2I3hIKUFFue+tXrKUqK+0GhZ32wcluHfRo1244KQx8Sivdr36LKkIA+wCXCcdJ0JBZh+Yw/4d
tvphOJ2Nd5mkTppAw04b/LLl26JTYNDwgO/z0nnjimdpUfqD22qcWsZQivUx+/DVJgOs3Pvp5t4G
6eScmYozSCtPWzoFbnIxO+y7q8mvHCPd9GVu5dSRKQoc/mPVh54w3xs2J0HpJ5eJYUrlp4pOMMa2
xhlc7HSvwggBW09w+RMv5O46pXFobt4chTLlSd0tUz9NvPQOiugwXGzDA+ts/6Bzb6xBQBd2a05H
TJ7socnKmOOMgtdctQdLpBhwkSKYQWE05uhNaSigVN2Q7BxVU1BBFALamWmrp9X+2ZBPlxgwj+gQ
Q/684roJokBZsvxaLtZwFxPX74MVeCz34cDPhtVXHbZhcy7L3XcK9JV3mEnU9vefbV3t41HTii75
Z4FZunyuxX+16qMuMnAUZ6vm+uPzi9TD4uEw/xdKBiKabfO94iS8K/hrVSE33HDyOaAm7edeRzYG
WiHAoZkAn2YV7evrY8bGBKSE2R6tt8pjuPNqQTIAlbo/+NoM3FPiTj00it+dRRkJjD+wKHy5IRhk
rHz6HGbIdDHcxAdMeM7Dc80m1Y1tBa48hl+ivvgXFJjjZjL1kbdsbw0J+4oB5C1GMQSG3LbxNVxG
8yL7Lw/hCIQCcQwMFHOFWWPXN0Z49l3Hx9yvm3W1/mC7vyMDxrVMhVe/24bPpKshZJIOV7m9BbJA
6+3XoLbLfsqpbJ9MJCTOTWYwfl8et5R3OV5aVA7XrdL6z2W/K+eFktasXYj/UG2WXZxwFB/5PEh9
UEUhSfnuP1gn9Xe/PpY1R0DMcMp07fDfTUzgDnfVBPs1bKknSOKeib3C9JxBW5gGWLHiyE+aYTRL
LbkPtkhmlq89h/FcnzGQzNx9+hgQkeyCIX+8zRHKqk4gi6wnMcOUGoiseAqRrFEzs5na0IvH0TDc
NJeViXFe626V8QeZZfS4UBMkfgeata4VXSMemtvNY6n1mtQpH2VRdCQfNfH/Bj98aQDaDIkQU1ys
LgTeSIIjibFnLTfo+lPKCnxIkD5zjr5lS6r6Yp5PerWMXrTSJGh5sBEvok/Dc3RcLWuUAycA2iIj
1cpARA8EDJXPIG1z4FeXez+87tajGviMx3js2m6nsU4Txh6j5RvIUuTz/kbCOGvUKfgCHxv0tpPX
pQnSkXxOTjwyROn1sSG4wcUv9llCngOR3xBZ/KrzCn0ndcoaCGvKXb8tU9GQOEoanI2bfF1H8DwX
wXV3hD7/7IaGwKuFUycZ4wyGmZaD3NK6NXT/Af47PMez0pMSdHHXkzyX96AQ8qgSP3tcmuGQ1tnw
cZglsJjl6WV8OZ52LNbEZ1w1LXAmeg/llll4H/TmRIJXxxxapRCdwqobO6QdBv1Sz0LnPXf1nso5
uMSl87ap/6Fn7SGQ8iCB1q5iRXfTaDd7ZheiDMJ8uouWKqemZ+DmTSKFMkhif0NTFgebG+8dxydy
YWABV3fhUFz+xwl260673NyT1FnQh5RQ5zJyliM2jjB4peQspTHnSpnUq3N1nuVSxI/IbdsAq3AR
K1GW3rB+erqsECz5TKoFCjc0j2yLs/Nyj8n/rf6bxZLFJcCbIo55v9RRaQLdaTpcn9om7wddVkK3
bM1XbqIhpBPUe+6HHzQqrmvfWeFmBQva3OdsDWKAvi8zy7FfmyUK63TNiE9wFC0DFT/1HJO9J7/y
aoKweBHnu3ycN65CEWYV+azlw+EDTbfnCoOWJhPnOyS2GtmqeiKH3JaHvyzgo3BLum67KGxwK4jj
wcJYk9twnw1lB8MzQrWVuPJhY79d3Wwvf4eDw7WEnDikAd3cIaPSPfI53LN0z1nN35GiVcj0vJC5
QlMtz+Qzt6DOhKoUdvgVxWDdRxcRqtT3j6c3jNAbPkvYn33XZy1JrY3YTRwOQjcL+1V+ZsCSFENe
CLNukYO2rsYEp4TWnVogVzsYNi7DSvd/PBWfu3CHYrvmLMuxS1+3AJUqRPZkEk4kORD0bgelCu00
ftBtGSkKlNFF302LwdpSDDlhyW+K8pXZdxPQcPjr4ZBeUpKlHLwqikHabG4KD4xRLvKa3+KzNf23
Moznu9PkIf50K0aImsqH8Zk//Zb+xrDinnQvf1vmXY/OXM/JFnoU7rVQCnejoTONmIjo/4zj4zTd
viroSmHd1auVoBwRcqavbngrjMA61uwwl5f7E3AGdwDZawp0czHIq2Xn9j+R8olAhqItqgxxmxqk
CYSqB9/eAPSn9vAo1wI34ZPvRPvGhOO7R7E1UNpInGjUq5fuAyoe+8xvk8bjOzPxoFXNj+Oa76rc
hTWeMaNPCSc4YkDXozx68W/tWdq5+f34L0e0FVkCFHNsgfXbw5/IgYzQQJlQFhmUBnGkgx+Wk5Ut
Rb2eW56GdVqUA038osaHECH2dvLJFqcSTLkaJRBdNfpkUj/3y/jun/Hwr/Z7+m1W9C8ZTEhnNoVr
3qDtB4OTLT2b5uDptoWNHTCpqzs/ZAjP6yhbYf0XcjeFndXlKaLzykYWXSEx6ABvqJ0Dr7Q1B0dX
qAM32ivuz+/hru+njlFvrHXo++pbXkeqivpRq3z36xAJdkX34jbw0FbStE5864qklpDheIIlFsIy
9e2kiYSLhc3gQ+rNsAfmXhHS9uy3YyvuSihU3Bpd3ACvUHz5NsIQW/GzPfyet5hCQj8LUiV/hSPf
2gonq1wU+D+PD+UKubhpqo6CDoS8HKZVFlS/eGpt9SD7Vsuq9qlrQS7+T9r5ORWShwR6bzlr+OKW
rJBXo+ZuUMl6DfI/1JSxb+am2mDlBW/ol1Z9a6/5nNsGtFmJ+hbV0HBBmpVCfxQEidUDTI+efJAD
pr4AZI72Pe4hTfqsHXEUFo8ZryqHbtYXFb4SlY6F4wTtueJMZRcHFnhvkO9/YatFmrA4vEuxVPCM
wUhkaAZQBokF6Rkj23a0jgDnRGkMVlkR9X4cqLDgJYaAU6IHBkZM+GAehMgVG32RDWTxcqZNHBRb
35Z1S2yxFYmUSLZSD839HH+pWUXAEMxoP0zlleSmmZEBPPlF5uRr18e8H7TygLQ6QTXHFWU96+K4
FGKs7D/kmxZs6SwD+lMmVxyppZ2lqlg97BMQY1O6pLZ1OID7qrDpwTanXVqIeThSbhlp6PjmkA7A
QWsi90FGWx5EWVzAQdpUdQeXqB6XZ5hTmGwADC5XwWB8I/f6OXJGDQmXrMdeyVW9UOAAdwc38ugB
pgCILg3ikrfTVe6YR4AX/22BEDBzB7VJoEjZJG+6CiEQ6/EbVXwqkZdCLoYF3+H+Ksev+xZCwici
E98jL2NBPuXz/GL44Px+r0udal5+XYMSIdYCjID0i+lpneiCBlSLuCSvSOOkPYDJe72vrq8KCoLB
5HWHDOpj8KBLoStwQgYdl3WBXHmQl9B81q/UL1pSSBN3mQBml3I2djfBSbfpAxT0xTiC7UeU/ga2
kPcR83hBjT6sf/FwrP/lx1Eh367cqVrkDa3RdrBwdxgWxRx2f+uSgY//TjERhjs/gw1iia+gsmyX
vQnaGUEqaUgFO2IfyOCBurui8g2E/lhXIF9ULaDKD7kJUenphAnDp+nmIOLUl64IuG7K0s+laSL3
pdpXGqGlr488pFeAg67/klxhGY7dt6p8+GkHZd6Lw+wPDy4T5VNEyCYXKMOys2U2QS33+7mRrXoE
/VwBzXQvEkLnteG8aac/x6RUY67tVywqM4P5MsCxMnZtx8Dk7CpW9vD/2kX8BkQyGH0vOL9KMj0N
5XtXEVdBIhRQ+N+St/A+y4YcunRBYcLTyrPxl14CufMIAQKm/UjpItZ3g5lvkNsaOhcgraEpif1t
YeMgY4OEv318NrTxvKx3yLTvr/GRPbc04VVHdjyZNEiOoh3c8LRZ6BlVCy/QEDY15GI4VtCfNwO9
Lr+l7Vn7dC6Bx0GA4KaDK4XKUTmVtVZ/UGTiTLH2gokZZtHIrwyaF/YXmj59BjwjBdfMAMXqufXj
06FN2G3j9/YMWWbXGF2R45BCKU4palIgbUqikC4AjmAjKMBdtnfmk6qB8SKDOB+zOp3P4axksyoO
8YZitCgW4Vp8hxHrt6bG82mPk7ICMyhL09llK7k529Kx4QZLvZ8k9PZk5m3D9uA15blnE5Jg2Q0o
bnkVMrtAo4H858sF6IneQXsE5arZVY6Q+3yS/rdtu31ZbAQaq2PvCRZ2MOcdvyuJeZiWt2A+XNL/
68OiU0joi7VsB2uhfl09PbeOZA66XT7/9CGV6Ny2LoF8HCjKrPpKpTUOS8p2ZuyhfclfW8WkFDiT
KXQJtoCOxcXbZMwjacLM9zvgQ1jEExwaV0Gh7QoYJEdn+g9IePQ8Ys+WfxEQuQfox2HM3I5JAZ9V
9etG7zIoapQLngCGxI75VIzdD+XkKzQTHODoJ5/W9XBCGJVu/hvPqDYgJUbl9iZfKhbEUFe+ej0v
nCQYo1OjMAusBoOgdfghz48mJ58F5FS0lqleDcd4uoun0tz4sSBANBHk7Jd2RggwVHyCO6zV71CT
suXyo7YQXvhsIFdepVemDuS9L86JnBymULleQTmTQBhVuICihEUktPDGCfoXBqgu32yAX9QnLhlm
ByqxbaNz6tEzNoa9dI+XrWKMgOhD14hX/T5T0cmLIKujtjd0xAzE6QONAAAXJbx6iYx/XGMLw5cD
MvYKwDD1VpIs2JH7+vBElKLaNc6sPs1HOeX3ZhRMMPeXpAhplJRmx+0GuZtu9Zf5bkWUTbFOo5NN
Coa6uJlRqVkiEZEIGCf0kdSjo1xZ1EKtITMWdGb/xzQZk30Jt5UsglgRdYB+KyQdLelUHZJyqYRE
W1nWiIccES4cizYVGcgzBqTv9oNnXYlcSnPT380Z1hHaAxaYTRcDlfVHdP9XYjKieDuexfJxkWRg
j81woBIR1YeweLHT288rZUiwfHBXGPlWxGTN+SAn1q1c/Dcx1PTM83DICaP6jYxT4NH0j7xU55Jh
xCbHNzGS1cpJqDPcSZNXVxmFRKFzP038OUMLRQZFBxLX/PKawF6MU2co77EBvk9WqGwevRNM4nR8
p63myL4CSMAOpXTCmR5SOkTpHREuNhgrwxHfZdt9c3e6Ye4xsu9KqIhT62OYtjZOb7W0bgaB70Zx
7oHjGLUfMPqVnCvgfOtw4uo0jq+czzEB+UCmapEY8cG757tv7mCOV1B/g5V4e+6FcrApOE1Wu3F5
bQcyUjjukI3EfhwW6xpDKNqFt6IXfz2lh0P5hER+U4EufqJG1t47mp7p+HK2QidbLH55o5lijZ4s
u4SZMwFtgRww8BwTxcksWDYOQlNRLxaLnmdnTOoPrtkE8L2/iCQIYMmm99opS4R7aQWAitFepEag
5kRII4Z6cx/BISFWfr/AFDlLxyi6PW9hp4CSzYNq0JHcXBISvPc0NFZkv25izppl8chCgAx5KHrT
jenHA7E12YqpCw2NS+Rar1cwGeetApQI48d5ms+KtLARvXipgoKWG94yYUHEWKXTHnU1RBxMpdXZ
U6ugviieEqBobunyu6Q/FcRfzsz18BV0VkKri5kzir/TNaf5rMdU5NZoYGJiFR3nulQIHZYxFOrR
mRFSRXFRu+Wh4e8vw46kn23Y6bzKIapWEConRN1REqtK/dhjONGdP+o7vbFuKW5TLeRkl+T8Doy/
SCQg0gHfcKq5cBGy+BFKK2H4SQ1wthoEZufJ9uaUfuntxZCVhVvvGMIfUvkMfNgtIIQDKvnU11aT
f13XXK94TH+Kj98JiyLAPjebRIIUC7ZX7YpJUzB51tVw1Djn7FnXlDQ8/dO+iMIp07742FYZkW57
6mog9qPHqjBlxuhJCeznMagsrsGDqc/PkkTQovEbUvYuaGvG6V+si2xDfWMT1AKpWh4xFtUyYuuQ
3fE1qXzpUlJgEPFg2ErE15Y2D70v3v42KEFPf4ZfiLBBSUqgulLxkKDzvst/IVxDKaWB1TImzvG+
RH0/oL2krO0X6NVnoh2TI0FPTv9DHjoJMbVc34qKjHSeUhb5l6XDtk9KUU9FTBn9V3EsV1Beooz1
edNv4UazZgCBo0Tukn/lDjm7zt3EsdUSxEexOQ4KD2k2n7rszgyxd3YYYglvmswt1VjSMgbOseJd
HWhRko+rLP4cWb5O1Xt3IwX+9dparJT+37PhCjozuG/ocdoKUkFLTnOnhj5qj5htLwg+QXoIf+MX
nFDVVEnVzCoLbrJ2WdDWs7T7a9qfmgTocKhmc6X6AuGbUmX8EulAOZLH2t1wc6ZFlb2DylZIMSFz
yWfcjHv8ApzohGs6boBXY6fblkD3zH/smkC6lEM2djTHOvY7sLkWbElSQRn3sZExyT8s+6ywTV2M
gzWQrG7CpQ/eeIt+lNnF2C2Xy3NazMvN6m8xO7L8nSIowRUQNCs+3SLRFC/drq6P+vshIflHrX/n
tssyoOTC0Y/HuxgaPiEV1WWi0T3DdqrB2/FX/DrQFaP4z0pAOB2Km28V1N0ibLjvLdiPCTqg3zP1
CaVWWC0k4VAIkATVUlSPc4RKhXWn6eSQfAyiU82uNj6X1RPj0s90tMnVtQB4y7w6BwIv/A1y7YQ9
iIh8soOZebyKa3bu+/ciXNjDjzmnJxd30K4CPLuJVzjrcsx7zbNUPkMpwQAzNfixvqZ5IyRtnHjc
T9n2bPMis3kay0HgvK3FAZ2RxkXW+RWuhirQ0oUV0ffMr5ibe/qUxoVUiUsjuZlZMIIIN8nTjDgV
2QV26KFvxUuRfjSPYvYmkvOAu1jUj3GcvZvIMAKHoRuEnjVScbzgPOh8ZP3nMylpffofbcBYZ2oo
H3Y59RMzW6DEFKhJ/kKP5aGhc3vc2TSrgKFK+tsBEZ7HHjiZyKeoSamnvMmGxwbBDGKJfD0Y5kvQ
loxfKy/9bcp/zbNquhqxXY4KDxVjPTJ/eAr/5ruOA/H9Exuu8MKnzgJUSVXZeuMVK4JSKi74v1JX
89H818dbQjSb66nWn76Y5pZ81PUIk07RLGilFlEVCwmHBEwACvMu3kNfm1FDTWNUrGOSI3ALbQ8p
liF9+M8bRpeGxg+A9T102BJIysFACXUsSLHXgMCNrUsA1SuPQZyRS6HytLnLBPInQ1a4u0c9z1nw
TxVF87DQr7eioD0d4vjVE2IBFNJFz/eDpBVz3EfHtYYK7gHG4ChSBuPjzfq5k2njXcyOB2GB8TER
XWQaAfQJEosPoisirsnV3TYiclNXPUHaZcADiXpce0tXl7NFSty3xzLUjTBhXh8fFPTbWMxLSPSk
AE8tasqgQPRilpf35L6rAuccBc7haTGEaXY38M6sQCGULWd8zDHLdpDP8z/Uc20Iir1xWQyMo4r+
34uKL7O3CieGIOFqcEz61o7cM3NHd6rQ+rkWj2dI1FOGMJQyaTE9UooKUVilUUiq152g+cirDfH4
3slD0u9DlY+jFRx2PsoJH1RS1CU7OL5U1unW3GPqn0qsairN2mc6bGtOEm6RjYlqJZaWDFplfnDK
laaVmo2SFeb9lsbdm65c9zi1LVodHyj0qit4KvfkZfJUYWd2FBFSfn5teC2GM+yzXDNv/D2J9key
7Y+Cl+2HsUd4ORB4SmETK1OSuXGcEmtBol2Ssa4M+56jHSNigoGF/gJuIuBH5uIcwX7OufMKaWTp
h9yrxQIf+sOSmJdG2gYfc9fHtL6lfOgwr+4ex6sJdgBCDw36dsltb3wpMlnujXjFvTDgtkBS2tOG
DryyJ86amx43Pmh/wsqxwXIkZ3JbvUL6y5DbUqgNvDL1iC8wgCxk8ZKaWxnMdt10UKGg9RSSd6Rb
+hgi5SQDRetOGEFw3eHKuXc0Aoo7Z6SroMComhp6Nlh5Gq7Si9rOxDIurcpQSaaZgG0BJ36K7mel
zujSZKe2S3nV0ECGHcFtW2YRiXH3xmE+6x6wiiXjQOAQ3CjryIrnRjp/VBL9DlnmAEQMKaSfcLyn
xU9Jy63q+bFb2R9oHIDo8yx4EpB9b29DX58kBfMAhcyn89p2vx+dlyEgHXUAgSYyV35Y9qBkQIK/
p5D2S41BFwLClC1+jKScNGj+GXaw6689Sy4UhC+DXdVciKsy2oZDKfxQqvbBL1xQtkuvW2mHh3y2
C6IQw0Uj5Io+wmN/TgikjYKsXsEZWBCKRJDHJHgqWS6fk3g5nKg7J7CV9Dqh+3oD0sJUvlFq5EK8
qTl5YFDlZGLKtvZhDPNpKWXmi3DnFbT0Fr30ypPiHeDVqMEuy4NFmHLV1g643bNgBBMEHEXK4as8
AV+qHbpuLUU6YKQTyEKAYax1GCmljbEqcSttsdWJOe9TPz+1ePlrwZhmLpSqYnbDbHDZqoErBQVd
JxVzXt7TyO6J8OZEYfjh3DsDENhCm1vcOPmR2rFApnWKP/UHzek5zvoshcLinquD3LsaC3BcKx3g
aW4g/7wW3fMgnzO9jiZHWY8LHTIPMKHh/p2cRqvfMXIhYwb5DoSw3jKOm7jlkAc9bXYda62ebCb1
gWffT9WffK+3DrKGYizFyVdamEH00sNxJ4Mbp6dmiarxdBV2RX8ZUZE2dsPeG7YKduHvok+FDPPK
r9MisNbFryO0fxKtpJORnh+C4ze+/E23tSHarKU58F3H5xlq9Ty5Bfw+VzyYDV7qk9WVs/ELXuKv
2/xkWA0KeozxeFlRcRN5XhVhaZcodbjIBfOQ3DN7GipilblXjDdEZbEajUKmsQzht0bt4mD1tlLk
tTWFi6SI87nUI1fb73tJY0ESB0iOdqpZusgoxR227RLRqY/2UXE3m/1Jeh4+nEtEXZaX45CmKpLx
K+FnpI6ebyyOYI4HI6gRRqvX9+cWK6OKYzZ1f/FRBjyXmnPjmyA8Wa1szP46iEjCgvbbWAEKkVr8
SZDm8YUp/KPZIRX62y//moKZDcsftLMAB7EpktiulPf9zS2vVxtt2vnEqeSIF5mwPOQiByFFC/vk
rDSckXb2AXOpkQwDYOEYeLRuPsY1nJEhIYqP106swQKwOrDt6JZ0FB62dvLXA7bo90MswT5Vd6RE
wQuR3D7sbcNufv7lQjrgCDjAGU4LcfSfdyhAOpBAp1c0S1OzFj8EjgheDjJRXKneg1wdwA0Zbj2R
6sOXp3HPBN03YUSzO12g2QPJMcs9LzZTYaBu8iqNiKKXQZuv4tUjdF8+NDMJNn+CHhvN6Eooa3Tn
HJFqNubn2IdJr/51z5gbJIIk/FuKsMauZ7NzTamLOdxBnaPpBiJj41vaJ0WBj3QdnwyAor9sUO/F
2F3G5xuKD8ZhwpLEpItcc3JEP3Rm6Y3kN+dXbXDtrawzpjLkh1ryJ8X19m+Qwl0mn4nBcFl6An6a
8eu87PbpzEEgN/2nLy47xDM6ObYoViD9b4nLkpaifxiDDIi0kLjmsNLjYTKUQimy/+yD1zMefjKq
KJAAwuJEbT5VbEQDOer6RFfrqU58jjzoSCG/qkBWUxi41GBVs+OafHMBA9pG6u1qeEtozyJLCFYV
wtysadKH8pnqYIKFN2Novb5P63JrITfNgV6rlLVFjwJUCGyunQjyG4LaYBUwax9moIzUI5/LQOUV
n+s+tIovcAMlFLF/SHqeHEKTb4QgG/aAsLi69OUJwCnTP3UArQtCsZAfCR3J3Sq9cly5u3hGJwIy
cI/5NoPSvjuc6m81ufWKbOZ55WRNd67928cE9yZyQVX49SsYSINa6NnKt6HKc4Qt57CXLcNQOLKi
8kYQLOuwJNOIazbzmdE348z9Vg1xlCpDQ4/S6nEjZFri0bAe2Ov0+hlDSfbXBntTRHDOvgVrkbpW
baHSq4ZpvOgwQzys/Rc5stAbGLPFQU4UQ1HXX+RIz18cEkvLbbv7rqWESQGrIqwaVjvqKrI6pZpq
D4LratUsVyAPDoh1TZOOlmUCBkoya+ZnvRsrzeeSDAFvR0CPXE5AmfuDuE70xpeje5Kox92HExpe
ojirTwmG4Av7NUnXJ+kZeITZGmYL3dCsS1UtCrxk+CFy7ILxmnKHPAAeXIrkNoKwJNSMwkQVs+OL
NibRVezZX59IE1EU2Wr78HDy11AVRpPIEL5CIWKFg3txWtGwkPcIgCMeaOZjA3zmEarw53PNOCWo
7NICZBXSp1FCGs+bxa1UuVt0Jxso3HImkqovlXx42flVvYahXUtjyjXPXXRb2cRD9W7pVOtURJ3E
fWG6BJbTTY9r2ZjX9WNlgg8+ZlEBZcLXwcqTY63uYQEKuTfyCmkzMITvUgO/65CEpRCZgeYWpY8B
CTDYNXY6Xfmg/YA3mr/0wnt6owHTMjZsy8GI5Y2nCyp+kHNiHRDHrnbGnfYGliHIpO66a3eA10Vn
GnQqgM6RvVSfyJde2I6tB/Q7tPjEt7OtaFLJyzNoboQKdTVeLTYt+r6kSnczJFJutSwOfhjGmtp2
F3LrN5AwBtm8hXeJp4O6cLLBufbTsJ2pzmV0Z9TempQ7tReqAK4pliESbJ1hfAGOEG6AurFLJlcH
RfGKe4RlBwQ29BUnilJjhiAu2C3C9MghSqVhH76n4eWjrQQSr5A6eouuA0QSn0xZpxmj/9A6dsKb
QjqER6nONdXbBlO+quy/JsD6QjymcuPimE+5XXAAzrOuFeBD5PVfzkTz6qdX1i/XcFcKNNq8xgcJ
uAdVTwkcAedn1bUmJgLWhA1a2c1/Ou/EkohYOx9AykKvc7njriLsv07SO/4V8Fv7xdO+rFP6JXPk
ozAHbKrKWXLNB+bRTKNGp0WKGouzsH3J1Jfkbi/cRM++7+2MwxN3FQGGDl3ynYvH8xWGgROmVBpe
MmT5UMO5Vr0BUuIM143o0LLMS4mnmeD+9t8b4wprOXpw+rGjK1AB8Qk3HZNVQXXZUjOp3fhXeeN2
PoO4WHzVcxmer1uUcVNdao8CbjejByL4JE0YaqnL7EaCZRukOhkL2sCY4t8F6fg4vz+T360lp8rO
ocFXQVKCtXZ8MZ3Y/BqS7lrbYRhvlFpz3g7TzK4W5z/ahh4jnL/bU6RFutCqHP9KqWhgrP6olxAM
Go7pY061+KtYm5/1IXAzpQLaGq7Dt1cTJxebQB2P5LdMRKY926OPwgwSG2sEqravgeVPUePvGtU0
zXGUFoE3IHbTztEd0Wq6AwE+3bCs6nGa/Sx8R6zD0XfvObT4YREJirAygdC5cmJV6VIl8CrciQ00
8KnB3A148Ni5FG3zEeU39uIdrE09fEG1rJB7PD/uPRR5vzWrHscpDgJsCCxdLnpwO4zveQFv32ZB
rtAgWrgVb20UjMK2wqjfWtxaD6GZ0rFQbKZvrmWNqm6pyNmhm1uUuWp07fEkJKfZSC+dw4hF3i+x
vW2l+FY3WmCLkk48+OFJhvIeJUbG0I8NiEuCUeYbA74g5MZj6nOo+XzGTp7ErBjIr7Ft7Jc6wAdr
8MYz72jLPlyovVmaxNzHQCs3vlaQtNunm8DFkPazENEq8vHVz7Pw242fyrX7n5MBQLqfqqA988/v
MVjakpKKEONpJcFktHBIU6Cp4rdpBgXNaz1FyC+LuhJKEFmMIidEOTxUCjn33/W++qoFf0kgfiR1
XWavOkEDqFi2j3wJBAIP75WczsXnh9r0oVk9sDC3RZfj+QJnYe2DhmfqPoL1m+NfnntQQets2b3l
pTZ5kP6FAfpQTfxPRrFN1dJ4z0ysWjDrBC1PAMIzclAnD6eAFXI9RuM/4v9i/I71ucgHcBijausd
/GyvjvZyg9eIDo44um48S+P9jHoLWr361rVXQPGF1cXG3fd20ihFpAdhaYsnIxXKth/mj3tev+G8
mlfjlpTt2qFKCIACHagrUIRbHbTHIgkS7+n8r2TvSkrmkUeHG9/pCdJSXJY6W6BPnx9GMbUZcBNb
OpeaTakiFL/PMVa7p4CmzXNFR2EuZtx4ft373K29NQs7KCKVYoqtTZlTB5YHuxUBWUfLefhdTALs
1OrQ6I663ElkF2XaF2OJ5FyBZiD8wzJVPxSY+fD64JdMjnCSu1ne7agTEkeW42PymaRQJ5pJemxa
nQJtrWCov1y0bD5pxKLhBSo+MvbLuR/iUV9rqHDuy2CRdNC6iObbYuLxnuiCuCtB+kK3Qanul0Cu
Eoe4Sf/iVxwK2NAHY4Y4MKvxcxWvVAm2sAo0NTZRccK/K4YXc62tfPCzNqWO/xei+eF0lcicGAUi
WdiUrwq4Ujxo3TN0vr56ayQXcl1J8MBgW8ngCVGPliNApsZ/3hFTRfJeXgq22EmZwQmJJzN1qTxd
u0epn3zgw24LgwMVZqxpHkyqTIXsJ7HyhAefr+gvIJzN4EHKujJG0wy7EheBLUOqro4MFelsU80d
ZJVSCTSv+lwFHEqqUh4fwqmvKqV3OHItXgXH2ZTqMQA10iUWABJR3Jtst60a1+3EFUCf7y2IP0Ni
W816cvwZoBkhuM6HYiOQ14NhhziXTLgSe1j3suKv3GILQeLCxSXHvEqYtsdADjh/Ph2TbdTZ7OvE
uyssYcaS2MJOtw6qf8CxlR1B2hVg8jBfavfBOOKHpjwin9LkR+PtMqJNAnMLLF2eQmClHwVovosA
gU4EWB+wy56S08+JyJcd74SbU4Gf8YrLzboVMCZOsLyyJsgkPts0wiPkFWkeCaC+/otvtBTApGG9
r+p+L9A1hE1IOZK63B+8v8bdQJlOpb/KvfyHh3zYslY5fx5RGkAVCr7KGWE82BA/SouuDav/JOzX
ac9bPDTemnRm4vgITsuSLvmAD688WEOzn80CzZCzHe4YjKgv+XS+NI7xoSS7aw1arlgccC+XjbG8
0rt2tvT32ARRwwhVFQZrTW/+tFBLN5rycJLZH3Iocf2nBJ/RTRMKO5DEkkBFewmLFYM3RvHjbDrc
d5yXgEFiHBcJk5wfgX/H842Etv1dhcmwzgyT2Q6bg6SF3qXLPibigGHzRbiSPNnGSUyuwMn5nJ+g
SpEahZjI6XpLj9V3gZ7qqfgzgibhuKfOfW17tfvT5CSR0tG60B9sNtZJVDWClAajlC1mBrg/RQV8
Lj473mJgMCki6hjy7PmOAgUG6T9I3QZ5D2VZQJLogI9ciMXR5qj07On4wTLvSTy71sqqSMevHeCN
YMyfNV2OQEGgiO3+4nNj7+pFalt9olBwRgMDyfbQ7H2QxAd25bHZUlxmA4cxYNCxFm6PE2LfmrJp
DlGpK9iKO/xYh9oEcNA8NavtCJ7BLH2Hc+lhiu6ORPNtw1HruffZRi90zUUHLJst2sQ25yRM3C5B
1+u4gRyiTHhK8wEYBy80+J/N3LxbLzokF6FoZ4ieKv5CYojfN4VTDdGlcXW2OqctZtBkPn0p16b5
4UXLjQ2KehAdVzeNUZaDUaCZarOmXIxfeVwiaenqR8FuQo+KZp3vGvtHRXVROpXoJ91fKyrPbdxo
WCMQYssTQ7pKRp0JX35vUhgmJWH8o1Dr07JEm4A02Tnj01camROY6/+oKruhb6sQ/gDVNUNkGPfz
ZAvlmQKGm9gR8LyjCczPoiCz0wWRcn1d8BzwthrZuJbVaAhQVtdow6ZrvseHrRONV37vt2fkOv8r
F/C+VkcEQarmYhxPTuHc8fyS0fqrA1JTlBSXRJkFNV37nJAvk6+/SDuAf/eYHB3dMC/A8cfVYrJQ
VZBUk94jiZ6BSjYS1MOl/uixeyqHUmZBlvMbbanZ9kWCdCX8kj/E0cb9i0DlB5aAY+/LP1DrLAU4
uuf441tGnFyGknxXnbCdAFShGhJ1Jqm1FduqMf2vKeIRS5/hcFukxAohRH01iUEtbOgQJzEZ0WJ6
mh7GDcfVVtHnAx3j+Or35hlOlalbHWysSvdMFFj5j5awyOp5jVS3PhKLP4QtnQdeJ5OV8NSpEC+X
xmBHjOfCRCw52rECxAOMvEyr5Ke1EumpIfXVajQNCJ/A9IJAe+Xxnps7FYgKFsh6ZbQbYD5wu9PJ
jeOR6yVrRwJzAj1Nt6wqURjr3uuT+W/d0+rVVgJaiIj0ML9zlsR1XU2UbITXUCyAXOMPCOFmfl9/
GHxC2ue7ELkDCzZJ+YwbMI2qb0Hc3XIYL7GnTKz5gMvLaiBSIC/7rsEbLyflwE+nSt3ELqs5X9xN
9FTSsFCjiOlEbo7WlXH3qhZsX116/rG7t8EaZEp386NJeUhJwUZm5jnghd/rSnImeBlw3Jm28IBz
ScDdlgPO5jxzJZThx2SYhECnI/W+qiZzdxLnCI4U8K0/VfCWpmeoEvcBLqK53yvUwN2wzAvWJxTz
WMdqoycH0yMAjSbmlYA2TXxiwx/iCVxtWj8L6z6qn74OzFzn6cNtyeBLiYgIfdF0cZbf4tNra6Gu
yMRKxW3jud78wgbbJ2am3PowhDXBgpsy//vOlLCG4uE1pl+ZdDfzXH19EbJIiB364kaJqZ1Gy58x
ezGHJ4vkBxJFV9oys2N+f7Ieq660GnqRsNdh4tEXZ9G4kdPtJLfQAhmfMzcOCh6hXgrpCMiCU1kK
AlaSgotKi5CStKbgrOuVwVL2u0PJEBxg1PXfz7sQUlziKKW7Dzqffg15cV5uaI4PmAs2EKYV7f8N
Df9IfE6F+rcOe/7z3cunhwCAtERWehvrOYBzaxuOQHsjPcNd2Gj6C1Fc272aGn/fkEkf/p17pDwa
lJVH7uhW77WjTvNEO8UPPC8/30+pTunkppCI10cTwpMuNnE8cVx/yr5WJI9u1SY31m+uu4ngCO+q
2DMopc47AsUlYsAS1JD/BNfaRsBbgf1xJTEz0GrWi6XgJ/AeaA0tkkLTNfF5k5OppglyRduA3aXt
gZzOhKkN8IzdDj+c6klFaVpviRvHlSHOi/Y9ugKuL/RdQ4OZAPceY37wzTIaKMo8pvT4OpkvTyyp
swW2aeg876p9P23ShiMu11C5oOqofkpH3YJyh7G/MuZ7FaEGC60UtEhqOhr/jgid0NKX+7u0Pkzl
++z1Smg7xAEq9muRfDk7DPvLv+30oVlqzqh3i86Gfb7lyp6coAarsJgwy8qoXZmYkC5jZXLqubLl
7DgJ451eqR+6zl7yD4xVXfZyOwTCsc6w8nEgevi2bp4QxqQ93X/0wJylZXPwml/R3mqVYMkVFBG4
USrdgs6Nwgh7Xf4oi+ArLQTOb+/RTxduXzbS2ND7itK6WHlCq1hydD5ymYWFG9p4lcTZJ68iGJUk
v5Ump/HLEI1hOaN091tXU4LwzktmdNucTao8L6gcUME6Xlu+V1utTB3A8XKJTMSZvsI8Mo+fiPR7
lp0LhCWDwniVj44FimV6EK8P2o2X3KlNy83pUxZeq85yHt2LWAfwWp2oAymQsWRAZ9YdiapM4W4O
x0PXLN7KbAvXY9SMXhHN1SDeUufkEu1a+wUYQ+oQ8gjz5aaSGitCH/+VGYZkUlTk5sKSL70KrZ0I
RTdr9GVtlE/PGlh7VDCBYiRtLWnnfHTnbWOXJ1SW0/Xx2z0ECi6ZyFeSkRWuk7tgBavRU1PGdYFe
cH8v+5KYVRKY6ynNCsmy/Wxhv51h6g/3naWSAnZbHtZK0S4oOfmrfBYx0/29fHMpPUqyswulZCmI
8pxOTu86m5PhpOoBR3wJSmgoQavuxSJc+FDAeeuX/nhC2aWl88WOeAR6PXsD0xDrcZ2ck3xdePDf
vFKd5dVRu8nenxmUT3ZYswsnd/n59pl2U+bmIws1Cohz2de64oH8Ho1Th6zaSjGJtl+3jxLUa6XW
wVNFZ0LlSi0Q05ATOQZ2lag+gDcE+vUim2B/J2JywEXn4INX1SAb9G6cERYmz1jHBZixYzs7msVs
D/7KEjUcxO4fYW0OMwE9Bori3T7jQGoqyKBw8t1CRlftnKwbgPkkTSyoLsuPt2/+//wdWarYZL8Z
M4jDhw6EB64NZCwKQ1CnJL6d5SpkrPU12nRCiMrVp87mIgZ5WbdKB37qeuJYOqVQQ/QR+vJfL4cg
atejJZ4k/7RKTLAxCojkdm1vIgwAzwSvRwiyxmhtCXd9nD9Jqmr5xN6BWQsc8qK+OQzP9UPH5dST
AHNz0F4C43535PAmm7lU2tdcCYj+Fyvf1oKlQr2UY+yIS+cLIBd6jEkrMTPgy60iioUD+cG3KWQ6
LSjERsxShUjzDZK1+bFMCpaAk3E3CR7O6dxqer9YS87gl2f1ipou6B6Ev57JnBFo9A3iNnATRV5v
8VWnCL3fibN23BV+LW3dH4yi+vd+2w+NhEsTlmPgELbrDcBv3NJ9LiI6kgcmQHHjqhDMqClbr+o9
dt+Vrxf7dBx6RzNDCm01p/6imKq4yO35HJ9eGxCXGjtNffLc4XgmnRW2TT5av24wkXY3Lvlvrzot
bZ/LkCdoeQdo2jzmZdwMkSOdT4RR1wV4Ao213dvLFYqBjbYAIZA3YChVet5Z1ESt7VGwBqE8ALEU
uQEjcGVYETeJXyvfmqwuMtZQBQkj3UdHMf93IKc3F7TNlQBoUuB/+gEJDrn3snZbbQzkSNxpkdAe
YOGEQWyLOUUv7rGSp6wsBgsMoFXu4WZNti67V/nzfoURn/nUDXVVE+3KnH88QWT0L01STi8GJbqN
p7ON5ah6gVrQYvg5CYxpWQCeWHyc8l16EVzcV40VGYK3Be0ldk8BZ+YlT9PUrqDkN3511bp46emf
sKmEhFEsbCbTjRAzQSvht4SoVqr7/qxxfrfr6QqR1/GfgCfP6oCNHtUbl9a1ecy+HgUvz5/d9IJw
Pu3RfMfExQve1wQvtrsm4wt+aW8Vh4JRYOM4mfIIjH92wTO8GK3oSYMHr510lcL0xI4Z+hfoItbF
Objdz1vFx3gDE4rZP+t0IBeb5uiUIsR4oekv3S/BgMw3z+Tp4z6bS3RDRoWaG81UKIWLUjW8J/1o
V59GVITAANbrnewxRhcS8xpEQ6Tuw44pmLJB+OKlUKjcXAU0ZxRa5XE5mUAvHDOnmSofO9VbSG08
Xeebwy/ZC4yycckgNo97VBIx6BCazxFxVPKv/dgCcX98mub5F9BSC2pVEX+OJM2crgsLCE2nba2i
3OeByxi5l2VCA1tkTHnNFo+y1/cvy14bKbjGr38SjRKcuzmcWhjcyssfJaEI8MiHWJt9l/7AWbLj
5BTcIkIe5A+6O7MAsM7f9/dlznBE3PaYIwdLUehHXmggxGQ7PXfu5vILpijVQ9gfFlFywFz5M6BW
PEwQgfQ79D1zmMTBAhJM8KWCWlzckyJsM23UNAee8UgppjSJbDOQy1LDVsQZSALXnjn6Ke4BXU1y
DqMAGdk2M+yuKfMeO9VRfbzmBe+nZZbfsROn5WuGsgHAh8bRvGLwNfEZ/NUBPww422a4Wzp/Znvx
4Pfz1bUof4xUJJgLIHVOQuG41CLRUuaLKGdUHMChieLQDu5EnEiTVzEuHgCRYS2iounblkO/UwL+
W6Lf9/Vs8ZOX/pb8YoceRb7tY0gVTU2n8qdO30VsfvXyIdEWmdalV7GdqdTHf4r6TkXEDyQUgJFx
VDeUMRd7WGuhOAs38LOducjxMlQls5ptF1yeCwY/krAc+Dj/L0axHXLpOJOcbHAAzv8lCn+pMwND
7Dhy0PGrCPb9/pEQCNJVbHumM/mgVLV5OCCZn+4YW2UhGotEfjs843gtEGVAJLp+j0WP4lZciJrx
GwWOCHXR6TOZq839QW1agCJpG7OkNKveJQmJGHy0nn/Inh/5tkLuEL1+8EdjXlkAmuvN2MVa07SR
E+W9Aj3iedZOkwNgrOlwtZEYNxP8bQtD78PEmxPu4xIREsD/6E57lKmo8s5xgSu0yCoUHSw9hdqL
+LFtElaDRHyPOMmRPxBqRaoEKMVmGqPH+SMglUudycxTuH13zSTyAz8qgMsYGbjr9sYjagsDiOuY
+QrUSYpKdxnm+S6JsgkdGx/ZA5VZ5slCXe3PAz9XyqARAgXWqV8lXmBL7/BpW7FRfUpkXPov2dcb
rk9mw12uF+s0Mbb1XFkuk77cvJPdWv0sNydNmJ86j+wy7Q+SefyYWfTIrR5qvecj4268ye0JNMhV
/PDyw7Q8JbfN9U9Sjui2wAhwlA+kPIkx6zvQjiF7uXEEgOtcpXt8DS2j/Bl1gMbmWQDipkld//xH
GvDKUSOjd++Jti7FRpY+J5CLizraHZB5eeMMEIvJh+ZEiCy8cCXJFaTHfjkm8JZO/OL7KC6MntTD
LYCoawa2Ya9ZyWk+JagKYKPd86IE2G11mVQd/RqrswtX/1OKRTsUtspn93Owyc4UGxjy3X2h3GkF
xoRY+blGqavHetBGj/qTyh+HMzPsuWegLmuX4kLjAh4gNSC7WtDQXp8o8PzF6sh/DJw6gWNWXXJU
s/OWyha6/Pq2UjPal7Vgyz0DcOdtwHBRjRaWA7Ees990JTx2dKFU3oCoR6SZqtrlLUxb+VSTyOE5
4W2tBpX2sHYoWXweYSGN/+9Ym3a0fzpf/5RAL9zq530NsY162A/zqgPq54cTQgvrINdXiS7IxkIF
olNSVP0DEluMaIDVhMrcGs4ZDo0FqKnjalLHgRtQt/8UYlPf4wMyREUgj3nSl5+AI2TWm6paJIX3
LzzIy6tr8KVDB2CwQ+XPCBxNFUY2Si/1kgYVyo3QiAqTUKDLCvXX+Shvlt+78EjgQNdVpQWW7Q7A
mJHZxLj6niTYJZh77d/op6mOjyRkEIf50RtLHdKAk4XsUBR8csKIF+zVwG/HcRmpfXNiMZtutxCu
ZJ+6m/wtvwCRmty9P9d3s9SsO4HRkrGKiSnpZN1ubNMosq2fyjUytmv/h47YhtboVRXdePthl+M+
YuMiH7f+SOgC2IYUyu5idSnxJ3/DcgofvvkE7+GfEgnkmGDhpWDafRBFLo3zaJcrMhzKG39hm3J8
jzlv13me7O5baqop+uNW+xwVFgprFdm3en1bxogCiCU6AYqkMX4gX6EwjvObZmTVGXO+GtBQNGp7
rEKmeCc64/BOGTgleCjxdjBII8Tl25HpZ93fwIhgc2O2FnOdeFIwhr7wDPMwUQgYewXVzrniLLva
JIdCV7gpY62QSOMQ4Gsb6RKmI8S9VHK7WvVAfFxk06yqmlDIdetMVTPCG+aTGKA+XYML/rIStHry
USBoEjVjzJ37WP932b6t8sXihBO7FOk68hon+1KGAy74OxrxoUme28sT1AHQKQxLjntaYIJZo+ys
Oa7S3KjlqAO0cq7sUaOUz++lcwGY9Z/riFhjWio4LR5Ea2cvoE9W5++ZtUWwbil8QwUK8IJI1WF6
u5xipSnvICY14bdgs0Xx3v1sF/GOzL9z2i28iJdYzgTn/EDQEQjOBZVKjqWQR2T2EfKH/PoLsTDQ
2gZ6Kl2dG5ykpH0LHqivIIhY5eqk7nTdB1+2hq097xmZduMinQnbW9U2a1MQnpKV9kjoX0gVpCsi
IKpnF/XU0ZbNGGuPljzXqu563PpYdwQLc7NYJW9FLcz8AMmNJR0Zb5/YHoot1rwojrhd9Ysd/i9D
Z3B19h23BYPiqZsRCkW7IdVlnOwCxZk/4MRCj6kHtKALXvv5fZsms4/7D4gSu3ctp/tLSQ1tiHe/
TPRgbDhUkNXGVsUVIFEKn83+iUEOEJDqaoVlCU54ySGV+HTM3iRKXNf1EZdjO8OcVh2MB6Zm8zXf
OKYHpjLmf3hJ83DvGXwZ7s08bYigtW3B8eilawwNEy1xKXCVPbJxUkUcxZbZxK6nSNAbEJxnkA0c
S5QNyiAotUpUp/bk4DSvYwik89sgXFW0xHER2moH1p99Hu2MkyslpVewlPAfDQItaSlVE8+dbkIB
BjAmVJ4LpDp3KTxOR5TfgIwUkjnAE14bkjDkwd6fCiCIoJTHP+Z849vCRD4QoIGfexVXFXeGrJQ/
uWwmgZhAi6W7nrym0hha1JCXmFJdB27Uixlvn3tBJW61FOprr3aBtwZMo+qS0NoHmo+NXH1mrdUc
336hV+lwKEjYaBz+xOSR0n4Sb/KCGFtGGqR3PDitGk7JQNh/SX3m+tga0mDt7qu0ZOFnDcoW/BWP
qXC2jYlAXulERD+aeKYDDVSlx7+3UHkn1nLmFr6i0XvT90lMq2vLls5BsqGP3MAUVyxorb6ucLXJ
yTjEtZVJ/MeIU+eqcSTTlz9psFPw3BSDfAgchlv671ad1xxVJiZJ9Yz0FJHjt0eR5c/pUTZI6uoc
TfR4sXQLs+P3qxqqA1Caq8jVVOVm4McIwkhjuh+oN9RXUQdZsD3NTLvEbrjH5u9U76t3yfj6GxWK
QWQcDyeLh4EqJsuutkEGcvY5L5Mk/xPMahYhCW7OYwsI6rD/IDLsTIndomVboUop0OD+UAncB9MR
rU7Ex91hRHYdCHiER+lA/qlhnhKcm45zrePsbf93BLhMUyQHdFMaPvmxqhrHpvIvG1U0iLEx46Kv
Jj4RT2ZFQ1+W8OZSS/YZ/HrX3WAQ7cInYBE7RHIGLRHH8WxNnwELlMvKfdFABR+EexEthFBK3isq
a9keuS7w2k8++grb/1awjmt9pgmBYf/qR/J4eIW6N62mcjpdSNwGqnXdrJxFcCAPHu8D9+1rn4HC
sCd3uz3AgOXbZvI/7Ouxk0SNJh2lk4Is5RQHYOFnYKVCsfaDZXkQmEixQNHLn/IKqGPv7MNHDn0Q
wnQAwupTOqxopWuhF0IP8r00euCeDobtt8aow8Ss0AeS6fQgb762kbRmgZk2rrV2cxsIRskkLI3A
7N7dQUn7+JC12HspnfaAJCCUs04cRfyJZ4jJXFRu4PKL4fdDE2l3DZ3CT8ZTeTQypEVJfCv7hnkq
GhogTqOCGeJ9bBQFIR5PDpqSBiQA1TLU8rW5hd2B3FdzN5ig/YgGLpX8bwYf9EyY7wcz3PCflpfL
9T70eP/yqDSMpX5os6alUyVH8OTAj0dFoaExadHsz5wkz98gDBKtoGCIIum9H8XBTAk/ytb81u9V
GiuT9QLHEr6CJH8i5Fgl3nrdn66WfQZLjd7zS4Fxg9brP1nVQlv4lb9E5hYx+V4UogQ9n0XZkMI/
PWBDTN8SMqpt0IU44cZsBYWvHLoMekZEKn/XoqQQ1RweuXnjl8NV4+DVAPy/fzFx1A2p9l5oQ2es
VmVLd20W2wTrChrIU8qUfbKlRLb7+FKQBfkLjm//NXuzUXQ5HWp8K/bzJ5eDkMVQXFUVonfvhftK
AIGBfIGu64FMv9ufianjYoDeU7WmhWEfAD/jW4Uf2JfPqD8vKByRM6C2jtVPpVSOGpGyCSFnXgsF
j4hbmszGujI1L2/2bCaxtoOjE8sMTnSQQbmK1InW4MyAK566q+l7OnNOfD5xWXK4Y21s9AgOHEsF
DS6g6LdKOVhBV2K3+f/yWD/PLSYQRoSCNpo1JcD1pcXCFiK1+kd0SCGc/GluPVH5z+Hu53byTzuS
I8+yzbUuubDfrFeqiuwH93o6tPuva62BB9cD5bMWRviOT9NVFcQr+ILsEiasRVdFc8EocOGXgzvb
R6Sp7WLP+V67HmGWaAWrwREBGQ05JYrRxhGDS7il4k0FWSQ/2yVXnRayW/ofHusO/uv27bI9547n
bz0Cjz80vfRWXLpwRAd7Yrz/ZQhLXlnFMrl2OkezIZD0D94sLj1TjQ8o3jHr4WFa+04C1gn989WF
4vDW9Fu8WrjEdnXboRaw9GX7RHY2qorhmKORMV9RU8ikZVmvJZ4dGM95YpVTPbZYWvYJaAzhKNTK
6Rl/+9ozv2HfPL8/iR41HsQNpYyoS2vVpNuy0yfoj229VCupc6eS8gX8MoGuxsbOEiSQncE4X8SL
vidxuGQPYjv9J86h6XZq9dUx/xjo/GrOPfWgwmW6HQh69oGHawkOMEFCWP01G1/yqzqCvl8otK3t
5sEoUt5ms5qZlu70B56tPQSNefZtY7mDSxdONNh45hBBQ6PJIwKDbFr4gvuivD8aPPdddKT7CTO0
M/EQ2fWOGDlAYnGFbuJ2LRWd49Zmn/0G3QHm7bAdS6HncUMBCvHQRqGCm/OBjDBvgUNDE3t3l8Bh
ehJoxnFanm//LY4VJT/fbw3ehomYBeUpBfEe7f2osHvE+tqBKPsKuOyz75+8tKpJSDqO7vt4D1mn
XT8dwepluekW9/STukxTPBp+DvRubRqmh+JDPR3ofSNJfnFycWR4YK8Zw/0oEUg+sDRWgIkS1ruL
W+xQdCoCuGSQFN/m0Q1BqqvI21U9i0Dy1ppbFIBprkqwLQAAYuJRMcx3z+DcolOd2GTIB4HeX9Ob
7r5SXzau3q3gokleef7o8C0lcfwLOeujJ6B9wKJBy2WAakJ8LLLaLy1pN9JoS2uhaCUelI8dUMO/
B93GKV5zK/4RcWtz53uI+g6JqfmPlmJsPrvG4GwLExbKHAY/lUrhlfGX2tCJzt/2ZxJ0UCGm6xdY
rMsSo0p0BSCzUsFMSmPRnhnVpfyzEuKtvWellr8XOskLVVaoU8t6YrsBRfFLjWJe304flnE7PXLg
1/GpmaGgbgfXbtZXh4G5yfk7ZQw80dk5p+H5jQx6Ubiqi7ni6NpnRWdS2EStV9MV/W0m6NCPFxSy
Evn9MPyWVxhUvGTP95nLsPMiY/3ECXjunIX9m7Ggrdj3HtC3mjdBJV4ZmZiyhWDhDjvjFKdKU85l
8GHCiBNcnbAaSlU6Ng5dimLNc0u1l/dAxY71mahppHDcSB+yppdaAO2n1SG4bLfimb0P44+iRvM5
Qx86EiAjD0AP0G/u2mdqSX9PizapEp39IV07aH5SN19EH7CfqyJL+3MaJ5xcJHtqOywTYIxTIu5o
ZxtiX102545IovwfemVKgt7gzDbJbTl+jmFJaPnQYK+MfIRXjqbL1IRkygJ6z2bSYzj2rJ6ug/ZB
9EvHB8MrViLEVA00io08/ChUviZ3a/eCWY0n/OfZQ4rEXto8ZVRowyJUCYtKP4yEjD5PWctP5p9r
hCJw3Rz+a860vorj6qDqSRvufXK+B93TJNjRligS0eoEpywZ3KWn0X0PGX7uIQ3uGWmzQ7nlYrGD
j7E9eylQv60PXwwei9Tt5YKkl5oVK8SCWeuurAeLA0GdhtimtOOhee280r+/GH602BpVGGneT79d
nhx2d8/KaQ7ZQ5QTZiumv38N4iaYj/rFSV5a9EB9SYwkOy9Fs2F+U+yQqCeRwZS84f/ZisXjMm03
Z2PumuoiXTO1nGdQDOGzQo1STGwDT2kUVEGTAvQymgfQD6B/s0jaEkfXKbuV/L8g8pfGbyQvaq+2
a/Kx6vUTTxZ3y4O7Ed+ajN03jXlofSC0OhWjJ3yG1k8/kD0V1J4224QO69GNYvHHtR2s0iemwavv
e2imlmxZlcI89LSEMe1PmnZ0fRxTsMbS74dwXo9SoHhG23M18S8tM7mX/TD8/Oc660JgI4sWV7Gg
LrVJUEWY+TjO1kQhucEGxUBMFamrUfKGqK7LklWG4g4c12/kh7lVar7Jb4Q0OkvvHpIG9k1e1igO
2UxO3njj2MU5sQ35ECYXQgBx++hlGLlmWQkEh+0ODFiGp8/pdbXM4wi+62FKALqWLugZ8bw35Hrv
bQ5/7JWNURrtWQD2j3aG82yE6CNs9r90snYB41Z9w09WhXbi9iTO4DdTp9vagN+ctfkQc7a2KezK
ycsvdvUDN3QrD+7jcRDEJ5uT6lRjtnFWGsovmirDJew/iFYdWp012mG9yLF6tECuge9tJLUKkBER
sZxL1KEWyGNrXKZBfGV4Oczf+A201ErzDXJyeduUgq5XBaP3qsaK++ummrPFtv1JIOTYoVGgzzeM
exRDXSKODyjStMs1VJlR1wZ5iu7lwuZRT9sEsKclkJdn4c4HIPDqeVqf0Ci1aJ1PWiDrgD3SZWDs
LujvnJH7uUnXl1OGm1zN9/iw7jGXn57IAKaThnpBfTqtqUWMpiv3JFZBQfrNSlcpDoez+TWWsZZh
CmCIzGj9x0L+fJsZrGFid38Rf0ZYavcLaxAIVPajQm4W0GgiaNsZnhkc2JzPQ/NX4wi2RF0WGATP
8Ozb0wXy18sMwQzD5jaszmfxhWns51p6yvOmJ9DkOs49/cfvsCDNRifzhCyIF9yKqKQtjAnoWXZg
ynEMbKBSFq/2p7BFtIG+fORaGzlZJwaUOM1gBMMXsZGkAqMEpH/IA5KXeiLgywpnRebMIk4Rosir
xf4RfTPPq56q816q9XXqy7+lXhN3ztNAhJUVoLWpyNT6BOb4unXVjjyeSJ/aG2SFSGDaG2KhFEmp
sPgGrOg2TahlQcFFfrCu8ebmiJpJZnosa85NBO52xvU2dUFMRKazAGTtKuN8oeqeJx5hwX3gJdpc
KXc4WP7umdEVVwapo4DGmO9ahwwoFlz7b8UKnWO4Fpzdn5aE9rhKbi8GlGMZ7U+OIBHE/oQ9LXyP
VYDOvTViiYDK8r07JF5S2loudmjNSXFxBZQkSAuJbQNpX2th1Ig9GylE+uc1WW33pIcLC7epqsLM
fjAwi1DgAs11/z3ofIWKne3Utcm2Pxyx+wLjYcZVDIUYrkME1yG6Ij+p/8/SHqP9XXbd2Qn1I5qC
d8AjcZmsNpp7p2b8juL4+mDGFoyrFXG28r/8bcZFVrPxmuQBzJGPInV4LfQmpp4TJcOR43xMq9lO
9G6HdVRvJ+sDltIXx8/k6wQLxPxjY+S/dGZVgThhThtxYdZobZAa988/GUxD7cShkQWg61q758wi
h3vfpWlt/PH9hN7Lk+uZOFkv4y1yYDFha7gwGr0OQk7kRnAuvxoC5B1A2UT9NHdME8azo3xOULls
50gShXAM1Cpfj8Lyr2EtgvZ+QlDua3NXIzN/9fjBInBtrI/nMAsKwzAuSxLIYFp4SxY6+I53AzaI
FE/CPw7/h3dRB78PYQUFAUGPAYHF0qxNtE5XcGvfrrpEGU16YmCjGcp6+fojZ/ruFmZCmch0hNIX
kr9qPmEn6HBnN+JsYxkow1Xbx9ieZJ4fYASenVKXn6ZjmZhJR0LhL1/eTo/SijYQdihoiPCv/G33
ROuOGrQpE0SHKvsBwzS0XQqMWLT9LyVcr6B55RsE6Ub01LUZOTHtDl8wkZ/s1jYDy5naat9YxhGV
7QXyGyuLumNS0kdS/PxrwbpB88oxhxoHKAV351H7R1Wg0qoCkPv/0ZTQzimBTuYUNWrNF9PXFoU7
DM8//URbEb5nGtJ2w17J+pTaVzBUykRwSubcuH7VSxdlvHVxItMcUj77UMdkcpGwNYUiQnTaJSpD
b+crugDp856r5016Q0+r9DfImxSR0+ipXE5jf1lQauG/fAXAz6NwucvivpP8WjiWnormH+g8y/Zb
vPgTZGkeCax6D8mpAG5CTRqk4wpG8lYum6IS0w6eP97ovuU29DF9fFPU7To/Hyrw2Pmzi2fmgycr
77pdC+Gc7QmkfX4RVTrU0b/IUmJsN0nAxjomKrvYKIThf4De8eCImCind9XWVsR8jpN4Hk8Whilk
MKqCBuL2sLewhXoPQbl0PRKydxUi9LQwcMP4QqmgmfF5tIniP1lWBE9fMYnk/DsqpTY5ryS9nprR
5oYBrflc0A3CGw7VDQlZUTdhDAtXpJIp6iXg70mf0gogh/WRv4p4wZdKkknJ9y4Y8QuwCepEvvtr
hE4rrTjfaXX10kMCMoYkBZ0QQIHCw81foka5p4Lli9SlENdUzgWywDOm3iKskksZBnPyziIkv5id
7thp022rDGTFRG5EL+ILdFjCyXfWdmoEZLlguyTj88A9TVHbDDWsCDmg/f+5JE1ukIhlAD1RBP8A
D8lZBV4Zb5rrNrOow9Ixb1c7fH4nraY6vHEiqEY9QLM48vFuRbiO5j199qz3g3suEs/6uSldNuoJ
A56wl9Rk60PC56FbdRWFMy92L3++7aucSGnU9xBSMU9KN0AWqbqtmOSymydHGGYjOPk3xv+E3QqK
9fRzD2YqqDb86evJQJkUIUipQX9Wm95fDSVPwgn3eFfUbagqNB8A0sPZ7LpfpZQeaOOpgkg5VMwN
KmcAsk+WLIN+0R3wmV9ZEtURpyMgrQTovCm9NkkfNHFZ4Nh1SQkZJnq2vbGMDsDZDF0v2CKqsr1E
IOxZhwyNVD9JABxlyUPTH7NmrPvJtq+/a6w+fz+nWQz2HZArv4dUPTryEBp9U1Yrw3ddG5mU5mbP
sQ1Dv0TQdfUUhY73xOu9EYo34NAdo1SqRgulyV96/S+IsQUqZZX07MJ/UGSMIuS91dA9m3TEZLfl
GtEJmqp5kN6ZnF84lVBiLNhbs0gYave0v7uLqd7/jJU3wFFK2q7LYMHxUEqOMTDFy5IzLmoatRkT
gSnOemB0AKmNQxzh3Oe8ajvYJ/4kBkJEtq+w/KBjy4iz3AsNb2tMxN6EhBxJ19buqRpMohlrXx67
FJiMx/SNUIAwxyVbAkXQu5/mG+9e+8W6ZJW915s72qvpJyUWTSWcU9bu3YcqjSP1/6qcraPXBTAU
V8ctvke4YgvxJN+FhLLd72Abwuwlygx5HZZUk8NkQfZDNNtJJGbt3HLKPACdyY8zHFjlgWm6qakF
/QfNYZkjxpUrb3gewbLBOuKTy6ENLlDMEqf4NTTvLmbO8/OLGZFizacb9VOLZ6y9PBhhe6SRhofH
haBaBLKHGAWSJQe8C9h0Rjaw2DhNMngFkRuDm9iadSm8c+r097LBCwPnNhRXItybZ3GTBh0tmkof
9IqniEMckytSIAbJ4WwGSo2YzdwM6j4rSCkf1roiiit1ilVpVPMha09+HIi6q8yACpaxFDXFkHZn
bSTm/k3g+6V3fudvbvpHHyPb8talNtVW09cI4fPbLs/RfFwGyiLy+Lp4nnzVPq8ZOn85+cFepWFF
K5BhEAfc3RsEvnuz1g0ykYklXncMZ8C0zdPnUpOgVci3pAd1Y7vBdFPTYt4g/IjSffxyfc8TYgaM
rAQhzqFpqxWh2el3wsVykw3u9j+ebY3A2e1NDhTUg5tB222FJGm6R/7q4Dh5TurTBod/S1/5HhiS
BnMpcuRoTdKC83E8NSOiDn6IFW3V0OQMS/++IeLoQvhbyzAlxD1brTGWlD3BxS5jb6mUJxJbEzVV
fjAMurQxJmjWLeH3apQKRT2E/2oHFfWwgN71RhmXGd1jCtUCdlipaZszf826wdrQGckDxHgP7zdz
jwvR0u1Jb0XoUg8Ctmrra8jAVzg7DzUaFBXMf+6I0DZrGQWipIArhN4qn5naAczfcGTV2EGkv4/i
ZjsAsAHEVk+oX565h7jyph5tunvB/gOCjKWdvzgdC5VYnWbip6bc/0BI87BJFhlXwH27RhxwcAVD
SS8v+25NmPK3jSBVvF5vQVFA3KZwd1Jafbrg6/NFDWfkaNeuAAmtPu6XemY8CghEYEe1BGI9trKL
GnGwu+IsR3h2OPGm4qes7ah1CcF0NHNFNSaB1opbkZPKdz8+rADNCVZPleBzsrt+M9p9jsELkrLA
P3QFAOzy0bgp4qSKJrbNOUKnNs5Q1uP0zqrmoIFVcktQj0lW7UITTlB8Ff7sojTOlANO4yw+SnW1
4mBupK2nWiG2OmbdfjBohCbph4pJmS85jJg/YSOACX09y61izij2Ts46DL/M+7NFvfxBdbFuSWC7
vdk37kMGdmzS/hqq/DzVykhEuSBZLb8h9n2Uv4pmeY+0brJsA6yiNzV2SHW0g5ELUqLl3oSGQgFF
K7/LdpJmp0/JfYwxr5bY/JxnUEwgFkJiLnW3fnI9PiuV8QfkZ/5BAX5Y+o7mGFVZUJyrZMrY6Q0U
y3na2XlGTnp1xmtuAoG/gRDNx2tS2yeGp1tjxmdLgmkkEkMSzRsBQnWWAGssZ51Rj1D0poIxRfpY
EzyZ34lHr3zWQ6EUnT3f93zL9HR+VYDAzf5TgXgxAuZSFH1le3NGrDdOJvAr0mHpLR7IzwUr9FEL
0FAXV7bH0C6Th4QlB2U+qddyXsobICQW667JCv4AXPOGSXZ+7pMWNfKxbIRTCLIyzoI68tQMlTv1
ENd2u3BmMrwstpkoAmNqBlrv7J1c4cJRhwXCIAiazImCE+TMSfUc+8+/KfuTqM9ONw0XkLuPLUDf
HFEAzasPtW6JZLOu9RFGXB6PdkYFMtLpHcaf+Y//s/h7mqeDIjQNeQBkRT1GIdKebyQIhEbBAjcu
rALgeUz5mMnc6uCdAmgaKnm9b6x0AcKv0qWUoH7UE9a7QeerlMB9dnPiCjo3G/5VcEd+ytlNDhUd
tceilefNDJ+s9ghdioQuU1fmprXmofreBtBa5jGYG8WkgxSxY3DA8x8rYq91uBYS8h4BmVAlp86P
lvDkGcsOnucADu/7uavTwkMBgFcmXpco3hNLGg4ZHR8WTLDJYwiI7u7B3gpRNj6slUMRb0zL5v41
JR77hyIt7sdAxUN5YaX0Hw/UUV3m2CoPuxZUmutzfqVVVhJIigGVORuvNoAWM9GArUhkFB/zaUrK
w51ha23uUV4XbxB1poDagvPi2DQKlitGsgBVZcFLUC52xFqOcTuU5Mot+CanKMPSjUezG2YiIEk+
A9Bb46ZkEXbbBnUO8op58pRHto9kxNvz22IQf6QHXk5qCkuChLCC3+QV3MjrL5ZVftydyubNYjug
u6HK3G7zXTGMHcHsHnJzUUdNLikjnB+ajSo3njRiyySlYYzeiRXJq4FBq/hBQ5kpIf0qLi32maq4
Hly/X1BbQ4EwKMziQuJZ2NRxIEOA0ObLc7VpVUXyTdHMbLEeKrr5Mi3eMPo1TqRqMcQEbQjWiHcV
p0GwTiOXmSTfxk8a7+tI+xBujLoRXgr+lcsmZFZPPA0y4WLCo+mSpRezUPjeRSfJlA/9YfNUTVzl
JrDwiw1tdCNIl7ZSJCwXbjIkKtLHGa4y4v1+Jl7NpjHHJ5aSVg8oqbovoDG+hUIHrH6B0R+KI8PX
PaySQnyWudP3pn1kfXy5ZngDA9khbq1BOWEesIIhCEPdPAbLu3DYIa9GFaKhAwxg3GW85hCGxigD
KiOQEumPeaY1j7IV0Z6HXeBQ/MOFQfTkkqgPWCs0qx07gZ8rxSwhbZ4s3f7kbD6nfDQ7lH54Iv3M
xUJKhHDOtMoLlc7zIZiL2e4s/nFjTDRzsJVP7Pu10NwSm54OTg4F9XdN5mUXdA8HmlhF2IlXC+7K
ht5UW4uFpY3I2sMi52rtKD9QhOQfcyTyPjF6yVKnSLYwGULb0wCLNmzqfnqskW18vix+aq16+JMZ
7lzRUk4o4zjQuf3Y7WC8t7soa4wiGw86kvEjO21vRcS0AmwrUCyejD4KgfW38NLmBpilsNHMByAZ
UeIsOF7mznJcGDV6pDklUFOkG8UX6U3yrdcu6t3xnAVLmEvfpQlpoQ3OEMn0RskPMcq1XfJmb6Uy
U0+z+Y81g46DUgNfOIFf+pZD7GQ7cksBWrbhzkjscQGLFsGrQsUzUOnmFX9+dUxjlWKhGH8rXahG
P6MGHuLvhO4sy5Wox9UpNKCe9zlNZgu8siTOZuy7VMThd4mdHXaLigO+MbwgpnzHuvowSaKCjAcR
mGoc0wFHHPkz/T5518+6PCrRDPcyGo95v56HNH+K6KBqRTgWabq4Liiu5UxMJclWtPTIX/bsTPlo
v4eltHEYphUqAWO49cjeZcMoSIa8wL04V0KOQpAhfZ97KhK4JRi8dDRkMEVZYwKHdOwCPH1LmGQy
1f1L/G4/c/6t8ka/HbShV1mrnzlEVKPkitUR0dkKZ54NHpZpEa5a3Q6JyL3f0PUA/0xkipB/pxKD
/MFkXI1s76pft4RLLarrxd4F0Fa7UnSpzu68nK7hOdr7eKmYPXQKNKKuNj55ERxVpiXaarKCvxUV
S/P/cX5z+fc7Mz6UnbHKugmuWRpQ8Qdz1Oy81XnJOBsrUhjhE8ZS6i9a0X0bdNO6QdDsOYZPkIzD
rHCiIctRuw/hUUYmslGP+9BUAzUzRMXIWSdDMAyg1AX/7ssq2KYdShbzKdXVRdvTDAT4oXIP8oc6
X9l/I53sVYRcd3FXDf01aaKm9QyiW4WjpMGW20DXuI+dcwqYOXJ0I6KuZgM3HaFXGIU6y8WoOQ2S
annTVXzbRdUsuZO6f02kFYrNsyQuoUIwlJhZ2qpegBnNm9rqgqEipSa/eElGr0jYWQ+K4TYrKMlN
C3HVrPo39L/JHqe0Mi1PhS6OZqTjsbrXlxcpxrWxZjMhFBTHkozJaDubym3iW8PpZOcE9qdKAtaF
Le/ooyqHdwK0vC/9uOGHRzEx9h5M5RxJB+5k29ENvNKPzQtNsKrnqnWKIUIZG9wY9cxS0NUIHg7u
EiqHN+1eSCiTCtxWzQbOMWcOQPC1nPCc6GRmgqVxetZni+VyjvZnTBoQRyUeKZGjCwqvq+r5KRHV
Lk8AfZnXk0raqjGEg1vMVHYZOKsUXFRmv/lJ1ormmmVtje8aRgYo1YTKlD5BkD1rBUlrhNUuC6DZ
kiaXfoVRPN47lPHxGM1xRAwMjHKSXCPBxMis+hSZVz/2zEeXVGnwFGGruyEMpgszSm7+jSP220lP
o4UFQbEktccjAHEb2Q1mzFjdvFdVvDwf1u4pvMQXic3bDo7+z4zqWFo9AFcZBqGyKR2q8KGWkkvl
EfZAtJXd3H2PSXU/E/01UbhMu3b/jRm/xScPzn7aWPYACD0/1tWpl1LOLjNgBmSQarInT5j/1GyF
EpyVzZ7U7QdInf1JT4xdtBNMAEfSPKSEQ1lf4PeldEdLB+hAMZoXWwJo0DlygQId9gcqWtEa8HBG
IiAGtwL53tZrlJ4H4Vs4PB3NBccR5CTInHCQ+/G4DZ1nkSGWedfaoMdKY/+LlbvyZaAMF6m37+u3
nyHHxlXmkvYMppSFzMzH+EI/9DQCg7WuH2rUpqhnsLtr841VH8ACXVqGXxjodxRE9ieQ8/8jr6qf
QEjvnce1yK/vqJ/v//cwxyjqRtximhYCz1TMdYcUG8IWgyYnvycd6cgoesauY/iKxYwIk6wvzgw1
34d5BkYuXIOxGHiDlVe4bxqQ6FjUNVPUfuSD2rEXmzt0sIeURNdV8hwSnsEphdsrYZJjcv4rxbZx
CPI2s633RhgeVIrI41f1XPz+7CveT74mMoLZGni+KNBifVdo1O+AAnmcrOvxq/qRssOExNeKDi2d
N1mKaGbfXkuvbzIK48pPe1aXcBUjJT4V/Gxo1l4QboG5XcpyB7G5eklFXOk00PTUQPUaHNYBVtdq
yjjtX9re92Pn+tB+I9Wv1UBNYS8vlnM3JTgmu5dyfvFCog901EmqeuPfE1/T/d2zoA93Xu/Xs0Pr
G15gKEXKcCd3tu0kqznsDNZh+++UzoXooR/lQT/1p95aIT+uvY4SSpu9FnxShRU8KVJgBeSi7HI6
GN0z2xtAIQM4Wud8/LqauKEOqNZDXMmbnKpJzaBmpRi48iSG1t79aksCyW6Jxd+hyWcobIygn7oD
gX8pa61RgndQ/9KQViayi7qyXvhTPd32ZJNJK2twL/YU1kVBlODgFxlXG7QOUuZQaXNje7KYbvJx
GJay4UVcQCGx1nL8TubjKEt8v1qhbk4shYWm5UJdHL4cMW9BPRi66kVwusC974u/fLWYtp9io0Bg
fz3FucOCHLsK6nr6j9dNKWp/mmG8r9PMua1Mww1jjgs/DysXpkKIkNcgUSn+7tELPbhhnu726RnQ
W+6q2mDXzORaARKr7i36hhyyFicajgeeiNg3RbaK9NhZyQ9ukNw0RcGbMiG+30SPLG3k+iPqfsOj
bDCwmFmQI2rCcTskEszOpD/PFQB8CSAUsunlS932VovXGP1hDq3ATV5eqPZL8cZ64CwCd9FCtYdI
SpoAUO+0PSgagPw4vR66VA5HpFzxo3slFRIH4mbTuOJlb0n9DL2+2MpSyD0XnIsoHRIClEuDpT0/
+0HuiJy/OrGQKVBDTA89ZuUzDlRGiJ06PdtVlGdxHN4KG/PADslJ9WW62MjGZbCTY/XVh7dc3Rd8
TvzJJDo0iIepZuZd8M/nf0XzDq1SmSK06Yt0CVjLgzfi+4MC/RPqWxEY/Eg1m7Q3kLwVCo768Ctk
Z4msDCNR+W2rOFuEADCrWo7+xtEyma8uX9ndrG5/2QKSUsQMwBhRIEpn5oA+XBNMtMTAyruU5V2L
kSAArGsyaR9K8QtWD+asL/mIk79Ft5fh3ZcVTdmq6+nH4KI3ivfPhTILYDf/I1cem8dm+i3YDIXs
2GlZzieHRewXLw+8xBJF8nhYoMxBTgFmU5qGiIpz+O/ay8M66L1xdNy0NvZ81msehBRrqKGQhOnQ
dgDGspxPSSPjfefUhYbaqmb28TAY3DZasB8TibXFK958LlHvuX/UTlAJjvqwZttS4x98u6N73o+m
8JH9p5Yt/ZNqmFBvA0t0EO6dH+KdzaqFUQ2g/pglXfCC9xPKJUN+gtNSmsQpxCRQzZid9I5p2+5p
qtDrYAI/zttiQhn6pdmlFIxIkvUSE4BBlONZDueryE94zs5T6gRPpMJ+oe897COx1yr4My5oDwTT
B3dcoN+f7hBjLj/Q5mKZHjCn5cQt+QKWEeJeX5aypoHApegFaogbS/meuJIGvETTFQoy6eG4JYur
VegMIp1j+Ww2wLQq1WnQHwqNbwL5SgzZhPSPfA3mKp5cWd9GH8I8OJ8+ZvgKorIMOD35ccj4hLTU
BtRuP02SVcteN13rc1U4HnwKEarW+Ukn42Me5G+L86Nv+nbuVv++cstbt6B0T8zg6zOsH3YTXefA
QX4Ta/k5OB67aV3hylvZJPdj2W4wh7EQUgfQm7epZx3igz3k5ZSLFfGqfulei3+Pue/9jp5AW0GV
aenj7YMH66hGojEW4Wl8nDM1ibgM5Cv0cmWg/Z7cikHRLhZrmUEf7nu200KA5GFSKChqLIFXouIh
KKZTtLK655dVMQjfEGOpRpAL/URJzBDNtTNjxFT+zXBvr7neXhvZIrcDyEnscAlDt2I4GHc9mmf7
r+68CMf5IwzfhG+KjjngKseuRSH0t81xqF1bCTTnRqCG1MRvYeTMFGOi+O5Jo1FdBsB86InLJDo+
5AQzNB1706PgYXmvwas7fdVWpgn3YAIquXtdZkiAZ2EA/H6tc9RrqblDGT4KJ/6R1foNs8jdlmnO
cYnowXpDY2L0M8gCJuz/xL4rsNuGrq/kkmSX4HUw8vAPPcRaApm5BQIGm7zUCUieg9bynt6qX6+V
kSJPxKi2QxGLtKSdKd9y5H7EvGMdiVC7bbmTokbVED8b/nB20mR/UHscWP1MzZeG+2+a96oUetAJ
6YfTzz8VfSPgCwWLM6kr3GAajH0pVIpa7/QckCnkb1C2XUOseqreNf6Qccu1gSqxIrySorJXbNVJ
xfM+2ES+hOIzgAOnEASVHeGZXSv/lvQPkn2IbilqQmOKz3X4mj1+frRS9KmT8DlhtOpI6616AXYN
20wAbUBo8jWb8DwcEPfG5CM1rZY3IlHCoXkh27ag2QCMdcSOXezXvk5rx7EKKkNdVgP5PQXJ57Dt
ME2WO31vHF2/izAULEQKAoyBaiGTGWO7ObUBP2ICBDseOJyW2/B70wzzVE7/aeNZA2me5kBJGBah
Mbqx8txbrRX/jj/dkp6sFlnyI78MpEJy6EiDDxztDAvwcMh8o35S5gAYKoJxFVgAw7mgqyYHSNCs
phVYy6I72V0HmwvqyiQmbuTKDe6DUzUSMrGnloANVaEvR+u2lXJByTh4VIdM11Nfx38RIVdeSaiV
vj2rSeBFV/joX0WcWuFEH0L5EUOIaXr5/LXtIV4gP3l8RowTDPho7xk9fBQBKikbQQTuIOc/2y1D
ixFBEVnxaHrtDgHYZfoL9MC1NS9ULY9RGOzreMHKFH9/DHpqzE2HFbSt+2Av8ZxMC+J/Pj36hwQ4
TX1L0CvaAtY1u5hIz+opZO5GmjyxFhbWCZ2HI0IZ76L0xyaxznM9ySxSrxMw+kbIdPAafW4QfDne
MR3TvUGrHGJQ6Np7gvyc86gEZCgfvaIlM4SvbQxkw/WfbQcLmsYfnpfvCGIRyr5imshIE0o14n2O
MPU2KrvyVdD0XXzBPKHx5nIOTZNLynYiKY4NtRJswS4AO5Hma12tEyFXpe9Cuk9IY+J3PKaxVDdY
JVugdO+hp5l1BQwIHwu7+votr0hwXCapX1YNuSy8PGvLSYRwPbsdYZtDx7a9HTCEWDDl1Fyoetfv
YLohQiUmBZmTy3lhEgm5RfpEF6Q42wr8/3amd067ElTNG73DYUupygxAap1P+PPwAZPLRBTCursR
wEySvik1YlNLA2TMjRmx3911lKVvjQ0FXxYqsL39nIuokQK8c9w0NsCS8bKcy9Ni8G+v+IxYb3hr
ivMEAoTQiEkmBcl7br+l/7l71xrvE19rEo/h3vu5mMaB90cknPUZt7zNYjSIgAnY49Lcjltv+kLI
f8QQUOlkcSxbAqFderq/aeQFul3iCKsNqR46U+W7jFazPtIAtrOwpdnIhdmo4ojsWyWiF8r3pAoy
PTPvxiXCIauTEzkKEbWyXknuy+wZu6vSSgo2gbL8SZCBa4gAez1oYQHu+pK87lG3GCzpEfO6So0E
R5yMkP/32ZNl1a5ozajorLCoXNnKEYBuwL832o/xJNA4GuqobGO0PYm/5XnILy36J2e7p4YxqNtK
CoLapq2TxGWMGxJ/HzBJMxz+uAu9zhZpvBVfiShNy4cVrOHLzdzEUytOk2wqrfgi33Ss6wtXt93m
+RLU8qyCN28X2Y7JqOPFyAxaXIdC0HLGh9ad7SJn+4s9jPPWY3J2avpq0BNm/rYfGi0kuuoNZmF2
CkIFyaanOwjUp6somuAQ9cUl8+lKVej4Em8I0XJlRdlVzAyF2ZIXbc12GijQf5HhwbTPQ0F2iUzJ
Y3R/4GzeuyPL874VC8Cv6O4rWShKSb+z6ZCXbAIQMQxe8zBfwi7/ZGBW1ZePXheg1xiROxE+7q7p
I0SbpDqvO+6PLRbwZLEgkkIp4NQnVWQiubWP5BcWwXQ2RAohsLfkpgXiPB5LUI3qoIF8LlAT7gpi
dZec5fuUzyQXyizn9Y8hOVI5AsiDZeE7+qa1oZ6FthzBndVlmfMxF0gUnMduuAFHtRtLcXrukpvR
S+CC7OZS2OWrLWvBK3f53dr9KDjd/NLhliWyG1JIL9jENELP7x0yN4SwwNQQH/PirSLbuQlcUlxM
cEEMtG850a+rzJLG3mVPVS82VRyWRUOEkLSrQAAEXVv6EmB09DYXpO/I8/DY4QoxCn0psJLLLXyL
Bti1bb2PVBO3rabSYNw3AwWYbQw0osE9mZf3Kkq5Ik8AcV81UZofZ1qVs6yD/VXQyV1buY0Vh+NE
uGscs/TEVbTJGjIAl9+XbFDiv8GIpZQOTzBj0BBRB9qlualyGnj7ERDcuTV+OHYde8lmn2kvK+ey
fdQE1xnDX/nhIBavhh5qHDjyFFMm3yXQ7KmszPl8eqb66L4fvtp/NVXNu5UVUpP2uqr8DhPckSSn
Pi8zrd5JaQk1EWzlr5kuykXQvADxZeahB1SUCrkUhyeYZIsDzeDV+6Br90tPqsq0Zy34DygghXU8
atSEq6ldfZVpZfgkB6mucd0PcZv9ziITdB1SL8mte4x4juKF3o6af7VmM5x//X0+CcSe6daMssuN
QVZwIZZiLwtR94qTBo40piy+uMHSDBw1UYlUzqNtBydb1T2gZe/DopBqUCA7u17WOvV4u6HILq9/
1hI0msQ5SMikNRyadHbAHWtOXQWuerZWWwqZHMTEJLgmtC0s5XSO5rZrPgHMgAtHJffmmKukpCBw
EijS9il8Cm1FZgMX/rHpru1tLBNjXdBU0Yoimil8WaCWM9RVtqmlXHLCP/yWLvqpI5kcyIkJhD85
lR5+uSLYqD+4WgrrK7F2yKZ2sIPUof2zSFBn3AWwotvsUDra6Pl1I19oAc2x7zTO//Ky23p7sf2U
gaPGSW2n6Mqbq5XdSJFkYRgymTFwTFelogvRZBYUEeEtFxLXLkgq1tkoy6Us3H0VQE5fptpPCXMf
Kspan3WPKHRG9UC7H+Y/9IgV9zzJyHj5MXzgJDLjto+KFtJew5DSGpSsr06coZacPkmsxVJKGOjo
GGNVFQp4FVifxmt/PEUaCedDODeEfUcq5eUB8L6z3xL84hC3ZOONZ9ioBvxPG7sKz5dO/75pbDgh
q57NpkHfMSy5Mgh1kconKDibQdHXKcrFrS10OulNdoxWprLRw+IHl2FCUB0vXSjnz/yWQcTqiebn
FDY50WwN5ZSAWMND11L7J5oKvEu9sfOsAqUG9IJrHikOQB0NogSXzFOKpFBxYOvYo8MHDNF/qk3t
HYPOyMxDXJfFBTSaEDmouz8tqD96bhuqQBlMrdeihcNLDfucNoIzBY/iuYqgbVwa95/H6IlYKy2q
2C9UeQNGin2rawsoY2ObkXblWIw73PccmQa9BouJrqoZpIYmlv6GDHmX5yIyItU1XYSxWpAbqeZs
sc7fHAhXe6oOAAIO2PkhCvGKEMAYluoARZllsL5yZG3C5+g3IEPCFQxhzYmZgQGM7EM8fSn2snk8
vyDH3pl8S48mz/8yxEaCM2/LK3Ku+PmHzK+oI63wiHpIqepKRO4SuIw5Aeq+BAY9HSM69nMGKtUs
LtqUnNfiqpKxIGD3WCqnkhqlLOeXa7iA3UPQdomPfMn8Z2onCPH6dv5sKj5xu+5M50K8vBlkRNEt
ZllHXLIyzrw6neoHKlpiis2svLZsJqwL2CwRTJWEIbxv48dD94skOEYrOLeehMJYwmjhpZtbgVsJ
G3BPwNIlTOOlU4NVJX5S9cN+XkcaQZMzJPSpk5Yvka/7VKDk5RxUtXV/o+rx+puW1NgHiaUWl4FZ
IV8HHcSlWUbT/TdqmqOGAWdxm2bkm8YPWltn3nFIoC8YNbgAFe5nc7WFlR8pXTwV3VR6svxsog7V
czZ5gCstsym+SeIzUhAXXA65Ont6Se0Hc6k95NLeH8mFCYxh92vhTolAOWbiqsmO0iLA3OwDVdfY
zmBMxwCkDudns8nD0irnVev+2iNjg8Ww9e4xtXgv1UAKu6ErNnAs8X+0oOwM/1S+cvin/PW7zRNK
RfrSMCJGfqJRdsF9eiE8eY+1y1oxAKCWYERv7SIVZPC9KQ4aocRfJImhNUFuEPcUY50s2xcseOUj
jd4xYQ7wyuRnYo5j6S+vgMTLOT/JlfN1f3hTSlGrmgcvDrsaUA6/URLgHr6gtUaKFx+8Lil2edvB
M6EMUE7WD8iPjbgcUBIoZcmhwFhu7sBHWvQUIe5iEBUI1R+bRYblMbcblHrZlzWa2dvy8/l2lASt
2fQvWNom8qivEO+aoHNxYvvMJUQ2m7AUE/j4w6G1YT7t+MwfR8SLXSFJF12oW5nlHW6H7r6jWn4p
3QPJtl7meGoGOdtDYjVrmgI8J5p8Cm1C6S+i2OYLpAMOHdKmpg37XQIUTuiwowxB1+N8VbgDQeTZ
7/+60eBK59bAopOUv/ROmGvbYcHnFD+GCbkSG0Rd5m4awWnkry1NYXD/TEmODTEiT16Gyt2D42bj
ak34jVxLqke27E30Lto/cmVB5wE0Oc8hmsI+GL/ZgijnSQ3dJ/xKtXrrfyHMYYRHBGAMH16A2Ri3
G+xE4auyz8CpfnkPRGqxOXoXmbzDa3IA39+gy1ZGaeo9CEVviSN9nR3QOMEnFlg3CA0K93DK38wc
D+f89gzhkhMz9nDNn94sGzvt/JKmwymmTVSTJR6MHFUmI61/aud/VBLkLwML013DxLgOUv3oKW8Y
51t9aT2P1CboatVxK5vmF26qPJ0sdCLgtvgy+SPNkMhrA16k5jx0kTUa3EbnpPEbn+79CJT0iFJL
gCUBQXHHoIVPIi36Q9xMBKqz6p9S/uYCGR1NsCqpxqaEeVT5q6xf96xbKf0GwTrL2bQt6+CiDorK
1hCluEbQ5oLSUHOMQJ0sdn+8HWnFNa8G+GRnP8Cl78zrNh+IVdK9CCqHt6M2RoixQjvp0HuAeCLO
/+csJOEuYsvB+e90Z4sDa9Yi89ke6+s2aXPEtVaRxJddB1M+W9o78RKsL7EqbzoTbnVKdv5L13ZL
vghrSn8KQguSc0CgN9ctTwdx2AV3FO13xww6gDc2xtpgAYix9YlRJ5bZB3r4vH7l0WDI8QwmKRsa
cZR/uSj4hC6wgfI27AmJHFjNxRSKtlGOXUmkhCLJmW8s5QZZMlbroMUgMa27YlKmG0/SfxwjzL37
b8ccHaDK4hEt0hJNyXCQ/N44yW/ml5mv1LcFm/gCMa8dENziUtwg6DDCj/PFlP9J5sD64jxO8U3M
sdEVP1yrf4Vk8q+AWIkbK7mTymWZv9u6IpcvDOTXYjz0HY8ouin7A1p/Ztu1311CctvmZOFF5zXk
Wox1gdHl1/xjDDIlOC7PLuFRjPnPFv5srBw3wB0n+q94gegq672AipjkUSqDiKuUvZIK/5wEdB4o
ZR//5L1bRXteH8gUSJLLc4pEjGpeFZiJObaUlGIOUG0C+iyiA9Ep6th8cYcVx816QA3k0NgYKr0X
JpX7ZoMfj+jJB7aMi++mj9eqZTD4aLEGSJzmgWo0mmUdeTu26VUIk3ytei4CYRnStkAVpjaFP9D9
9M9ODnD/wYMuVOb1S7WxAtkh1fPE5pDvHsCqJcYFZhmPHMOspWQyUYUDvcim4yhu6ZA2QlP5vlMm
h7kp5wsccWjQCmcBzDaUGuGyp+2/PqF5BaPcXGV5EV3avBYFKCXJqnJFUwqfui/rVptIfDI5bymI
Pf1BU47C4B4Y32V1hKcooWv5nwOCz170fS8ixztTlWu620WfAv11AJ03RCzN4NfamZq9d+0olA8k
6WflFt+YJhWKPI+n7iGs8L8poH5tQgF0V6wQ+/wPy9+4gVcif4vhJYtDMrXQ5tu5fTtv09h284Ik
aEn1DJmnhnetJv2MycTMMa5zSRwuN59FrcjJIEn6bPEzAZFgi1gnbHdECLUKi1q5v2eVja4e3/1u
Pb0ReyK+xUfOeBzh5J80yTRCRUMX/P6fW4UIm4C4QrqlVprS5qhR3axhuTgAC9IOWcceKvifVqb+
tzhpTC3eFt4IYe54cUoS/wdWvY0CfwtNDr86o4JOmgO7Vzdaxwes1JWuxhzPTvFuAGItzs+CUGn4
EOh326hYExdmKltVR/N7DaZftfJI0DcuSb77yRwVDg/aLO7Tfb1CQ8gEFZjTiAWAkrEXGe4wdfIP
edpakNniqxm7PByhGA6ndYgE8xyYM9uozXA8UTfl80IUSXeAbYc1pQHos7GqxR2XLJ+26/sA7O5K
yo5cnG9MnztzFOahh5WrN9Vi6FyqRSnJ1ZbDp4M4cUqzNA/D5XPCC0mlPaMYR6QkKsc9oZvZEOxS
mbC/SFQGu50ZPuQIdp4i9YOBPOKMrdsBos1jorjJhdC1+v1A3+lW3MdjlQs5tslmd3ReyCJ4AHGz
sxdKpTyK8V1nbcvO35aP1cRkOfuEege84ZgknTCPwXE1B4gUp2OkH5XcGttyrmb5Ke9o36yYFL0+
TbsnyuNZPpk/EPvKJQT6W6otBrkh/KB4xbkcrJECOMz86QgW3CssDltsyGg4xHXsNjtZnrPu/Zr4
RBdWLbzTUER4TBmTkm9G9zdWi09vGOzT4BxVFv4OQRV2ySu8UigaG0nO9jiUOQkQ580eaa78P8oc
Q+Q54iH5HI4qGPMIIQ4dd8AqIpNHone5kTcsEZYOj7Cl1Grm7VM41OBzBgX8hblJxkV8OSuplDRe
xqD9Oxii8U5pi3HUa6c/7yLuFPpIrJ17ghhlaN3P3G0fTnNLZsUoh6CqdBlBYvjnSDB6N8MTdAlR
XC4mjLviKz7+ooc8X/T/9wvbaFdJKazymuTgxOXxYhqE/Dqj+XM5oMnj1nSx7CcxpbNlbRVCxb+a
cnJFOB6fycjamqr7bM7C9oL6wzgBs5ZLoTm0k9rWOA9SM+Njb/r5M+mSAsE7UvsCe/q1gAKpBxN7
TRv8t1KLtlm7nRUBjj54d95PWAuu62Auuh1QOTykaeROUFmnaa1GsamRK4nXUhM2kXotm4tQ4adM
2NugxYBAmTjBoa+Vd8o6HCFz6VXG9CCoyXS1mUOOsTnqSrrvdEIAf4GiCoyoq9VBqQtoZuEzLWdt
UuQILb+xnd/uxSy4RQN6Zp7CzWXD0/gNiaaU+2E6nCzKRG0vyInxBLtSBhn/ITrtAQBCLzAQy1NU
0ALsXT6oaKW0bUy+xpUDD4zb3zObvM6AlpEQ0GTJIydA+a7UMqCNLesiV5dyatsrta+q8tr5+epX
ljH4kQ8A0YILOrmvLCMYXSXPBYnOxJqzZ+/tJ6Y9ZlJPhl4NqiIJPScWeLMlAcpAmoS/k5/khRaT
BooTke8hLjs1p8Y6rl0UoX66PSPbmkhj0Q7F+DJFDoX8ZfSS29YOjXJDqdzhnkoB1609ITTWmEQr
hVVNJhhikPbdJmeJ1zqYIcas76td8whSDTipAGO0k/CC2WuDzVMRFvTiXOOJPfA8U3czeJl+PyOr
T7KcuOtMqyDbvA0uVVhlxpPote8ifA/vmzHGe0FRCPL9lvw4DzYwwi6e7cC2pFFoqU2hTIVEkHDe
ePD0fEtZRWysX+jjjpbF9egfYmYVtn8SccSnE+jq+9oIBaX9oGHEyOHc/FmnqqkXyoZYtk3BkgTi
6mMR1JI8XeOrrJu69qMEiOQGjOCFbv+vJchI7CFtgCU8YhlEe0eMAkP6J45qUGkAUiuLn6IPX6rA
KlZaWKJanmezB39JvO11w/TZlHr9uXqHWhUjdHI2WJT3oDsw10v4HhxqONAd6WFCCXBT18DQHfZ2
h0Rg0ivxVz8TCvhocKttJebZgS7w/h6C1n1eqfGSTA75jn4MqpOQexU0y/tXvG3Er4929l2e086R
oEMNy1i/uPKoUCqZkOIfXuacqImAKuimKjnQ8ODBtv45atlPcAzNS/bkuUj16D6BryAEz2ieRv1f
HRQZSf75T5HWfVQ13fASB6E0aOg7EiLngd+2qgdJNeW8LQwJ+Vge4WxWbJZBdCyP/dXGf6THv097
L1HGAPbtKDjTS9Yr72/fgiVNstzF4GmARiKQ3ZpOfxcLDdlaLTT/o4h7Wuhl4PTaTVcsnvSeiWdJ
WQGuaoDDIhI/SQQHmYClAtBQESmTmvzHCucYmfeSxhlHkBAn6VgtxwrxLwUZnm3+snn9fNqu/XkQ
48KA1yuGIo5r8p6L20WEdvrr7YkJH5QCicreYPcEKm5tBNH+1qEvF1zxetya3wUVpB496KkjhJYT
t3SNiGaYZscXkAdujXEeZCkZAGhkHAZLN9TA1UjVHV9J0ClSrnCb/NNGZXc9BIwNO/BqlAvHQXO2
eMzromSpeoDHePxX6OCizllmP1ogB9uYr4feW2u4Rn3AM90dqOtgGPqxTHN8E6D+Ie3WySJSA38s
vLeM+kFIEZyM9jpJ1POC5p0thu+xYKIIjC4VI10wfwq5+Gdq07aRI8tUlGA+0vHqMAiIL3Tp5Dp1
2dBrsczXRB07kODnfsvrBBxGWHjfRrFMX4TThfXhQqfsAzk36bqhL3H4ZuQRXBXpq1ZqTRTUhDJS
CASpU+KVwTQlWpiMi66KiQxCUWavD+vwmvc+y8h0cPBHOR/39WgiTxk6SNLsTlNsaKshLvGPh1zA
GTbGqW1BesExIpfYeEP1zwglGe+4pMTn41ajr7b30oSSsvC9k5Ll3mZdv48vk4exRwtaGjY1ZBxU
eaU+I9i1WC2rxuePtmY+s28at7HNSIN2cDOrP/DGq3F+cMNj4hLbfRlqGR7hqzQBZpWDlcFNMTIN
MywwCfdd2WlhYQ6gEksl2qkkQoxxO6Sgk5vay+CuzNNPPPzWPuRyauuR2ignPciFOzMgqaqVY6Hn
hPyRXxQRoYvwk+2ENoPotdVzsUy9tWR7zjp21wrGXG07R51JEU4hbrYG+ra/cpXYbb6u1Wyn9zxB
IoUgeUzxL+O8smZVpDjfPz4sePH0O+6KquvgNA0/dXb0z8JvofT4CvC2UQBHWnbrD9hHhHFQTuTl
NW5b+FgtLa59Mt72JpNCSSFyust8INYMKp1lOqg7M1VggkjjsJIPCIoVR5fLY2nlAsYcuRDbZYXG
91L62Vce471BI6fnPE8j0Mq8Lv0aIEjh4hQ/v+FjDynAgazFhKP47s+Hiy6qxfQt+wcQgdYsc+Bk
OHskKVzVgjCSWLiXfXQ/bZTL3QIyCP7y4Ht1oNip/BSSXa7V5rb1SkaZ9xTUlFjGbIUV+QBbBEKK
SfMPc6g3BS0niqyV9J33PCT8XHfkuo9dULmunMpnqieK+TO2Qf9ue7UbgpKmSQ8LDsLExCcgiXrG
9veJ86wOXw3kEOVQ8Bqkh3hK69jJDtZAUuIjqIR6pq15L57SsjmMDHstHdRd5kqnty4MdYtZ/TjQ
Ubu0dM+76aRIW0qrS+n15k6GasvDBXL7tauO655YFVrU/Is5m78KIChu6pT0WR/g6vISCB11928O
xjVV/4GLWmqH2GMNj15EDaxPXhe0T9rdkiaK9iufNfkAYtZEuUzGai1y7/FnO2kgYwacoFgj2JQr
mR+JipZ3UTeySq193adx1udda+a+KKog2YoXCoP84hxOVtfXqeAGSkjBHHojvWHV6tp0ba56apNC
ViUoXdamAume6k2Ye0qPQnn4j+kMeGQPJd2dh24uLvgYf/9v+qSfO1k5t0UslienLYmnQ3nPMPEA
kteJd860kCf1D/XLQuuqsEagyTbdprDgJedETQmkhxH6a2DcfwJAYE9XJ/IrmYv5vYeXl4uPKDck
p/8RzrnliWWO7FMQknu9lgRq5vMMdXguvyH8TahTe1iIztHSiERY8DMxVmsapNLdxLK297iiZexH
3LGSVSOQk4xZcLBH5IF0PE69eTVrV/sb3iu6MQwvQpIQATWMw3/i56TzQ8JkFvDMhvS4WHvwCPFV
2ZLiM9cRWGbto2Al92CSAGjO1e5kuBnMFlX5xpVFpYhSZpZxg+yVn4eXMlqWbotmdcHisTAM9W7Y
daLsL/r9EXuhCMBMBu4mu11Xw2hOt+czuPYlQTl5iHBXvDgZSA0QzwsfCgMlxFQqoIpX5vs/q80I
7W23R7JBNaSaoXzPpLH5JTpn4xiZf7OwZxVKk3lmNpUITeOG+0j0Fm3+iiB8LU6xfu1FgrNIbaYQ
72q7ilpQlb7Zxp2LFPVylWIcH9Kp3fWysG3G/b4ix1JPaLRiLgcCBwC+AHH/t+vchZKkANqpMsVp
apO9K/L98g+v6ED1kG/s28EIoAAna8b0MbhlrPNnkqoA0Q+TmrjpTVCNnfYXg3xqvL90C6M78rmv
GROPM08cgprpp8cy9YwN7IR71hjCkSM4FcrdqcUy6kjr+J0rFARPgKBeVoMYFKuJTl1/s9yMpYlb
ITRBPI73czAB5YRLBmL79inlxKlGfGsHgbYUoe44Ai8RJB+x+zRkwOR7U0ojeW+uuZ/i7b1jQa6v
qpjy9+GbiL/FBuL2Xo80jYkFhgt/7Sx1CY6MdezTLQo4jTw618S/uYgkWmsfzLPOzzPxUNqkf4fK
Eapwsno7MOWIZpEYurIMTECaAyitY5IwuAfUCUCduAk5ghHWlq1jEGIn1VunpUtONAC9zox6xzLx
SdB0Ym7hp5CRPYD9zBc+tHsVqWdRfRMYgizjHpWw3nGffL1q94yBCXs9Q9BPiojE9T4Ohu1qzEAh
5946XORUtuwMaZxYA3U+bTi2uXWhCvjjx81sp03wPVEe4gFbwo7lzOQXPH/xi/IPc2SACyH2A5Ce
ih9aWG4uXY+H6zpiRmhjXz7gUYvWdxDdC5tkZjqXqPl3yqzEaL+hxfkypmvgXEmjjEPxmDOu6q1p
1T2EhE/PQc94wHDG1dgihFGbgoixWSqtzlB3R+WF6CTUQj0ouuOwVliex4tK+31yWyQKp/3YLaKm
Hpo//wnHXauInE5lvC+CPGO8gS3KcwKM+K8bs+Mbu/RYDZwjwAmddJeu6THic/3Yleu7/mOq3l2/
FLj1jmNfjZ0p+i2aGCCIE0JqJyzdkEr+lVKqjw7nJbo+36dZ7ixCVnzvY4XPZ+yxFweNsoin1hi8
RaS8pMk1QJrTJrUFvaR0mpB0dgmOlqgm1deQYyfHHkEQGejnEktPY/Of0E2SCIX5Yn8ntXe5fB9c
6h/9wp6oRA4TIZ74sqbni+ZuAOYY2aZ2jdAWeZqJZ53W317vnHPJF4nx6U7j2xbXvxavvPJJYVso
2MUW5YQKLEXAr5B868DA57WB2F/jQBOVp855KL5slN2uNPO09Ts6dH0xwh9ehGk61MCiu19FOEoA
XMY04G19QI4HVHEazRwuy09dFf930zXVnFmkwHnObSgktnWZG7g8Dc0mMJgubCSwN54VoEqA52lb
wEs+HhsoPOW4eLOJxXeOS2t/da72xKkLyhngDDp0PpTixuPvrf+kTe2UqKx5Wctpx7za6MlFrxKR
8AY4mAPOUgye5Wy5e87j7kKk5sj4Me+UCYYeVh9Tbp9SHu9F7ihYADPXDG9Epmofh3LwcmTqEsnn
ya01K0hQGfsn5lkH03bhXykN4PGU999T2fY4pLEGab/fECtnRi+MhinduuOIBcf6Bbh1pRVEvo+a
9lA2QelQRMxqQHb5ZHFQb1832jWA/IbWXGj7TVN4NoVV+Xub9JekhcvxXDFESXlatsPPvQv4wvRV
DpkousJ8QtXlMY0UqPNVDX09FhwSDcW68m76DYhq7eVYwIOBy/P37OkwfR7E1reWHjPU5nOMcNos
sU/y3BaFMT+5PC4/CbTQZy0wTyfuUYRuiIHF+KgfgNiOhNn3HdvbZcz1cD364LVlKLlccEytH9A5
FlT0m2unlCkm7wxfkpFhtDmSoo6dvtS2uAMMZYd1pTSD3ejB3fPFm7AROxFFCtk/AAvlEBgCfGV2
hs/a2MOhlQPSEs+1Roo7p16JC2BafFjOWpwS2hCplVr6Zj/+X5DwvBJwaGROXUOceLRFgviEmw7g
TmEsmCH2VYFjxKA+5c6nIipqcqYw5UJUgBaZAi0oMPTFxF75nqWHjnLmXd7y/HO8RNgTqMC+fXla
zbJz1F2rqWqLQxE74bycqffWVLqZwdKfCJFbGZyb6sRKcdfuTARAgX/0NK+r/F5tg93U1oPkKPOd
h16Urc2f1l/pXY2qiE3nYRZQI5mM0658nFfgob5S+9oPfce5VJwwqreGNhSGYNLcc7Bz3LNyIvZT
HADaI1W4HPZsraobIHAij3/klpSBRh78zPz/ZovIyhBzbCz3ZEo106hmgseqBUMh+rnAprnf3eva
0i/Xpmed7xPC/X916oCv/ZUj9rOaMQLAdcK54xdN1KiXLIFxE8fUNGHHTlAmTMbe5DhQOMogUuAR
rcV74ZmZgaXXSPhR8IxVXtwRjRC73p8rljxvN23gVu7DtOMoFSxUBeNG4rcxTU+KPYK5HqiwY/cX
8abXq9qDPIxGA2WuG6+Y9gwWGYMXWTlxSpqvqb5U2xuzyZ1iGxpILDAb8hMee2nR+h5ChLoG07S/
KwXg3TQEmZWRmz3O4ssjgZgMJffDWjrRvRcJ1/Z/8v4fNYpQ9JZUmyjcy3Gtx/jRV8g8b9I+a4TB
QBSu9Y5bMwM4/MQ0TrtjFOfHlq38Cm0GAoIU3d7bX0aVP6AZWDw0ttXiLwVUfGdyTrwLZMnpuwQi
9XOVbNyf5ItaRuywt++vCH/ScaN3R4VJKqObSM//TYohgMAcADNJNLFlkYzmarqnlAdV+5JYKnuT
hVCZ4KemL2Gectp+ROFdv7R0vKcFbfwQZk+lPCLkIqIp63k9yno/twwypHzMcamje/rHTMm71DAI
5n5XMOrlibKbi2z0V80boEJ8htH0A9ZgPOtXZfYmpAqH/KXYIQKlUlwrwmwhvRCc6useFQWHyfwE
8rak4AH8LPG5sTChYZSwEruUygLOcsr7YuLOISojdQlQJE58nS345Zl8KVQLFUBDZ3qlYJnFdt3g
ayRZ4kOF5EV5ckFU+lLOxmQXLI2D0sCmS5xoEMTqfYC4hhMXpngaKQGiQ7GoRaagnUvkAn5zmPQH
m4KB87OA5bFTCvpyAvwDN398lvtnpVKM5jC9UxtddMGSfVM1rdvEb+zp1Y2zQTTkptNCdUnTzVDA
fDT0PBEbzZX1wLqcf27K2+ADekeTF0IK/qzELROfaxdJN+3N2ID7OjgNu5jXkaLkpfJ8KR9E0eVX
oKY2j4zdfpmiqab8E0SLPTB1vsYNkB66LM5eBoLAaeBiY2mB0xmEXNOE9xPGnQZmUvmEg0w4AoTf
7SO/23T47hYkftw4EwwxD2INFD0odcy1qRJWSm/36JygKltA8S3pTfZQWr/2+rHiy0JQ/Gg2Xrho
KlhUZLaKLaNXVHODfVbkwuXBQKucaRYwuHF61bbEBSKANhxzw5ro0AH3iXPAWccXyzELIinBhoPG
C2H19QizmNF2weLloQPkKYlXdQ1aMnljrAedw9/lchZxXp7NSOdzbgK5vHTPKj07dir0MJrEPM1e
EMHZ+5RouEKQT2K72345rYcgezre4MH63HNBMy9bEyZxz6W0qpMLtdelEucxe8NDtj93qyHoV1e7
cvhytwPrTOrnff0pLjfcTYIiJChchecsLK18rkz7Aez0xqtDUXxjIFmAVh83Lv3JyQLRihxGBr4D
Ry/2tvVZK8ZvziguOe3tkHDqfv8+EPH1NfLf94afcNmiV59RL1RBZLyD/MZsdXbq1u3sLGt+feTd
/70TC1D/7iIDyAhqQYt99dxQ6W/O61lYJqnwLOjvreW0+fTFY+zxDTUm29zZgTabjLv6hnPJuk+B
eP+UkSy2ioJSZg3XiAPQJvOQOSqNrNlSRd7kMd+QBogihcvByh/NvSfU+2G4OhSFxubp6x2Nw6lo
cCvG1ue4h/7ev9ttTbXnoYj53rwK4UoICzAZy0so26Vcc2wyLg4jYlwt4zH94b+BacMdtA+PhooD
+tbi8uNGAP7VvZi+ZXUCfui7MZlMNrjSGv2GbHUnVhcCDMsfZ0oTJVOMzXevJI7tG+Pthrvr+pvC
qF697W9/J2sxzKW4o9iE1qmCj0dFulbtnF7JPQqk7HLPy1bovg6HO6lnU7gG2y4jIhbNEdlt4eiN
eUBR/sS0+wGlXlNC+KpBUQsapXFY55uMG1tbwFk0TlNAg0/aWIGp9tNH28n4ZrUTQDS81te7le+U
KNhTb6srCvsChAr1eM2P6U0iYmE7sRzI5wfolIdVE/6736ED6pziqP9qqehX0yfb4/DmoFMIRv7f
KNpDNkHSfO8UpCw//jYZHaaCdMgjMhPsyhv0luK9MLRGEljUbd5H2IttRnlOyu27el5X0EdQeeYi
RnorjPOWi90jzo11W/AY8QjS8HbgQVRfaUPwTHFl139dkzOYX/M9jskiaHkSxRzOPWkcY86STNmk
8OS3jv5BWVtGHFwhsa11EnqIKHtHeJADveNE7fCMkcLPUnfneFuJFajbyxU/J5bALTF2Mjj6+KGj
VsaAjs3I5E3jGrLxmgfGHa72PcFY0rd5eONkIjn9+Nh9gjrH8HTXS7nk1Px+T0ytVsja8MKZSv2I
/heFq3UgFLtLvm+6LKnBvAF7TTWfgM4z89CMR5qyGrVWKbd1rnjURoYVPKXIYV7nJ3qbo1eCVajB
mTwuWxQ3EsYb8j7Hwm6Y98Gje+CSAvuVsfvD46n0RiCAgA7ON5nDoy5mz9kQTr+H9Vw+LFF3hNo2
1B8MEjyE1SEZIXDArwMPIz8qEPeId7bFHbaBPYnVZZrYa3jpXDH4PUMtHaEOCmMONNshGLXzF40H
UyUWUIIuqYmcpZMOzCJoYLmGiuYygI1QIThu6XmF16xhlm7Tqzok0Vs+voyHpqrb3BNlhaW9sOzc
Q808XtrL2JIPSrqDirTHaj7bVH+vZNx7QHLBATPMGdRjFkHHNJ51fT+JpwWD5zcVA1hFyYS9scyS
sbmNb1+X3uoWr7Q4FnIy7h+5a39dNvEOPJYQPrPmpeRNtrLJCv8Knvidkn3qgMf3f2lODjPMaRvV
IXtSGrT9UNziMpGjTpYW8CPXCM4ZWmPljJ6qYPwQueDmMQgOKCAqIQxAA+BxPgkHmEoqUvxoPWG3
El7uUNgJzBdeStLQAhrgDP33ChMdtGYcYAAdx8MV2NFVSeodjLpxj/tVhAwR4HiJbYEYYyOpGXft
w6FS9ZObdFlVdBxRHvsZAAAa2g+vNDQEYtcSNwYlzbqEPFuA+rCl/FQ2gp6p3ZVX8t6AZZJI2KNX
nFg9WnX8aSx4Y7UmWgrHxdiBWb6rOcYZLK2KdBcuuNd9nqPoazzy58ZXBsBrQF4hQMTxunfjSpj5
MOq0i9pSo6XbRDstFFS9FjX1za3Z/xaR1T0gYL16OTY4mxOiju44qf25PsH0me9jrNrnlJ0CECyC
bLzoHixhGPjQujXtJ/CmOB1RWnqBWroLXbcHt2Jq8a1F0AbHCiAJVsuKhcd93V1D2+o4Dcw90vir
Uo/O9Cnx07YCaAGgtK+QxYpo7C3/4GhgxQNavqN7ZW/6ruGCxngHpxtMjL49xNoUNi89sP8+w7w3
+s+Xv4dmptfiMDJZIV3tH7/x0UMCg4Z08EfE7DCq6ZEpso2HsGobE2bade0UjuiZcEDoVTqhVMbU
ChM400D52T2ECFkhducw6shuBzGNKUD6XMC6UgUzCQPMFQZ4V+z4rYek97Wwx2CtWyyDNCt8qmvi
Kw6UApZe0XPaFlUz/E3jBFzzogoKBVXY9nWfwMNSKuBWKHUCc8baPmxsnK+LhEesrOvGUvA3xe90
GnSTRm34coth4emVH59IsqAn9o4FnYYQ2B+ZMlc/Pxtj3xSmmouhGKlPjwW9sKj/EDAVkpmUcLY7
g5Nfx+jeq8yV/m9+KWq+qAjmO/8wz/zUyOi1HZStNkm8rBreboxEUMyothmhd7z9ayQxuGBzKiIQ
npRBhN0GBCtLVMw8KvAfi3f+GtrVE9UYGxIBpDGsGpCloKcuNK/iaOJs7KGyWTFo50bmwuStygfs
NqEYleI4aqAD0Umn/P3YtJgKY/HlNErI/dyN+gtyvY4jfMDoaQRsOQXKPyXpkxKGbPZB8V65olWs
yX9Ewvsd6EU0BfQovEYPLzicLwypEvBknL7jqjEnl3wp7sRXR3nBhZcprxwqvIbsjmrerVwbxfDF
ozgJ5T+xEk9++/sB5dRQw4vDOZQ4CoaoBTqbS0vuUESe4X384huiJfFgH0l8umjB6jDkDXQLwaw6
ue/Wz10YemCZA5ZaXvcOVSvpMesfSpwb/jmZPwb0pwQA5gbdI1pwe3+AivwCohxJFYRgmywyGXFb
65hmoE+QVX8AYe7pbJ0YjzliaiAXnMrgtobPcV9mlIoOCkq+J+fSSgpsOboJ2Y6t3ZewRz284z//
+ZEelroEPUTKo6TjwGezJhiAXRTZ6iJKzEc4VJCE8zIoW+fCajQt7xhcUrvXPCcYKWIZ/GzedBJ7
ozt3m7MCQ47m3DY45shs7TqKR7XRp+afrhzxzzqyFthqX0HHNs+Dus6d1UlqpjpGju4MEX9nD0Mi
9cpGX7fopEDc2J5IscdKXUHFZe471mrcNLK4vrhNV9aNSrKZVJtHSL7KWdiVVnzcxlcWwPjEPiTD
4hgPmEoOXoay/+XOYIARcA2uW3wqRaGTMwHmh+cueUiLHOvdnlM8ocQ77nc/GVJmcQLYSVRxi5J5
mrWoO+yAFPFweRXxvUPd5xdtmOvwmUsjuo2tB2Hrp6YXmzGpfSbF19PmxMuLwvwARz9og71IU53v
zozkKN1nZRBgGHbFjDby2w47kdlGJBJAq58Wqu1Yeoa/MB4OMtBjQtQio2oMirmrVmaRmH6YkxyT
GjZpCslD9xPVOGVVy0CkmC7oBn3+HwgMvjGRL9tv7qOBC+bjOZXvxa4LmDO5/pPfPDk1vVe46otZ
qtoc5FDXo9tjEeg5423T3faoe+kzJ+VwbMa8odDN+ohzr3G2T25wrU2eRmTjBwNDSDHdODNPY9Z2
jP897CPwPfYFJ/2wXMw6fYEKKnHkvkVZOKQKjfTlhpQ4Hvfb0thHDCTXl9KEu7+/S0Lc5DJz8tuN
M4gXeZChgwgVBr0IEAALlXaK3wahZrbl+tUjeAreTNaim3cTzlBW54zmE7RPhtmCk1kV5M/kcQ4H
w3h1IUw1hzmSVxaxchRkqFq97v/79AZEd7FjrKcvzhX/VAw/uKGkOHeLFn/08TBFAdenuSjZ5Fi1
6Zcr6VUMSsmkRuLMtF0tqjhHXsEBCxHIRrVGvBOab/LXy40YXfKmTNWh1EyV9pvmSVJci+CRwyZj
EHnVBaybD37QW1QCony9BJyPvmpJ+EiEXp57z7fOYt4JtotKteC8Wz74Li1gQ+nrd24KKUPzYMPH
ye5p67KJp/CqFt9I3eP4LSkNOknGKR5vJELuIdt+vZCPnJ+5j0f5x3FF7EwGvetlodj6K4Yg6PF3
wif+/sA6/aI36avgI5P/mDWAZhNxGw4IRdB4bHW3j2whg1bSrHYALwb/PLWdOCQzFxAquq3bv4bV
o0o0UUsabfjq+leAFDqRYKpM+yKNNOdwOj057upuuIMR21EfdF8YBen7tsAGSZ8t7v06cxCFbLZD
ardlrpgxTZ9NsmfpxZQpNchsNpiZUjKQ8gILiWxz7CMgHIu55H4awF+VBjK7T3eqFb6HgjggfSLF
kPijnqucw5gRTwG6oRsimPRaG3sOZVJOvNNPDXHV2ddg/rIRRfVbNi2jwgqhhbD+6iXNNsybVDWm
egnCTPN8C/ZACWsege7JDeB/yQflF3fPpsnkvTVfA2eKSvzjHWOi+6HuBgUx6nna9EqCozCXteaF
PizjplOg4I4BS8ulJFR1q1fjyJkVJbe0sTkFzYAUDkuMdNlL3Pc0aYBvXNxHWiXPOjBkWY9SgbSA
suvoTLVN7HBJDGAzw6r5xRpWPgWEH6LnIZ8KM6XXSBMkbK8be7YqRdqKKIk4SPH06cLSuBR5Wk/O
WaopcDD9ww1A9TuTfmuS3qc0LJvHfza8iVM+64/rkYzy3ZtQLTdO8Olr8pgGWJxPXJ2o+i69eLrT
G6jVIB8ENTdVsH9t19YYE3N7c/95xGDkXyWhQEZJdhSr81u11Dw+s2IRe1BxoWBjBqIDLwKeE7T5
qjmwwhG4xQzJLE45Tqk7RBO80FMwMJ7R46o/hCsLfqGg/TUQ4ivKpLMNPCAcvIuJmrQBZ0eu1Zxg
akgdgJut5f6T0BGWWTurnjeYmO6vg0VLndMOyCVnkAizz1B+jBHC21aP2PNfmjONkIgX6D/oOZyf
0m/Hu5mr75nEqRwowOuFIaf8fsPewzo44hrqGyzKQo6dsdadnplfi5iTMBp6KqzQehwG/Qmck9ZF
ZpKW87CIikXe87w6H7HKraZhNCIe9SSL4GV5FrQvv4wFy9d8l0Iw/gso7tG3nyyp5Q2DhqEhCTFa
DS6Fftfw9054FN1XnKIewFInOUCBjcVhi78BxkG4kTjQaPAWVf7vth6Xy6zJIp5Yktk9R9WiOngP
9d+Txam40o/IIozgYwKpfSj6WERt/GVVWfsifPogEMNcW5h53S9cB+CloIH0a6CHpWPZ3I1HF4bc
/gFqHuRN8rsWmnb1YdEcrP+CyJhr94kZFIQEbsUozqTJ7fmBymn3Rb62EVo5f5L3Bt4mG6r8YrnY
gIbGv5XA/gqE8+AmWPd3xMSkUlibyDTsph8xjjxb3ipQnsJnDrLVmj9262PdGuNoYcF/zVABnsQE
hnLdp3U8RbC1CfjODTkx3x8EXaYBJtnDveLRNMZ7Lsb0n1fLV4vhMnBnAP8HThiWwRCL5pbaib29
/XAlech6CdnWoByJ7FATyY936Ez/KZksRhNwbwE5KZEWGvJvwCp9JnPDq/vJUOmJCuubuLAPKeiK
TxqspOOHj/PhRt1J40tFrrgsUKtVo2Ue+ZeMgFkzcbd1EknLFEIKEBoe1X0YvZ7q8UiXVQTUusL7
plxeiNfrs5rjxyxAxFRFFQXDoZTjwjvmKJ23V1miwczBxMZMwKslpjGA2g3BGQvCeVVpEngdl/51
dHUmBkxaf/Z36RY8hiCtOwAOSfb/8yaE9SKh9J8TGBs9z18cgluwcwSCvZnu4Bc6yh/Q8JL3Ntlo
wya2KWnAId3Ek/xs8kkGEkAnC1YasErfwAdGWcur5ugjx/c9hZe/tsFWvJXKjwRUyIOE55ELc6Qb
nxSNJgjbJSnouBh249fGgaVjM/h58gujnjk8p6+vNl8cuv+z8tIVOuYoIdZH9ae9M2glx3RGXmDJ
xic5IdMrjwhSOtF5/fAbRz/uQgjPOsoehD9gPhELTRT4pfujTbi7QmiQacYWWGrxY0w9TN+SV/+A
0wUt0c6x87jCrrn1Rh8gkce30xxysk37gbv10nCKJEJ3YsFW0fmp+pnVuLyFVpw5Cov+H5NqMtcm
sATqwg84XY2+V5iVW6OEJvx3ppr+nhAQQFCmbM1tZw7YEcIxzcoFSxqn+pacV/+WsKcqE8Fv831o
5FxkmUHyXhZFLQnc0aOtIy78jRZrdQWI9Gn5iWlF5hz5LKG/dN3ozMCuf8wc/Wza3nDQBpn23ev/
TBnynhZ3NAY2J/dLvquyBuuB77wyop5andJWijSWb/euDLujSfHBhFyS5h5VoLbttm6mK//Svg7l
CczFKres0aeIxEfZjOMUifkjiRCnVEkeci62QYCgjszUlBChTDRPoD2WhcWv/SLJRJ1dqy4RBKRr
aF7zAK015aUq4uVs8jU9pGIZw6TsN84wQS4JiyOAkk2apJuujbmiX3LRYHe07NfSp37uGDvAYjB3
59W90ngmnjLLc2buZwKzqtmDIwUu7RL1ixQdIIvQGoUCyi2kY+la284PP7RK0rXkxdllV8fgAMiJ
GGsMYKiFOUaRGE7BH20sgTLAxuc82sV1KyJgL1u+PEt2l50Rl0MZVY1B2r9hnLtG30wpiuMxYQwM
KgC6Qvxj/pwJwNvOKxRdd1xW67uFYMEiWXtVjCH+75LWckPGHEyDFZeN8WX4QI9cZYwsVLug801O
1U3lzn66gU+CroKU9wKYOUFcW2co33IMzcIryBe5Pbst5ONEkuOM3efWza4bCZyJ8DR7B/hkrM6S
L22VxrlXPufZcsuDhO2plv3NvKA+MRtuuujL8XM6dziVoolQoSIGPbev1NwiMZjxeXIJUVHBWNG8
RmQ3ecne2XNFhGEF5tOA7FAP5QsFBocAg+1HS9+4S531pbekCamyzC21lJ1+VVloPuqix9cwpJ6D
/OnhcTtEfmLOH7SeMdhuPgH7bobkDJRxnI2xpbcwp79+keaAB5NQrEMzn7BgHNWfRUSCVjdneUwu
g0VfFi1/G5HgdaIipFOHiEFZoKt29j4nB/Jb7RpVwR0A+PMhZbhYtw4S5LCXe9F2lbjruwKl4Z3q
AjiX+HtS/BI2x1cnCvXEaCycb+VYnH9LqjlPMZcOI4MuES3l8QArF4VEJUIqjlh7z/k7PXacK31b
Kmc5LwK4sYLyOkUpijMnG6HHQpCfcSSeamEb+lu8Sq347+bfFhqJ3jjgniXkuytR71yDyoQjmF9c
oix0P8DgeN0XlMu0xAzrnle38WPVPsWoBcuwv9xKcf2zppwCaUSwnDAeM0b/8KIb0HS0tiFMr57D
WyAF2oTlOUb83BxnKq4O9ozeqVe/zLvdFOSo4a3qLcdGF27jouXnDZilm2NFa+0gdFrom19i5oKe
y+Cpvgm8Fxv4MVqf9F0jlDWewEnt7dXJBZrGmXs/DguvUkNZfKuBolOLMLoWrzSuUzv92y5YfwHQ
KifXWX5x558/717PVb/2ZSKrxahGyn9Wn9tArC/ID4AROAaqmzcZSYV9lCpBfo+Q1z0syQtZ1S/p
mkQ3k2JX6jxqC4AuRcojYNA/2FyC6JT3Mc10YCZFetjcrzaUw5yBCClhtKOVvWRhr9zK5vBeBnyz
e6McakcPYu/eY+U1LuVXeUvpPIyA0D+e5wtwrmRwDgnMV7tIJmEbYpW7VYnR+PdU/yRsF6dcVgEh
8L9B28N5QaGaAGKh8/22LzF0lCe2AhJpo7siqDF5Qy506iRP/alhn1fu9XGG4FrQ1W+XqFVCM7fi
WW/UzwG95ZwPcYnifEMwgjSX5ru5sZy8NixcdqUMnpQvclVsKUdGndFvqTtzeRWOAk7xEhBojw5Y
M6gWxLrQXn3MBABfe2PLv2BnawQ7EIobm+uwRULtMNmPfbg22s53It6nxU0Sulhb5NwLTg7DnSPf
NdU0DZMzF3NqOZQx2VmrdsUqHU7tdO3PuGAk9l/pgo/pO7jqg8W667w+Yeo2xxMUjIhPuQIB3eGU
0Yvfvw/EMqnqGN/9wENm4A0djN8u/K25F0JS2aMNZdOE55+uIq3T3Owt4QTG8nOYEgUnlDcbbt4b
/Sjy+lfwtUjrskbxwcpGjfVdFW/l5QlvGPmlJjBVewKv5zw4VQhQujFJTBqXfY0dV34QfEGyed2q
3pzOX4S7bhaWRCl7dEwvWkIdVMmyOdbJfrw6RZaVNXlWNe9MDIvyzx7z7nJObYBrC052yrNVHx+w
khz0yiz3aNGM2fTMMbmAC/aH47VMcaBYQf6DXQHZdwnuW3W9kShKKuj2mMjzn3/nzn8/VcUtHaQD
qZlwbuO/apBjagBZF437nhF6FE5NJlko1NyOe4ubNTFiAPihqJnHE04lCYR3cvpLWQyqoxPrF9Jl
XLvCPHk02DChd9fh7il8DHYY4OcmkBLMyA7nIwPWjs4TCyzBo4OJQnOeRsQrQVnoR9yTI3d5Mq52
DC4TwIqjrylRzQTRpjDLKICBLpkBioVE41GKDfGyEARgk7R0Ljb1UxBbegB7MsVoE3v885N3a71T
UVAFcBjCHYOdk/YXWkX3x70WK6aBv9OJsVntv2nX12DqH8NyZJcGYyGPi3hoFiDBdCUYRaWl1eD2
pCR3s3sbVJ+wva55z24ChkDGvf78HwcEpZYEXIrtj1CVBQNUoQGyS95Tf6prUVfb9bwZSqacGHte
ClZ0xgy6PrImKGQJW0Wd8AOC+FvkQazAKp6H9RKZY9RvjqHfKHujllzl/o8TbtYxfCITwwjusnKC
ophmEABTBLl4oD+xcswM4oWXEtV9Xjkf/Ndg+ZEPTdHHaLmpelbdvz7qFM4Ewln6Gc9lB9CA3MiF
i7k53BJrh2NDHYB0CVO7ZQZ3Q+H4FMKI+yD4UZuIlji8afqQnjj4DNeM+Epn8r4liwCBYWfUXRuX
95pOE7NvZSSGgioYkaSPlwKDvbDTTG9aHFrcG5VGugPv/bunoLgd1xDsySf/fSJcbvM4FLNPTwTn
8u0E/po3YLJpZxyMMIWfvZ9v6xyZ/4/IEKEouy+CyVOUZgPUoMW61F+9kuMLFJwLEhLh1AHGL12D
LH6uRwzWkZ+VLBI+SLCqfeFvvoPURqE+W4NsW5CfGFvd73k80+FpO5T9WVGJTZhNI7h2TWpIp7J3
7ouV1wfMR+YwKn3pLEtn3YlMOLIyyXfUmESs0V+aIniCwPgtotLmNdNTN4x0Wj9227iDbVgt9vGG
mEOqDLdd24L94BFjq5YbZdq6MLvPcdvYtW3V1APgTHhJW3sUEFTrBTCn00IxzCj7tHYYyqZd5l74
Fm4YrHUl5es3hTq0aI+FZpCtRe3hJ834JMS0tiNuB7nHG1nt3V0/eyATzJtv0MIBh8glg+uBh93S
kngPrYJjibCd0ZJ89UYre22sMXmm1BP6pTTNss5GWmV5KMgIYV5yOmrwvkCN90HkHLW7jGP0RZ6G
2q5OfJWi4hwwiaLCcuxUxTjDuY/WVQ/tG6/8N5N4Bc3PHSKNbSNjaBbdwaflmGBuOCbAiRT4yU1Q
Dprn29DbkcHF7SwP+EcxsYD/zWDxYX7JSI+HriIvPOZWep0yqQL/jI8f9J4h2YJpkh36XU0zzTEt
KmX15msZler4SGBtwqSpxsW0ZX5aybb+nOhiV1ERZq2vcAd9esFaq+hAmzGXDqmigOhyhh679gH/
kU/ZBCnOVXRzwIBb/rTsCWGqAOH3KIW6TNc08VyjYeXxKrujC/cpXi8h7hykuaUXr2dBSg8sAvmx
8YRYdJfs+9minSqTY+GTtl+ACkJ+U6qKAtxQPmS2LNfojrWxNOd5whBdnnYnhhPu481zvOVrv85c
DdFRN90Xl/4GlSa8UsiceKKlkULUYjq4l9/wW74H14s0UqIh3iExzWz18I/lau+FkY8NcJ02irB1
xFAb2ZkbT1T4qF4zsEq0uG3YrnG4hJsnTh3atgo03s7gXRAM/ky4j1fBh5dg7hy5bMRZd6dg4HCg
F2Vf+R2cL6tDX8XkRU7gHk2YWggu7ptosyF0Al+MUP1QSOH77Jc7cc5mM8kMkV9vNpHHLAHJ+Y8R
dA5AfrQaD046qlSIICNnomIh9FY2LN5m4O031RnA54EWNQ7nNyaHpnJgnVzDvGi5pER6xsMSaTJB
VL4tkTSe4fAzfi2oIcM7zGjNVZzyWzW97ADw9Ha8oBRJVZBKWJ4rG+KZnOxtOBe0CGLjhoqJfsvC
NBZqvWWeOv56oqLdzXgWpoUnFCF7kxTfIkTmEBKjzWzDLqN3EfBayr92vC9fZJfoNGRrjUvz/4tv
VGsDiVYrXaSOGF2OhGAI4WxE7FgSvwkjJxNGgVSAj3nleM/X2TgDy2/Nci1jdULJPUps3pDllo7C
Tr/9x5j/b+VLNAVLMhQ35HGyS7UymnErk53nEbRYXU4FQWbLj2JvCX3+dD6aXogbNLQgRo9PZ9sj
6J1tVv+MYvxAhlr21f0UHZKwbGzGAQTltCSe2LTzsjfM3IpjsZOcf3EuJvavlgMxkJB857lQ/2wu
bfjrN6xQiQCOLS5uyjGGJKoC8FQ68LuPnAWKwzAeJ9RuTTxOhOJhXs7o3aMlOrJiqTkrIlXpuNon
pQ8Qgsgjfm7YQpaDfbBc2Ruv7ZYe8Z2dEFI+wQ6xQDjOMdoWugLegAX+KS7yEy0PWzpBWI9mrwFH
didPW7TseWiB3w9AUtp5q+xPlk415Fn9a7jB43bD6zyt13ETERcGFNh3+le18+ETaLpxlAsoZamG
jDdTlnibkCqUrHR+yUE80Goj9lbkeZL6jsc7/dYQYD8Ccr7ihiIi3IsIMTurLoSW9mIeAkfIbrcd
365vZH/qM7PeobUhyNFEJPuBMX4r/vwVophvKlJQm7YNlC3SeA9J/eE6agX9Cvm0EVDSwMXQ0TEh
WJ8uIquCPteLGlKpu0oDNhqXV3/jIHJkOy6KeIfDstB3SCjpS+G2/kDkuj2voUA1EooO1TASfgaZ
/SGk4ZKY0Xsa/D8wvnpx97iwlmekZ8u9BETFf5DWLSwdPN/u62NSfb6ZX1+bqZgVH3y78ZwdxIID
nPiQWTI2cc4Vk5YqitaeurtzDTQv2Oq6MpmcGnyYmF68cNQmVYHqA3iCw/PfqO6IVZ4D/dQ0WG+z
Yjj+gtIUIihu6IDQm9Xe/RGMrUojTHwIbV1ZleCc1+djBugyhuPNxMVcNA1OJwArHD9iHsp64vEf
dJw2C/uOkHNtZZXgcpll4bsOv24yMHCAbCA9v7X+iobbs2xn4z0FQyAenH+uknSaEAZUoL+Nkadp
WWJ+yQsCp/PcbSPIk+j8MjBasxf1Wmt7IXQXKoX2w4IMTsbO902BZHCaIAZg9eGQVefpSgvLSQjN
GZJNsuHN8/72cTiCTPGNKNUREO/qIPCBCGL2ezFjJG6xZrbQLHBH20sfsoV4685xeuvKLnblsdhU
JU6Z18WGO3l6/7dlFXc1AYQupdjMcebCGF+0dxpMGWP+rz97AsptaDr4JgjNjUyQlDPOV+510p70
qGsHv+B/vYXxt05dX3N6uZbahflrC58uRzHQi5U2TA1yXAz0D61wQQV6fwe+CAH41gI8VQeO7jAH
2/JSRpZ/+mtaGgjPqRZtDTN+iJ/7Jtnff6vnre1EZwXkg/r6qS3fefWClNYUbjWFCvmDA3y+KWxe
lgjW2YD6/Zacu5j3tMOfLzRQgyhuu3T+eKNZ6YtL6ZXIL+c8V14WfKmxLrxMEFMKYMc6n2rAFXxu
ZE7+o6XQDfhiUPNtFTLUaJ7lSVwek9H5s/MQdcg1GU97n9cb2qnjRS1ezMN4jcoUG6Jgk875Y52r
idZxsqks06Yt38S2uojvkxRj8QN1jIUEIyDghinQE1Yni0afuR7lk/5K41bj3dNUsFXzDcWcNUUL
vvMSfbrKUvtsZpJq+giFrqhIapUQbc8opDEo6uU8EqH9ODVTmmrQcf52hY36x3pgxRu7PEtXK0za
X7TUck0+NbbXI4Q4CBTR7PLzYKpgqaVHWwIq1nLel+IAL69YmnTY+KSBzI8dAcmE/gSnZulhvGmy
67PPjEbKz0aTEaJW/cbetx3rEWXTjevDTu5GThi8TPzrayZMNJAtWQgCRV5RMhlTHP0Lrr2AJL5m
Cn0vNofKjHFd6Rq+tHrgfF+Vn+M60+Byu7oXyO9c24UjFldWZURtHMSbbuy8AhsT3IiOydVUyj8U
n0dPh8o5HezvmW7gTZ/xPr1GOhEfaFhDCNrMJArP1eZ9Xt5sgmtCfhiVD9GJNMBe1+ONciYtxfs1
AlAfxlGnJaYo8xpfNLYh2IxXcTc7g+RdKY0D8DY8b1EknFyoYnrNYsDzD7kaxeXUMNtumA850WMI
AelppkwNqvJ7/+4WLH2ue9BMiQ6c1PIvvI9Z+yknlnZocipVQF8d2ALuCHbXX/IlxLMp42jj/5mr
egPbxRukE+GNQMxlBmMDH3585u6ISqkkFKkF7xwFa3VIyLrAzA2jyDMJLB1uFW/HpojoqdS3ba8K
rRgRgEcFRTjX9jFqbu5SwSB5jidqOQ7m3li3R22+o5h9yqQ27gWNzvn8/niw+KLrZTw7NGE9SMFG
XcauqoAIIiuvS+fHaFvOyioo9aSe+rEJ4ZH1YazOjyCpie3OACPCyHZewqWmSckgBlxOTPZDJBfj
Z1jbEdMwoTkz5NEGOHupkLg6WeqbpyC9OBAiriUHAVO1W62lRN88JEuhzQwTn37yfXTIDE5SmKAr
nsYf32KQrjasftR2s3iE/KWEHwJqByMpDpYyICqxJxrTJj0SS9tFy7Qczc6R+Y778ugTxkk+Dy2c
/2x+b8hqLHxhATtGB7unnLQgR21FMhYaRFFK7FY68NmfLuqLKXKM1dqkR1ep1jlgVVRjSM9l8CFs
bTlDFAOipGoxnaXPApMybIUM8gX7NV3MZ5fjkgPjzpqgr5FXWXBlwfOEPr7uWihBlAgOGvVdNIst
Bu1GZQUITFCGs/k2Zxc+fgUMxtT/SIz90fH/xWm4HiO5UbLrGXBqOJXf0kNTiSsNPz+KkDZ0KXkK
Cr22xnDRED5wa1ulWvkRGnHVix4n2hii9riObPQ3CNUr5ykugOEAqQfGi0R28VqH2rRSBTP5Y6KG
kKTGAhkaoJLMatwsWyw4iCmLwZzxRxrTCh5u/HoBdX+HbXFK6a/0TSerU09I2lW/ZQS5U2OG/RK9
zTBg/EkozDiyYtXnJjIEi4tTKf2DDX66NVP5Ev7GMOFRK4Xntb7ocuor3fBzRo6s+7HaOigSSPZk
JWuY4g0OvIfDx9iheUMMXJn4X9nfkPOb6H/w/F45gNmO5M6AG3Js5JCYriZMudd0n/jsNsX+wzgT
eUy4nqiH9Ht7Wzk3m8KWA68z3xQCXWcUbbvd+s34dOQcG4UcMKatl+TD28hAe7yv4cC1xdwi30OW
OuA8MIo9ILBw3viGIqPL7B2no2lPMM4A0owPgrT9PYEEmOwqNaGghPukEO5ZY8ZLssDU2fHVXsNd
GiumWhiazh8ZjyXSNwWLzABEVB4luRhTGre00GaBLUcKRfHZDPfuoGagWgA94SG77Gsy3Xwajqae
FJ8tcRDcOmdpWmQX0wn4Wd4Q8MCwV7xk4fpJ0eoSbPSkErotUock53zGd3G2V4+Pk5gFGMYDHH8P
7Ab4vB85E3FxA7VH890tFV9X3txM4C2czmfOleOX5mJ09HEXmvviB27oAsyo6k3i+jGrXmeoC2Rc
Nav5mYm/vuIpBt+tVXnQ6hsTPHUpFXv2uGDsbvtxO22FCb1NFkT8dHJpBt+Cy0EAy6t1uAlwH7C5
ZkkGhJl4jh8jt8fUnexuQRZM6S6tavE5gfOBqorc80ql5fZf/cJnvNIdTQxTJUCl0j7wJP1KsUO3
Hro3NTmWTjSP+J6sUorWQt+st7BkLJzrqbdN2DGj3+J6bO/HhoBUDR+c2rBskj0qG4AxT0HoHIit
+0ehltVeGgI9FhUmTy0mHRRGnPYv5X8sqXLHUdjNtQ8qrpwwOpQWcbA8QXCH0FMdxGTMlJNuOIeD
e1lheLKlRzZyJbXmIMFZT1BfkREUWJv5W2WqzbVl8+0yQYkbST5cCo/kuXiKTJxYniwyPd337ImC
OI+u2wR3f8bDRLx79VRv0L36lEdyr5LpKzK/S9DdS7CA8+aH1TTIxNlvYJgoTBesmvBy//SHDl1A
CA9+qZDdy7MwYBLfHA96ifMJHtFZCsgjBeiYOGtSa4imu3sGjAB4O1mQ+0A8TK6oWEKBHplA/BFu
s23yhddWmIpcnuqTehtIjW6hajcWRdA+ggTebn6BCEWpGNrH4xX1QiQNfYt6qjoJ8OwsBqH6KmOU
csV1X00XfwTZVZkfYnIWminTYBTM1Ii8d1nLxeoOa+hFu3U1XJDfJtrVrMn41lnLLYmMVRA8CYGR
yn0Y2L6Xayg5MwBPxx0973AqallGPuGr3eMNQhLI8848xK/wGY6RqEU8pWbzpnBymtxjUJbYRYuN
VeIr5uqWNuiqWmsgs0T1btnx/4Cz49Yt2oisv5/s8OtFoPYxU5mgqVUPqob0qOxoGmwDv7ObMXB9
vE37fPLqwHbpbAAlCYnbR+r5nP459iqEZEn0bfFD5I9W28vfjulyN3fr46r6ZQxmb3kH/inIOGKA
X4dui3QVyEI/P9RMQa1r4BO1rexQaY4sDWQLmvbM2DeM4oU+q1z6GiMouUMbRpgUJFsFKSPdesg6
5XEQajyd9998J4qRcMWp1+lJC8HYuS32iIrsiFL+GXilwxA/liNErzPF/sa9jgumU42dgL/t2VzM
avtfs6iybTT5joOALNryXGXDZ78vvEKNBbcMstr+UBGAgpJPCREOxqaEnodsVknPYyNlRA10ybxr
xP1rUoCFGtsAUg4mhYwOgeEiFDoPll+i4fgQB2TJgCdBpKEGYints53zRCNfbPt03HasHw7xFvd2
ejVF7JinOEtXyI4erVfD0x2HzhBqw7d6/euI9gs8NBVPt/QKjKjAOgx6aA7aJCVIQFwnLM8noCgi
RzTOJjn4lObTamSzZjUvv/7HBhJ67abPDCiHZa+vLqXxyKlZQUBq/D2kdMhOxE2iUSRg5Es2fCiy
NV35JfXmg3jwYv6B1NSFyc0hrLDF5iI4DyJKFn4qDFCxiKivG+5nzFx37tOKb7llUvSpE1Q3r+IA
rs0zDKP8llrWOm1Rdxp1EoJ8X28nwOEB1ijTWxsghl0znzOOmB5YZsYKVTYYbNNmDgThZDHKQrQw
2L9vuAmgDcoR2V85d9WkwYlPt2et7Menn0XtNeB6Dab7x3D5lLkISf04SfezuOU4s3BvbZi55PV6
NyJDAwzizFWgczTLBD8rtM+VpLDtUEcfFEQK0lYGWLp5gfyDbkPIQ9TMOTvqKkpnUCm1a/E6mICO
/Hv0v7UsSNhghrhq97N4XaIcBTzr95aV2tUrb2o6i4lczdZc5VsXsVd+lGBWqoHD3oZpEURQiPSr
x3vi/K7u7c16pA0Ignj78f4zqhG2Ljj+8Te8d6X/uTD6/JL2Wl1SMWjH+nF3QJJevhbkOYu6Uf4S
nMA/WQm1rc0j4RgecXoCb5FoMsefwZzrMVDI3W54pgKXAEP7Uzi0N9ryn2SrVwkeruCbxXgHBUnm
zjuF80VvCyGcaoZV+Ca/3lxKR7VyrMsJGpZATe3pI4atBDwuL/OHN6+YO73/k4Y90Z9Fbkejwy+W
MMGSUrOepqo3k1T0XRkbAeL80Gl989lY6HDPjbAjZYYUIBIiW6I5FJfeLAm0GutmizAGhpKStQnb
iPGNZZ2Q72YYKO7LKug1W2gkPXZfOn1J1vHQaF5QBLH8HptxsusaK4l2qEr8hvXzaE7uq5ajB79W
i1H7asi/C2mgttSVRIp7dnd8Lmy3vLXY3SPadQ/cRTdIug4z/TOeMSQLMbdvhrQtVT4+U2hTNwuI
Z1NP941y1nlmdXhItNcCLwMZXSFzQTHKj4VRpb8NpVhunOhPSDQYuOiBtN3hN/7lFa3683XkHxe4
5iLueOpQuKI9YhbTXYg08A+4F9qqvbK+uwqVJmMr0Zjc5ngmdYhH8R92riQdfeETJ6Zwof3dIT3U
WzgKNtccwJ5QhjpJssT765cq+iBFooKzlsGwcUc8ERzqDg/UsUgoEo0UD++tqFPHe4ON3zeOvJkq
iIdR3QUQQ4W0Q7i23y0tKpu2dRUsN+BtK1C0Hnv77vba8BB0ZhBImr0pNjQPfz4ZHZ/oq3cszBZU
LGeNxoNQhdiJI4zzuT62RzHES71PaKYplMm6QwcUB/EFRsu14e5tTzW6s/BIWOzA9369HAFPWZpt
wZ1ViMIC762rHr5WDbEh4FHcE/1qt5JOD7NyxJj7ARflZD4i+kKimNvCLmwQAa3q9EXZYKpGHuZW
LtyrStjRp2IMzVTnJBhW3BRx/sn+f5z5HGbMIB6aTQN9LezItHXlYUjodVOjZXf5pGSxfIvRdh4Y
aGeiftthy5ezRkMNieLYWmZALjSe49Eq+Tp5ild3kucqgBa9W2vU8UUUrFiX0LLwLowprR3amT6z
nOBkctf9wRIeJnazqfelZeVQMAtUkaa6BT2AgwFrAxmgo/rXjSnrRFXDdLR24UxfrjJ0T+IcJGfW
sbQ0Ep4Bcy2e8KFUcZH5H6zemOs3e0CEHGdDlWcHYMI+Xhm4sJozeYJG6AF16gpyNBaHBSLRtJEu
IFIw6gkHXQu5dItHQ0HtzpiKpoZ+vOvUAi6VhpJsdlfYfMCs07adZrvcMq446IhoA2y7V6VFO4YN
WkIGkAxBDZX9/EmZF5lIDZz7S/os503bI1xCfW1iCSmBYeP3y45JdZFleIbtZku7a01w2vZybcBj
SKA9sLYuZGgEqTrkpof7uWcWXS72OkGG24e2vhFGgJZSdvf/3ayn0q97NUaZmyF8GhY2JazKpigo
7GJq8rfPeJdyw86GwjNXPECi0k7+118OJCireWxe8Sf2cf5fHRkBvwuaBvUZLaF35dC+p3m8iM0V
YabfbyvG3xBy7S/I5HsZuZTf9FtSsBrK6uthofsXkbXnan+aGs42sdPMAZnpuXgPM/IviLq2ZSbp
ToHkckTUv1+e3LpiU+xIDrBCn3qZjH97py5F8kZ5Q/Hjxsu2a5HwasBgSz+yp3i7pb3rO8F0DyCG
tACYqqLxjBPh3PEdG1KJuN6QPQ9MeBzRk11cizcSeCNzOXcovKLK6HXN+sbCEwB3Ne/kKgVSmzIi
AygEmzuxY9WmuLQljtTq/PRP/KyPvKOsJL7fPNBjoH0iavNrrP2P8zsa2RnTOhtIRQWhAzosFTk/
dlA8+tjcPEJBTatkBXOT0dWHBMK59mod9ry79MsZ4bq3bCG+mDFl1Oga3L0240fhTCynUDLhxDdh
9IBo3fJdPahiEmQaDs5/relEt/1Wtwa31hagZ7aCL6ZoTI6OD0Iqmlc/Kkp2ZvE/+C6d5AD30EuP
WbBCZYXHXSmUhdHr+NCcLBPqNInlPpG7InG+Vn6eP1GTE8NSS2szlBeovcTiBbNA7k8FLu9fPZSk
gZJWkO5VqT/yX/93tHXTnH3qhJpOL6pVDmQ+mBrDSGwNJOfTg9rZjKafw+pvh1ELYZKPYjrRWgU7
MNnXVmz8kOWwhebnYoKWLd8owjy5BPkCA6sj0ELR6C46++r3fOqXgFKOjbF28jLzYfIQj14vrTlx
x3HGx5pPmbjMCSZRYx9ITc9vEA1FCKu7NwhOnbjsmuJHviVGCaYKgonP6eNzuypDJDCsb/5cLp1S
d4fZPrUysyIbCHNtnm6yAt+AZZnsWw/nt4kEAomnGimsZKuOtqDNUEkIgPSZSmNgodB+bLMl3Bc6
dQSh3aekP97a+Ug55KvkJiu4jV+I+oxJfPrw5QeshLaiXCLUgdU58EyN0/W+hifjzcXcbSF8GH53
Ao/jNHkFLqLNJHNtu8ozilp7eA+RFwf4zGJSngjfJuMvM1m//olO0JAVE34r8NoElje44T/4Uj7v
i4jPi/wqrnEb03z4ku9XYQ4apquia4i8H9lUI+fXhh8PgjlR5RYdqkqSe0hgiHiNRYAdonHTofE3
okQIHr49RqoOFAQughK03GQjhda/NtWNNBp69/9eCCX6/QiteMBs5aOxd5Y+Kk5aBpIBmlObaUhL
6/Z7qcspRas1SCoqUWae+zSPQRfewOvxnt+SLOivf8X0++8hvHevAhzVcrl9RsiVbvwN34ZhtIp8
p6FBb6Qr6bOevJJjuTSoHQVI2Z85TaiSRxDTmSQe+UjZ6AYQm0KAKofgjZT68ea23xUyqfckV9yA
8ZFAF7rNBkcDJ9N7tC2TX4BCMs1Cxa7kgS9qxkjuvZfdPFabUV1ygpiAROcwJ+Rx72MZX0gqSczF
KeUCbrKqNS4pHbvWvUIZYZaSLM460oQXzRf2H8FFvrfCiUbgYvcnWCXofTKU0zOlPLHu0ioXZ81A
wiXhr5RTiTlZvFD5Z1Ssbu49BQTUPSgn4D98mz8Ka/+mCd3JkFEmTsuo/Engca26OBjj9MmCXqeL
Ak+Z0EgPX1D26TgqHF+VeuAAri11lrpBQqHq/a9pUilsrO3JNXxp7btTlxq7O7FurcSX0jDTlU3x
Nu9AYEgs9fo1p8TtPkqlsEI5pl5blXFBPCW0OglPvnnh0vTLMaI4qT24zYYIoQJlWiRsy6B0MSsy
jt2d7I+biZlFqJfjGDwhWOSWDjym7iOP9tjNmrjTVgpApkqJsrAGmln50CiDMGsrDbzphe31GxHL
fNM2ycKMQNkBWY4Y3nx/tDofqqcWSGGOU/ViWmobxc9IO3wteXTeCNvMP3vf4ZksCDANc0psdhS8
a7gglRCUGrdbA5p4Ma9y9mlrgpwvx4uFz4RIYra9Y5EM/7axaIl8gvWwl8RQvzWIOrz1s8bk18Vg
m/AlLhTBtq2mI9rQeb2ieIa49pwrx1pNVKm03L5gMComMQX40yA27b8REh+FmAtd0G1NAQI87uaY
V3Ww+DoL0SZi1NS0K/4Kiba+ERM1p3vKvkZwfPjsc2lYaObmg4tNY087+CRmVvmchGZynE7Z1Fx2
9wL9NbQ9Z5yWUvLT6odv4Avf8+XCgKhHaqQGH/UFrylRkANI6D7WwMIkYBTANxzghFfukUhp6ZNX
PlQUtc0bCYcA48ZGZ0Km4Af4svaU2ameyQG93I63ptLagr3cHyHkr9zqy6EXqVmAjaS10YVnA0qx
AUZPrE+iGVO9Bn0gfDL21nQq6UdDqpjrl9JpnrOp0zPXMxngPng5JGZPZ0IOiAT3JcBpbU/ZEdkU
XFTjE56YM4ddCkbLUz6xoArw+n5VWPBMaCpzoQrBgVYCwuJPScLN+9pYPxCCBwsLgqWGRN4/D0CY
gO5gcJkOiNrsCmqFO+FtT/UT0IyA6yCbSPv4dVB38ZeVLs3funKbDLeLZptTEajFmptgX1HAs80c
rrcfzyonUU2X21S9Bao+VY/hPO5sAnpklCJWdF0KyatVQxnYW97Lx821jv8IQ5h5WAP11QeOCwiE
qA6M2K8GI3Nz9GDUOeJufk+xF4c4UUO1+mDatK8ZiZuy2SUL3c6aOPSUiS4p5umqwhIw1DDypAyw
GbhGI414iWfvNt5LlD719Fp9mOGMVsV2Z8k3YyqCXLaO7rp+W69HNyQMlWgE2RbJp7b2RfO3hA8u
Z2vXTRwAXKtrnHGfsHc1Zbk/5LlnMcN8vWxVePnN9RkVkNaN2KrEFT8t28dguKagl2IjmqTqXHr2
3uk9xps+ep54p9AR/Nm72q9V0Io07JyI9m2kTFNX8kaE2mqYSOIVoxWY6Fb4rDk6v3+7Jupb8FdL
UYXoKZyyOhksaMANF31U6mtcb01JMuqHyst93h0fO1Sh5khbSk0UEdU8Qr8Kn5m3C4h2/dWfRYFU
1LH+yrVixqSX4ZKbN21eu4zJTsHvHhuTwnmZ9eRL3p/heEPq/DCwr91zSvwqDCVLURfYrjIXqk9b
U9eSw65/g75z84hhLbkEa/hOTWMxxxLa5pNGTFD9JhCjaQDRfq/PEa1tzXsyUmFm/HE+SV3nOvIJ
ulSmEzjU6fq00XHZs8+t8hlOj4g2hL/f6jMOm0KZ3RTkItqmkZMcaJ1/gnLi+kZw99nRTSxKc4pN
8xpTAfsfVWqOJI+D5kiTZQ8NbNhtj0BNGEM0gtyx7Slyob0zBOHwl7v6cnMLd8DVWRvTiHighAZz
NreDnke1llgHuRSPJmXJfmpklH8FXFKrgJqBUohDAJQXMxfYAdiPiQ3uGLZPbHCvMs0IishVRX8x
AevKKQVmc3FG3/QamjDmp97WlzgGULSZSAwOX+fr1TejIUL114l40EFMvaxATYC73++InmsCOQpW
UTyUwtnuLwHodJu5+YvWwIA2XD9DQsfK9DDOOK4+FXFLRpFMmWMc/LKYLpiwGIfIsT49prhmb6zI
ld0MFFutL2PiMMmnFIN3uSN7kVW3e0302ybl0qh09yBIAm9MCgRM0x8o+ovss3Ra0Vmg5Ffmvcjs
F/vmPkRdfBKbl8AoiWmX44FUeH01edERGzCb8bRjghTVXfGXapgPiq2Opon0Si75YR/yOkDtFYi6
rguP3sUOPx7spatrIcYyLJPC2xd/YEft9GWC7YcuMQowenm+HVh9qlOUaClrHtnVftowR+anh4ru
vDMbNbacF2dW4D/IPdfsjKanunH7zCMjhbJUGWQtrtMSVobICh4huw91Xj7/tSj2OqLPCADzTVKj
HCEM3H4UVQEy/VGTIgroHIlh7ekkWPE+fkAYX3lNZXOg4TYQ0GNvl8PvQZhuWm6TmdK9pcbU+I+/
iBQsbWGH2rEE9MT0Al4CEZgewe4NLq7d76yFJRUoNuGuiYUFTNf9Wubz97LFmeVbDVJBjqoLzIhF
lAbUOwSYTdRjQxf9hAr9zEHLWYuzV1fL6ZD83A9/j0YsjSL7GkRdy35BkU4L9qLwBlaQPvsQ4oNg
wR78QkfehezmlnEvdK8pdUDVadSaEi2pm+JHOq0EOfPF6NL90UnmlKIiTeLENUEZX57GyTZ7PYVT
JTZ3dW2EfIqkoSc7i/0/yneEeEFz4k8GOz5F7d5St90MLuPyacn7HrItMkruMpiI+ukRzmyYt0e3
8fB0xOaMhiVw52ARQHAXv+lOkOGKr0P0tYaP3oMFaVNgGRRy8svb4LIdQ+yeA6ATDHcF3JvD1lOE
k3dX49GJWEx9suZd6YVdJIe3ZQd9aoDjjOErih58Ndblo5AQb0cXhfYqO0gWOewW1ZlNYOVZ8m4I
TKZxV8O3TTJdXhuIJRIGJPkoYVnAy+ITYVROzEXBetq7ByrAzvAPh5Y2T0K+Qfg6BzkrTxC+x15n
k/4Y4cBG1HW/Ih3xrT6IcWYn4HJABUtZGQkhDBsUubpGi2IAqPzU+5wYXAgik4I9/JdrIbW3S6Iq
PkgOjHgBXH70dXt28guXMB+2/MOpy2ixOE99dDf3GxwH2kN53sLgZjt8n3q72dKx8LpgTMjCsmdS
PsfXHgoJjCTdM39AqZam3gEddaJPhe+ntLmAUasKnLdUyHn7ukKIfA8ULPqhb/fOXV0HK12stnOJ
CbXez/n90Ejx1Ho1KknxBlZ5XBpDCXLHKeIjhJAHcMcxskMiMz9O09aYjMh4Ol8vogUS8byjnti/
vCOM3UY+dhbt/UukfSaDZEQPmSvtxnNL4VnIbuC5OzAd6sTecQHbe4tZ3TvNhTZVvIyCMQu7MqOm
6EouPuEgzPot/ZT7OgTsRdGMlq+DXJFdHAJ6T9aL87kfbIqKcvqbt0bxFKU1m8URYljGR165tWrZ
s/5IB9PxGA9OIxksopWnY4u7PU20hy2AEOWTvJ1Sx0E9wiIdj/hqSmTvvr/G1K66Mk25RhR3Katv
2qTc7akmlWw89e93yubsSZR3ge/ZJse7fj7Sgv+69gmV+DvRD9P+EsJj55PtDKFm/7fDfLzPbsYD
2ycFksCuhocbJdz2ldibBYYsGT3ID1UJE7iRX3thLt/bzEk+V21uRPhq6sf3OBDtgRwb1CGMQyUj
c/SRCtRQFOUDj65NprJomvC0wlx/Ze0iey9JkYk4N4r0DLALhQUgJ6qY++9JXjebS7r4qCm/4NZ1
PQvmbA5HywOGQ6mJ2EHMBOMscoGyIFtoSHX5l6BGDT2tXQboIQ7gj1Bp+lP/ElulaYjBZ963O/OQ
9xMkfyyk7CEciJ9AK5KJZFC93LID3EqiZCWzPdFfP/Z0VlR0zsWdL8Uo2uJO/ICVzJkzZylIm/28
X7MPyKCSwbRQL0Uh7BfUtOYSs+neU+SIAaa+5kSxt9MEaAVh27l+h8Ls9DIJa2NN8+S2OMJzm282
LXmKmTWXMtgwtyGsqdP3GOO5mVTpbToa+V6ODkl3YFzb+zCJj5ij9jgItmdTMtzuUOV/sdw76J2d
Q9xZ5Q6xdZd7GId/HVo8HHyZVeGvDYIXD/GE+VSIaIEkGL31E97Ru0JOyV//BMNHG4gGD5lIxc7O
GAteb9dYAc6DB7qgobYZ+kpkCL8YErsEzR512XlvV+XMPjlHZoAxgxiNG8B5C7eA2wCRE0dIjQl8
zI8KOy22y5oMjdsiB8MHpibUngRfN+HYO1PdfwK0/LsTaQdTpao9gGnhJyFoZveAWPG9wrMXQ/oR
rr2nXkL4tHIPeasm+Ec2l6+h3fVvWVenkT68FYytVnYgTMMaLXS30HbVJuB9ol98mGtHWfOMW793
nM4rIqADHXMPZ4K6V72oKaRl/n5TblqZFVDTVZ1p1ilW4LPOs0BxMfPg4AH36pUq+2QaxWYi9jZV
9MPR5UStdNWEn/N8LR6/sGog2dnIF9ikGuUZr5Fuk6+EeEs7idheLZJbOj6t6psa+6ZkKowd+5eS
LGxh5jWoS3mvxM9BlmsUmpEQvgiLOGzoORCdFzzeeo5L7zvdq6i5Ku9m0PMOUKRoEBFJOI0Z7QUz
tbZUOl5aXsOeCWZlYLpPB4Y1OYsusEpNaRIdVaGrdRQ30kivvSVQfJZYzpA1vaS3yLNBr5LpGLQx
12MpZo33fmHQcKdhDhbty8eyBdlFTCtGsJkbG//VOeCHYo3O4OWFY554KEKpZRC9c8/+mWmRekJd
9XiuhbKOTcuWLAmBHp99JHvwGfmTKOcGsOgk6rgAb9ae2upjFrcmaBOydBHbUegc7uD0sB2iP0lf
vNBvJpFaNlEbCuohsFh0XhSviuK0H+/8uxIprGGEEu+SX7iNPLqUqasWEWjSzQf/4waAdpK6XAfH
V5llbCXkc592G7v8eEiPipTTDYoNArAxdz87gWSiHwKLE4mmhnf3CCe8t4cmrGfgAGDtgac73m6x
jGMmUrhe0qXg/w0h+G0iJqJOER1xAC90WHqTaQfiUnYudhAfstpKvsILDvQ2EiApnT0iviK8YsvD
L8XTyMaTrr+kVW0i4SZXYTSk0bYyvSYCxkatHB7Kkqr9TWo1AU9r4rejItCsSU01ewnIt7TCedMZ
3bVLnpfpxLoic3DooRmJWRwbsy5TtqPuVWwz4oBg3qVbX5SOuinZ1pJ5Is5Cs5E7OCili/CBRJeS
oRt16ZmHzi7lNjDZwV19d+UELD5uGa+Lx15N5jcVJjVNAEODxdxQPiOPs8YG7I70hrn2UIqNYiHw
xonDFkwZLTbwmYIwtctXSE24rJ62oEfdqSJ6xv49Clo+k409BvCIr2JFOqlk8tjk6fy4WHqWoAgs
CKorQySpfw9LlfTQwxncXYoFPryqh9mrqh9XfGrnbe2GvgeRuK6GehKFUDS8fcRRED/Le5tMd5YK
C7eshM0YGKz0N6KDW/zmyPDSKvBmR0p8ukYE9ao3Fbbih7J1szdsGJOg7mBLzGs1VNAxQUT7bo1X
agL4zw9pRX6+WXKVw1+0GW6M+DHev6XvvQ9Yj5bimT2f/6reCuju9H/ShVPXH0WzsLe8iZk91c1j
YuezvIon0OVpsbKv5fYjyRlCMmqRqFpU0Zc8iS/01OYPjAbEZf69ysmhpenuT0MUiLoVYJ/EdSJ9
E2wKU5qkOwC7XAnjiBU4sSfsomajPTMWu6Nw6oJyKPw6pN7qoUAfW83M4EdRfwvwYVO4DdRbQlpb
71gpNN4BkHKBccQpHUAwp+YYJ7ssOqfhflCBa0TL2rx2G6iACS+aUIEuKX7JOWqtDhz4R3YpNCoH
EN+6v7ewCARZb6bkGGCjIvY/OU8PB56mbWeZQUsvWEVF7M2iLFH94MZrvCQtUr/WijnuIPEJx/Jm
KEqa+PlzA8r+gG1xfObro5wEHiJaGzvTWtix7/P3Km2xiSdbe/o1F7OA9OC5VMBoWOtxFt7tX7xD
ORZAMHFylfOoA48MghPe+Y1zFKHc2ISEYvkaoMzKT8/suc5VW1LR4FEQlkiWR8TOXNfszmJaHYd8
j5dFZ2GtHRMkZgmdmsV9qt9WBJrg/H+tNM7YBOqLTGq/GUFT3P/aHzRyw4Gkk+9tX8aQY3iG+38u
Xzr+h5HAnTbZ8RTUzPTjk7EGJm0dN5KQNvTRp8WXhcQJRlhN1ARk+C4Iqa2guFifZRpOKiAZuiEf
YL6nTCNJKlaFKhueu895NuxK5MwoxjbjJ2TnCz96QBYFPpWFkNyHuQVydR+F6CL+KNltjQE1EZTA
IXoRzSLqFN73VsvCyCLmNGRq9if++anFDVqZWTMQH1DtZTzWH/IE5AI84XUZ6GV+O2b/87MPOn7s
yt1NyM4g8En46jG7USotevatFUyW/Y7xwtjMDVP+a7h1qf5YNQt2zIzk8Ctb7YMo04DbelTxzF/i
kVCH2VaeiuxnPPn1LTyO7QI5aPnC7T13mTVed4RoVFwascIryMxkm1XvvRUI6QwgoUk5M9QIE+4m
vb/5OxVJFUzcNar2sTfHhLo8aGFjz424utyGp7rPunCmrcHw/tnBdbBPNQgp7q8Nl692wP8xm3Ie
HxYXyJ8iFa+uJG3sp3KH9nh8o5wgTMFH6jggerGK+bKcolccO5wq5yzPmR17b7xyvW4Ib3iLqDkh
ElCTUZHkwPM8ClQ+1f4kG84PsXoTBPwBAMXY+pMRWFFO2IP6fMPih64V/I9dz8ltV4f0/jJJw+Xb
avD/aSHS3rFtTWBJuLz3r+keYNjNDAF0Hb1u2/HenkWvgbkweh9OORVs2LskBikDZpxH/eeOcNDW
51NDeKmpq7LOvF8NUmI7SXw2PAf+TrdHJeXpshPh612Wmo/kF5VifeNDsgkPKWIQ3yFcU1/KUPMo
8eMw4IHA/96N33162sCST5QRQR8vgajzfJce3OZmHRBgR2Fs7ANKZ+kyOIBRanoJ6AeNSB7InwVk
ThM/myE05lvK3fBVckbx4b/Tdpw6/uT/7qHI+RT1dLYVHe78Pe1vZ3/EmdmbaBxVqT+bg3VRNmxd
hkv0D89Lb/aD7OYZB+dUC377aDRbJOzxpZML6yCJR/6ZXn8Pco1IfsU35WVIaeU4FfDo737jwVle
XRaYAWpY+s/u4X3NOR0hM5MdN1/GbuhlqGRGNy4ngDQVxSL69BF9qti2o0ORL6PPJlmcW8S/wM+l
EASRDvubR6M7Fv2JoavQuSmjYfkEnX7d590Z8/7LRnYujEhxRWfdG4V5s1L96m06qFevojz0ZSHu
T04RHZhrzFwceqsLASjG5vxZ3Ns+BnVC0UjotcDaH8irgRx/Jt246XtBMfyVFDkaENnnrrwDqDM9
zax8qs7shX/A7rlvd7Quqp4WWfkA826Vss45nMnMwMU9tZh0zxBKd+MaMsYGCzwbTyFhx1vnPsV/
FvWLgF/JKYiD+Qb+2JmHkAabSgG8LRUGLnLRCauX5UoKn9whQmag3xUj79zJ53+o8Y2YOz5S91ZN
6r2/HSxpxFRk4p9lnls8N0VfrpF1t3aTieN7p/fynpE5agdRTMhFx3SNVZStNAJUGIz4Hp8eitiE
PBTPinm0L45IziW09tO7uOmVzmt+ZZ1YNlGwWTdbV0A+MhMOkTu3ZYzafpyR9TTk+EcK1t5ZdioR
2F9ZrguVeMGzRGWszAx0jTZW9lNbs4ZJmrXzyP9ed3OBwH36MXdht5vsSVe1b2quXuWytZlXRjv/
d0zrbKNak31HKQBf4Uh27E1bYW8u2CWsQfYa0rVsAID8u1IqwZR3snKR3lK0VP8QtrkxnXWBjyW7
3uyrOgRp90AYSLvr8Vpu9e69A057pRVcXzPp9nSdDixyE5Xsg7o6MxzEXUyZyIzFVzXafDtbcxZJ
j6Zq9eWC7QOtUioIAGHmxhygzRBPu4Ed1Uh4hfR3NXTXrr9G55LDOxUHjk6j7NJ+GBi8uxYe9CLE
Ots6mbomQInr4mKV9fZO9Wens25GfSakCulQ/f4GXrzq8AhdKypBYUA9RVHmLsUz7uVqxfoVAN1u
a3icj5i6Txb1arIow0mpVw6W+PxZdq2udI4Xyobcj3Z5QU4C7ZqcSjqWALITQTRsl+HSxs6a5z+P
hJeW/ZVDuvQV0BVD1AnJK/PlR6MyW1cfa9ISNJStvzephdZr8n1dlSUEjSjYDXKItC5gkmxtV7Yp
8oP2vyY8iufPUn1wDbiuJbjG7sckYeDVf3MJZ+h0Jd/GU+CGRquZ3ZPANtpQOZeQhHE9E7m3wd5B
yms3r9DgT9ZutNSeVYWYvL8pETfgpGityiEnx8jIO694bWrSVRXeYn1DmluZmmUdJyxbByUtjSBP
9vJRwUV09eSEE4XvFsstwS6RL+tIYapmBKO16h4sq3zStAuO4197h+WAmaj5JByylUro0IXrLxVK
Gj0DWMu2Rn7SeRgMwYt4xb0MpT1Iv+U5jan5SGYI8HMk7zKWR9zSnfsViH7nmqum+wF37c5qTUAc
m1Qy0tne3Wi3f6AOSd2VvEiK/GkpDCMIwXtooN+aHv03vsIWsLa8WLRN+jBaxRvW/LY8rIb0uIfO
8vGyue2CBUgIUgnguojjgozHlF12kPLpW5AGfXPrVqQQRjTW/w/P3epqU0WCwUcpLZnOjmWCCKjd
6oKtgBE2x7lLfAMW6czG9IfUZgt1TvGKu5wJOmAwJ5LpGBO/Rk9oqpcFTbXYYeoN2YzAli82USee
/RUbM8kn3bXnPguQ8lOuD/wEX0O1EzZAdQkMtOmSjBCV1FGBLfpa1z/vidiCcqJU8Ff+y/pBiSWG
7Ei4FXqLenXrH+mru5Foir1QfmMNDgjPFuoSQ4V+FWv+1A5POdlmYi3a4QooBqWEyXdkx6QsL++A
YVfXt+coDwQAoYx06/8K9tSdkEI+tSkWxun/EOs3XNJu9YqRBCNTdeSU2FU0EaAx9sXhcu7F9YsJ
KdB9tVrLwOW8ooclFK6A5QS3+SLxSTaSftt7N45V3Adjr7qIbcxoM8t73oxY7i5841yQ10dO/7HC
49CqKjQkhhOPIkuSEnTwhOzmbm5Q/fkAD9ryztAImbcUtliaXgixlHm1HMFvVeqzBmGYm2jjDrcZ
1VbTV6hP1g4GzPgYOWyieJBDNnAiAqzH4KCAnspg/ZLSsFGGu4mofil0d4IVXlNRlK2WEPl/muRK
SLNQ9AY9UDfNkaJWd9wmb93etQHKOvG7fe9llKnY0EseIguqNNMILRhFfEZcKqn96T1z63JFTRhs
IF8V5AObWo7pSQQtilF7TJT5JRLkH8yiskO5F6g7jto1PgnhBy707eyIba0DE0ECzU9unf9tsosv
KiyCo9SMBbHTUbOLRraTDkOStzOJVv2pC3fL7qt2o5TH0d5kp4pLaK7xPChM5kUhu4L6uNgg6bfG
bY5ccJ5joaxkiQGN4nPN/cpmKEDcDXGmEPvNZTvOGn33CDcBdL7rP0ozwpY2jn3DA3bOTV61UhY4
OVUSJ0a9GBJQbUZVEiEu8+Qfm5XqHYqOCLY/EZBNC2yeVUjsfJI4A2tKxhlLjn8sfXW5AQeyVCHM
fmm2z2njwmiza4wbAvAbkLSBjHeBL5Exmfy4o9AZbds1D7zYBxoXxxT8byuh6aY0E7ua3UfYSwLs
kQ5YalDs4HOqjiDT9JiGOj2vf3x9RpQmDjeU3JvLccWqycgNbsTqyOLJZAoO4yrUe1KRwlb4jEQW
pdTz9XfA5c3RWlU5sK0HwEqqNVsdAlMQYKod7cyOuD+NosSrDC+bPPx4qNvy/9acOtayLQof/zMd
9s85Zlu3/HllET9RqmZUx3zSIleMIAfKdOU6RkvreM4/lm8ObMSJPYCL0tCZNWIxTTJV+P+H3GUP
Q5tiow4OfMU+3ImjZaOgsoBJLwarmnlmM+0KsWp7lQRrNHmQO3A0sNvUUwTXWcVo5q6TMRTE24MB
3RrN503hGUGgmtT+xnVBLNjJmi1vJS7lJDo1YJoNvr2xfq0KN8pCJ+Y4hbAeUwLAfAtYdqOIl569
jXerLuE+/K9RB+RfPwHMiWROB0Scx2FyhKW3V7LpxtgCt4s1bNtWyOJBWOjZZoFpgpbLtALE8rBX
2HwZCPPXXvURBRtbtSLEgaCD4fPcSDVMp+NzLhM3YUj0wR0tJygR8jn/uza1oPc7CYr84iFU8X7d
/RuA7M0WJDEz6hz0pkEWwDCCmnZXfvs4Gqz6IVAO6jRhON3sc4AZ9PBdhH6YFP9Bt0Xj37sXNkJo
x1BkodfCW363i/N0VDxdQheUtzfcuT5rpXhUfPtWXO5kQQIIgY3Ju/M3mn46zZtMXwWHtKEh4hzL
jNaloRU46ojKfGT29gVCsHvkjkAtMKpAk0jr8s1dPGDAWbprGjonLG1zsx/iX6fu95HcY0OKMPnF
+V4HwNWr5yWkHYTkjPEKR6CNg+FpPjKFkF+kGFe4GfhfOKzOluKW7QSpVc+mA5wcw787Tncz9g3L
cyaIWG/r2sK5tW7R52Iu4pQsVZ8BBwoCZi7vhd/r3Wbhw/cMwvL+G15AD+HPozUpfwukDqz5xulj
qdDF1IRTFBLF/fUKZ8ObUJ1V4DWnj+KHGBRfZmnHAY4slCypN9lJpT0iHTQmSuG75025ziwspwDp
ZU6YXs9/lptYGrvUY+BC3+kqjri4g6DA5A9n/hbHq7BRWIEzvJw+Qi1d8Wx0cIE+sZ6mF1AHiP8u
5DJ1Oy/M475NEk/FsZOyD6xmmdiz+mg+IiS+fpqSRF2HsQG+avqwKZsRtQuyX7rd8JMPeBMBxY/8
ukynldC7eaeM0JRj57NcBHPedqn+YY2gE3tq4P7tnEZmjfPIWNwkTUMdk8a8659RDP7PiYnX5PJM
rs3hzNjHf15mVpHg8aBk4ymV7OM6B3KLi1NWIpk7qka1o//5doVqQmGHyiSyz3q4d2MhqvpAZcZp
WU8xfHMPTPAJuujfdIl1sheJu+ytFqgVYyVO6tOAAPaxzvmyMeaFWXXBL9q8gsICRH39eu/a9Byd
7X2gV15x0zG6/espGIpYlGeWiGtF0OvRCTIu9MloxCYdxlag+nSE3CkOnX7U3H9RuhfukCBS+XS5
bVG5ULTM/uh9eyHuDWB59op2DtD+h+VljpzEnIoW14FGkLjOznoWBcvT3S87xNaAwA1IUdknWvlP
Jz9J0bqcZ2Mt1VR6h66NaONU/rCarb1kPVI8vyHIJCDGnuXT6mwbG7qidaO6A6T5h23NcKUEt1u8
d8NFgW/xZmZZl/9+ku/QgOUOy2WesLojL48wlSRXx9SKY1KEOAdcnBT2mfOBCtz1gQBHSBidCWkA
GimpAbV37WeWRsXQQVYjiiaBJ8QFw6c0oT7KdQoWwqGzj4qhpTOmxn+HrS0H9MRpcgYnvjnRXi+a
LOweHcdPVPLTsVLeGNeiR/MwSBjQWl+N7I5feuH88ynO5hUeatrjI0NkMwSUIInMUANYdxgDXEO6
rN1juHHuKOcdysWT2jP/Bk9Dq/jRWPtRpN0XK+OyXHYld5KUzIOXIH9sLBlssYjOyzdyOLdpwmRN
AMTqu/a7bYjy9TqI9CYdhJMYrIYQTxajx2y0NZ+6qI6h8RB8qDpmQXIEjoDAHHDIUtH/d7du7zEz
vCkW32h3SgmqHYFn9T9DJ0IameDbv3MPeQlvxEDqLzwvkaA0vWe9kUTRZAvQuIBYgMMcmrYY4VGY
lNQnEUvyFUbrUkrmFNyd8okau48MrwoYXdLBwCd7D+RFz9AgqhdiTW541WDln7ff7aatE+rV5a6Q
xiNqvtMOU9IxyNQCKoYRs9es8j7Ppnxs2bIn9wOY1AglGVXXAssK18vlnnvkiwa1JkpFgeSw9+I5
gkHrslvq+SU1uMCKgGgfKsMiton5SuveUP44jdDmhbfohkqN66VudrzHPgeVMdea4aMkBpHgsp9q
zdU+NdU/3x7FMuhNAmiFycBcxhH7LVVvKR3hSIeJKruE7x5QHi0l34XbOvQ2BMKeq9ZclPkVM/mk
nG0yY2Gorfg5z2EdqLP4WPryWIOXOi4vzeUt/PmytTEEj1FmxhkUC3xhXbH++UxJ/kWEyFl6DpBZ
6Yg/j1XQDpFmKy+an0OFm8ZjfTnmX4wlX1W1KFaI7KClVdwzRRxvq+O7mW2JFCxSFx9kbDMj1xIb
3BMtcI5yhswJa/aLP3KE+sxjtBKQSk5lyiYuGH0+J2G+KCI8nx58dqEAvkQ4Cw+mj7cz7R/QPK9a
LL3u5AQ8G5f5wL2NXqwoK51agz91yck8pukO4MHLYPLwkuTj+dQ+ulDOZbFBCxKE5dOxX2haNp+J
n6HIhzj2khT14IepzGDlTkRMtA5VAhbIcQBXijaPpSgca7HrEqSLVU1/r4jV9k7A+t+TcF6LY5f8
AMaQW8FewTuxcmVUUZrsxYK5vg9VuglqRx0Tn+b/kJbeVtN0lmGCDwKwVh9CftXIkCeNt9cjwopi
EY7S7wzfwa8StCSqjkxv89+IhW1vrxVIlj7Q8/SO80QEaCAM+xUhz4FsbXGOgWrabt1FPzUn4Pp1
fLzpOyWOKApKGh/+VVrzFW3DZO2rr1gNfrd4Hq7kEMrCU7r3SpgKPHGGwcGLInfXJOkA8oHjuW1d
SjKNFh1jtnZnbcBmCZTZ+A/LFKJAyvuWyOm0OiFgkBwDyzsWUwi+R3DiWiL+DvPpuibsxao3y16t
f3I9l1vd17R8gAupdgSFWjUV7ahw7ewpgkPYLXcuRF3O7X7CKpgx40R3y+FrPJeYROsOpimly+zK
CMeEsw1ocTD3HYMVyug+uCogg9ntPUEH5HahA4LGeOOO7xWAVVHL253831uhbvaBaRvoA18lI1mz
oW7UCZkZOvb7NjZdl/rh4aAM8Z5728e2K2w0ROJnOaI+0WHQUEWP4xyVTh/LbV9aVm6Qm/q52Oal
rOWP3yZEjpRHp+6t4VBp0iXVzH+X3EZJ5InscRmlPj8TOcnuvgFk9O/0gudpd5K6Dynv5mKVLbkx
RrPeV3lorW0yW2xAIOcZvohXgUmCrevfmVRFq8MkdmO/FHD/j9QPzN6QA3AsvPGkkNU+f10ZES/T
KXMVEggDLN0WVYX5VoxlkQD8TJb7patV2ILNnGfkAQJUFzY22juTUSFkHwV15X73JdUfQKUb4FMK
2UFm51WFOLZihecIFezD2isF71/cQNDwIiPFj2DTeGVraebGQeKGDiAgJUzmhnS88U12pqfDjmhP
xR1RYCxxg0QKWjPuN3aDBZtJhO7uMOtlqm7XJP7n8x3X5W9mJ0a/CAYYWYJG8zaN4CD9SUtMcgX2
if50g8ZiwAktuT/IgnbpiRzo9tJfXScyFaic+TazjYG7OQ6zm4ittaX2bt/ko/q25Rt9L95AO0jg
yzis2ne6byZLObkvMqKfX97wQDqfOAJTw4XYXjLoHfvjKnXKN/WS72J+1oz8IaWW95qZWLXVNKfs
b/ENoN36htOvlyFRXEYt/ySGOLAcf+ofp5zlhLLntTXsA8NtHfebu1a0y5soUHxIfO1sho3DyjK9
CI/IiwUHhN9Z8DJlDMj9SDZ40loM0/88wydCV9Nch1MO7T0vIzLckwDBz0KurcmuWFv2Nr6TE4qr
rb9d1SJd0ZTKuZQ3ePFjtODiWuUbLr00DXtXyLcmjLW7MUqqs31QdOEy2XFYeTgr/Vt96dOPl691
F5MMHO8uXpJM7zUbnx1z54ClROvwa3AOvzYK48i4ciq9kwdyl0VD95ZoTFOMDI7eNMdg3xQVHIk9
0NUtWtuPG4V/YFqk9tsNL/5lG9cnncP8p1TbDTJ0Y5MHfpwana/5fJMqrLdiemtYX4IQnlAXR72m
KezFkSAsH/WHxzoAlWqXB7whEvH0Qd4fmXkILIienuWhhdZFDTTmN4b2hDeX9647Z/NmikZYCxRk
GlXiT2aorDjXWHRqyC7lWDuL4wr3/U1JQerJ+pQR98FQpKMWWIs01Ht1yMgQuI8jHObflO49HE4u
kWUfh7wGLGQpcC8uRfKqkvJpEbsUVritgTg/zjSJkw4n5omO+fh4aPXYKmzY2VCdDUjqy1puFBIG
lH+NNarRm4JzQF7yMnML2c1/a5uI/29xoO612aeHT+2WaGWq2ySNo8y8fDHe3vldBRdsKI9PL6Hn
gOpUPzUaQ6N6Gu7ArAm/1P/+P5dUyn7yjf8x31hvsweKrGiRck5F0g5KaKGVu73OkVC0L0ytvUou
dEJKDICgUg5l6KB40Jok+3gf/nviDxjh7wR5Yeej0nrEIk/pysf+9P66WjApEKvb8eMkhG5ctEd8
MvGXYtgLTbWAA/5rwVpqRCsBOFhHwgGYTpaNeSefop5cFeQPLQLUeXIewONErKgYmLVq+moOEhr7
CIMfizH6REh9AkWYLHHJB7r39Foy3GNQcVg5c+43HCr57yJ/4Ml7RzLmTx4SxEBfx8J48ECSLWIZ
JAS1UlmRG4R6G96b53xI/H+Oq1moXhUfWZOFHriC+jixuuOCaoM/wcUzmUjnGXGPeMEQ87rwvj3A
JtanIYRKJWhooPeLZnJ6fXrMGJseytfPaACvQafldoZoHUQ/Fl0gPWO4nb8EokqTObz0cXh+I58L
HpnNjnC8ZQjM8iqAzThzF+mlkz0quzQEcF1GufLtR8QFW0ZUL0BlQVTpOn8sXz9UL6/yBvzuaxNN
cyEJgPagw8V7yMmufhqLjKnUq6eHQPfJ0m7GNVuuV9mAQrqjXzur36hyyV3gI3B2xBi7a1s1XYOX
G7MA9J/68OTDjjGUGx+4ba4Soa6GplXoBr9LnufsN2u+nW8MteHOx4RXuOgdxPJ2g8AxqbrhfEeJ
fU4q9kZ+DHUDVCM0ZSN8iSXHi/EDto85yPQx5Ye9sMnTlZMLUsqGKgF7fs93lwB8llODZibuqiPU
hBp+lc2mxL9/H/dfBLWPGEwHhEJyRomQd5fofJkzTOEE+zPTOeNClBP9zwSf0xsn7gj8j5YRxdDP
kRSWAu0uNhiAyLtVNRuew01FX+T2p+A0bOPZM6Ob0EPyoqcjw2YlDXkQFuDQiUOoe1gl6P+QHzM6
llbOSTerZlpGqnBzYE8MUO9NZVm8ooaVnyg9EtTjQ/gsHVVkcck6C7vjuY0z/XdvOj4eiNGaTUcG
qCwwEQymzbcZ2Ejc48H3Phc2pi6CxxGWgvFhTjq0G6Na25K1owfdMqIKIF1jaD4TOf9dNIkf95Ny
hBuwvDklJn2PvQ+q49Oc3ADvaJcufeO8St2SaPvZgz7rhaSxodZ+YiAJjOfFNLLEmViIKLBiZNLT
XXY29D1gIzCGRxVe3pgCSiTRgYMZQuo8U7BmezLUe2lHSrUebEB3WI787jjiJLQAOmlHna01KaN7
xP7cQhboiRFH0BK9S9gSKUTNlz2XsrXPvCqwd/5r5WheMGr8gCWxFeGqPFqJDEhsuWtvgOb3RUQP
TLUb3TAQYfgH7/QMnfCnO6ZapDV3f/OIJHmLj4w+asnSV2Ulc2Hlr3vT3UjF0F/KZ8bWI0E3d7RK
EtNZaab3U7Rqf/Z8TFneseKN1X4kLfMlLy/ebE+A96hGqj76SmKF3LF+kVW10l/TARQ5OdoBrQmY
HrVp2Bd9DSvmdUAKg36owmCoexSryBmF7Jhj+rJr7huzSbZAawEhU7bmFyvGw14G3HcJCNrp0WRT
kIidEbqupxVAOB27Fcp5WNc1e87TDxDJtF678h3J9UEgBVmPpStclkFHBgee69Iiy8G8KNg1BbBL
FCxFrjFXXu3h0LaGJvHFSv66WXvmZP+ko6pP/5ySFJA1WbCcqEdDbUEUfsxX4S+l47yaKOBiIjLo
40D7ziDHssi564190UR5hmHQBCW/LPWtDThSg5gkuOwn/FpHS7cDdVxmRDbEQ/YKhFpHJXdkf4wR
IXJLGNYf08j/JnpdGbKDbIM1/OeAt2FZtVI62OtckTFgkyl8Qv6cwScEH229ppl5ylPbneKmHxks
kp0T2Ux4SRjhLZ8XwgX6T/JNDop1cBaS3QGgklWWAj0k3QKnhMIFeJ9H15yvr3AbnKiy0oYRpqpS
qoqUiVvHjg2N++ec74bGRnqoOQvurGIiIRz5TjB0zGTta6NraY6mkY/yeOeDjbLVG+wZA3NNmw+v
6g1vOZj0ffzGXAaowsTyxsy3A7fgfsX4NW6f8uyWWsL2xQEDQZBsjnE+TBccR6Fi59LWlh+5FiMR
UFzvJTL3wWV5g34RTiQmh7dr2brA3CrgLUtsafF9n1+LgU0Mh31GaEwuMR4KdDERkSZ8MupkcJtd
LRM96Po2QLl+FUGgUdtW3A6BffNmo0FpNO41rZwZFVAzEnlANsHEKd87QVsj62V2SzKWwCT3u4l6
G40n3R+8o8An3VeFldDmYsp7/PDp/ch3HSIO20G48ViG2NMRfegeeHyhXP8V8DtErFrH1GAIWfAS
I4wh/beBjUrF9pmohsyjRGP7LoexsevUsUKoWehPWq112aX2v27R4Gl3pTYyet9skAo+d7795Bzt
O7qcV6mPc9V0AkZn0xYnDjmEaYKsdpfdAZ6wby9n6Z/LgfV35q6NjWyIuV3SZ6ySkmXFa2JP2V4P
MTpfR1P0lu4WhdRwGuhtApBp94Jmj7bsoAniONQHwHveiPDWqvGoQWZ17RiixfZhsC9jMcx5pYCa
tMMLsEfa1M6C61qVcNyo18uwGMNS5HdB1KRUmpDhe4KE/JcVE2GR0qH9puGHJNmmmO/+qsk0uyii
vPMD5Fco0hq6Tnu9bpz1Kw6eb9fRC9q7mCM4IEPwiU+VrlYDvliXWlgrcKTocrqqLcfxZrdC3eSO
qI/pI2R/qy3v3Igh4G/LYAO4S7HRmUugEgSRa1zG/Fn69x0JXAN2lr5uYZ3h7Wj2qhb90QzJ+b7d
4ya8rIlpte8gRxKQ633YII+qxzloXhds3mUCu1sgA0UjiLQM2MthkQtu80RrCuMVwuNH5+NjKCJp
yIkqogJ7sWRhko6V8UM/Iw6BUKo6F2ZEvr2UzPhEf/IJjL5BiBm4Pcgk6OAuRtjDjXEsV1otavzL
xKgCSe9Nh45mnNlM8TasYNNEjZjIchnM+7U1AsKXnSBQX01663w4n6J5R5daU3xv8js/Ip1oI3hO
+x5duiR5+UMGFtZmyEwki+GoV5vnjitXMq+jf0UdRIAJxkDTYY6yy95pcFi7NWiZJkg6CEpxxthv
xDIKpLPAfLo4VvrRknqukwm05aYFSSlkPEm3DEZR2le4YGthcqFudfsrl+vjDrKSN6X8Abb+Phnw
nmXwytfVPDUOj60dEwf1IhxE4eOs8njIV0RUjaj4Tmd366uvRGs1UZMnCAa4NwTq6nisf9fEDuPh
imxqm+X8XwaGBAyCTC56AKJDtcnnWHlj7goAToDxsZNhxbqa/fjj+CcM5H5XSj0BLYc+SNa9jsa8
W7zR+z0zktI8Wo0O5X86mTJd+j8s3F1YlQ24AnMnMJelTStpyhxmJzRufjLAE7bLdJvAYPbsmYBN
5yw4kNNyaklp6HV7dMvNENRzsm3Bt0tHbbv6/IinGs38WsQMEunWyKraF5jAvAVR7ahHAXIh9UAf
GkpiMdz87xjPoAbDzfOlSiMwxAGZ1LyQXUPaxf4fO86XlYYiYueLDxyzwb5IOlPNVfbIuIPbLPHv
y0O5BEmjuZD/x/r5KpgCprqEOCTpODxhIZNfuIunpJpaNpvgdxI0ZneojjOL/96vj147MwKNcCCV
ou5WJ2JFbM0Ujaxlbl0ybNbg72mY4D53DR7piXjGcJ459kW3XxBoNZ8LLcNIXKCtHKB9dzpPzpdn
p0C5cfmSPd2eE91RoKiS/590drxl4G7/0NWLEGyCyHVpCc7tXoFOacCCnZlS96OP+0XdrNzFgywO
zEuqERDjpo/gpm0QFrkcsS7r3Y/Y0pDvPwYaG62QVPprcwSoLu6EwHuqRYxeuE9InGHnJ/7iEZlx
DBYEMLMIjpWA81SEGcewhL+DUrVSiibRyaN5s9hRdDgebtyyPYRJl5DOKA3FvU9BE9KNN0N0PFlw
2/0m52cYZkV4YAL0DNC4ngySG3WCiUhKtG1KCkxY9LD1NygXTw6Ht5ny0auPz8Ya/uhzNwJIA66G
U+TbKTM45/4nphaDTHUIrHsfSVv/tPPPeP4WMjsiFI/IRlSMarGqUbojRWTvISZexEx/268xumNC
EYEzpTTiaoXy2Hc+l1tbwJg2vt8g2UAK3Zs+VU9uZNRYkcA4z7U96hf4spQxHLd6/ysAfb4OZcX0
sdVnkY1PxY3Zt2SEFHLLFHTizviVPkAhfaDAbbEP0Qy+tmBTmJOm+UCTjZuwY8hvDo1S3+DMAslO
2gSM2A9NdUTI0GmBlbYCDpmCp+elAMWPwtUGgwW5hHi3TaKjVOYIar09E/36jZf374tEU5lUZP6d
l1X+2Hz2VZw+bysxfoAffdR1eNIWoTAulR1eg2NRvrdqm61qq7ReukQgBlYTZQVtWXkq29ila0Mc
MjOcEBPR0C5U28Lb0M4Ws6rxcu9TnGRU7Zf9WzMqERPnWvlkv2Hhq0UQaNHKnx03PU6mWMMGXlO8
wNYUSdzq9+H14Lzjn/M20+DspXFqXrQJLTIak6Q4jk7zkDWMcN4sb3RHkSHHu/skozoCgHZFxk6u
cN8wOZ35FEPeSx7oZLIIZBfDyjMGiizmXFUSmgvL/FCMOyv3dBaVPeU3++EnlHXRNfnXbje8MtRN
TosP80pVNOu63ObRZew5+jlQZErzT9zRvMB0ZQfl0buPbWNS/dZVHRD97gt9tSi8YAzQLOSzU1iS
YudqXMX2Kq7u/D3SxcGhwTrnwdtT1tRNdA687fc8WfY5LSoNmNlyz9f2K/dTt78vfmx21hHvIOZA
L4XWRMaUeWGpH0I6R1mmX71jOsZMkT+7MvSSNJ014pGyxGPqSWdE38nUYqvfE2nHiA+QkLxtPBuT
hG1rm/7ZrZu5x2bEsOV5GlszRDraUm2znM5h8befRG9FInQ+u3ru1m1Dq8pBrf697Er7RrbSLf0M
tEjzmbJFgoPAOL+RA7I8zuHFTanMrtofFsvcveHThoZrf1H6gr+DQlQ9D28Fz1fnq1KLaPyaXtck
JOYHtEjFeinkrpqdUtvFDrHGGdzy6HH6uU1sycjAcphFB1wHOY5WHPbF23qQJ+8+7rGtpLT0VNag
BX8mixj9x73GeZPHXQ5N/5iCSuOBi/YR03sFSprtdFvSEON9Vxg1DqaWTFLTII2ucyvda0Jtqchq
zNrevHF0HN1jbS8imuaIiy/8d8ohtG0ouT9bEaw2KID2YAdyGo/jyazmu2mHpu0qvYv6H2FhUZQy
zzP/NensFnZBe7glqPxiM8AfO4vTmb6PuRyXjmf9nn26Ak3PoRYACoam4hcHLelI1cj66ai69VBQ
NG89T0MRYG5B5OFsjO91Tr9jtBfDGOYosvzq+SmNBJvv98dX3mqK4S0SjAmnnwuIQKDahvUpT9fI
nC69zIuvz3CbuyHEFu+T9gr8PIj4pA2aDACtgixxs+k2UJs/4fl7u0yYI7B5xU50Y7WlSP+qoUmy
efenrcIrTuVVQ4bvwh/ZTMEa52sVnKKKmvb/0P7zsehpE4sGG24DX2Vyhrts53hXDZr2aaUYuC7M
ysVTAkh4O0fhc/CbtEmcBlcGS4RwMZ4uX80yke6jnDfsBK27stRl9DGRt8S2uTAS3fES8yna1tAf
3TcXOhTfqoLDTwyLRaYroNaBGhW51D2R2zXHuBc8+t9tEA/f3clk0gwdS8EknZTVyGa/ovfAfXjX
V/blb6g63jbRABfYGtYknpCA2AYt0GOc9RRQ2ceqzvW4P4hhFy7/5/MRizmCuvclxGofXfzoAaQh
5YaHrH+K4rVuqIwDkQd7gZdDBU6pN3TIJ61AI2g22ObGoK4SotoozaU/CVH/3S84Av3Md8N8KT6W
5DTsIc5YtpTAfEXdti7eWz7NOzbWxYUxOX8gh/TrDcOCbccxBwG8QmNtn8TfGbYSvhxqlukf2BP/
dVZbCYIvFuLF2HP9LLWlt0h3ldA06+nlaW+GckYxnTWIzsEa8IrJJPT3XJUQUqg4WuScZrPmVAyg
0hLHiiU8BhYASLwK8L7m/myQXX4NOYgmrLECW9MGaz/hTROkP+m+005+qV/1ndoKw0ve+36n7BP4
KMjTZHRyMAGenM9EVMUlZMhMI86D3aSMSUAD8/JlyN72HiqBfR/Ohntpnh/E5Ykkrb3IPj3GhIiY
mNvPiipD0N3dvOrouDrc25HtWAmw70ZWMeR+D9N5HVZoJoOWh/hRiv/kJDmXvnaqh12s6ZmgyYuH
NqZVhZKFulEoa9DggXK86s9JB/aCLEW+R1rLmkHQEQ9lO65brhvC+s0En1/zmFHA6vF36WYvatVr
8Tx0cxm3XAiWi9ugnGhL6LwlA6YG4T5b7o8tc8Ce0lrS4WPLIeEvjCgcw/dUrsDCybewNk9tZihp
i9etTXncCn4VxgpXo6VD4s904BpXXG5WG7s/O8TU9acJrWXn4UFmAcK31je8EhFWDRA1ndDxn9dG
3Ku/du/5PXf066KHwhy5XvB9ZKJpLZUjRfJmrH/9tdxNU1BGZTB/kpbQx6l33FA4T5GfQ2Jcsbl7
gFS38iTJnA8uw+z46a5sZ9wgUsoNpgh/A25OYo3qCgH9kK5ZGPSnnu+fT4ggfKDYYE5owpk8xhuD
BTv0oOLjtc5KBfj8/FoF9n4SB2k7g+71e1tO27jcU2JR+srVYvdY4soE9g6xJ0Kban03o6You77L
GenBgUQpBtLXK2mOIP+alfzS6Jb1NGWBcvk2ptQor3mVOX670ksME9ODFxgdmqLiiQqjhXloszss
u5hfKQvHhJq9AosA9rBldkWzs93miIP3gssI4Yqd1pBna8kAiqBUZqKrZ3MMP0MtaUWY4kq9EhZv
Lfrcys2+XMU6NH08SwgWO54P1cGmjSSoz8Mt2c5W5H1S1Ves4nxRopALt5pt6KLLrEPW8zAkXnYO
JYjQq7RWuBtZ/gFVRsdsj5dC5QeZBmJnzqGzmeQCgFBZHLPmyMdMbwKVVfR758laSqeDHtQyBJ8t
pplmxtz7IKRv6HItBaO5Deb4tC/u2gtOBrRe/0NppB/2IMaxW1KBKxT/RtlCasDcofCi80igfoB6
Sz6fKlq5O1ppXF1FcHPgIWF1h3az/F6G8pST/9ESjuelsobeLW6gejivIqgK22ZugAvNVg2Q/UPF
BfEiCMRFoDu8Tt8vU1BzZqPrV9dw4iyZ/Hu/HXcTzSHneLeasDA6U5338mX6CPBhQCNt2qv+hFp4
sHYKZwkFoPBNMbBt9fXVW0svK19NFsmTKa8A9NDvQTKcOnZB8I1BXB5qiDklf8TNZSaoqnjWrzv/
rPZe3Q9yvE0fZ5pc4WlSKIc6ksDCy6emCqOY3FBOc/2eChsD2bGIECtgEnsW0FnUH7mMDCNiBd53
eBEOK/YmIl+r163cKSUlXAxWwbFBUF5+UWeuXxiqp1cIB3n8X5PxljfS44x5HKA8u+dTSa6sIzJT
sXfEYutVY4WTJFjsUt3/UFbWmyumO9OdZBpGCTbYheggP3QKH+GHuXcX3g/VuiAcIFB7iWZ6oSPL
rvwH5Vo5tEgD60Tj9mgjXNIiaULXb3wpdyEwuRBRWa2hX/iTkp92E1HbEUPLPXYtCStIOGrxznYc
mbZpNPXdIz/fa+y0StUjx3DSmXw7qYoFZMIW7SqGk2H0KdlRbrQ4tHxQR9tMdZ/m3vFR2ZebUkUR
+W8XSQ0+5dicm0vCWvaA4O8lA4c5SUrFcGumpN9srWeYIkCRJikF4tgIuI/rrgn37xMK6hU2pYH1
ssz4TJXqSMvrrM7T45hE9qU0qOAQyOGpPM4B8LfA6znyBLMVw/a6PoQOQ3IIsv+gsKImBFRHJD4r
WIfdy39u0GKTTnQp4SL7w2p0l5Cw+2x5RXRgiE0SCruFUSeckKwIIiglnhGP3c9eE6ckQXH8r2Dd
GylwM+qhKAMRCR9YP7mELeOYOuU8nu7G7GPGpofgMltildO98JNTGWlG+RjvGW503Avn0IEEuPcP
dLVEm04tWFBh1Wb4WsddiERb9TpQ4ORz/9q8k6D+qH0hfMrsxYvbZLynMQcH5wDylZJN6He7Nl4k
6LSYNpYc4LYxZRtxUBAL3f+OBhoP+S0pBFzR3Z8YEhshymUifCI54fZlJxLGpdeigfp87m+U1+AO
2LS1vZLUjMTCSlDdu4rW7jQYggDiDM5XdL5WqjSD464U8wI++mli4M/ehTuAJg/UhZqlWoGxoanG
hBv9ZDHQZYVlpoS+tm4g4zWdJEp5ef9mXDoco/4vrJu1lAKBzmbLbdMkB5ejX+V8FySRYQ0r4Tmo
xH0jZ8FNYPCx9IwGBHEgraDaZnEkAYZO967gHhqEqEeCQ30PAbCpUyyHZfa4F0bgGHLu7AFG1ei4
V1Gn65qTHLv/Twj72VjFPHeeIOpqS9Fm9MQh8Oakk4070l6sR4HjXyMJ7NyhVsLews9bXyXhszqA
HqhIzDyLdSl0l6lrlmU6JO5z0Zw4VTAThTQiedYtsDljwWc49MEz0fhddtUNfgK+5M4Kc5HcqpIE
aqNEpUPmdnAZq4452MRnkjm/8nxfh2gu7PpmsEQ4go+wQv/e9ykvMmWO2MzWlfKOQmNTeGeVt0cr
Q4uMqaO1/AEJ2AeAHpHhbUafZbfNktV6RFTmpeM80w6bKqncRdqX3wIIkjekCGIFvi5GkIaTqd0E
IRchU+JwDN8+JnSqpAjAijrSyfyAWvam+pPpDFWbgowVGLDCt24f2puCsXtot9aubayuGA4xV9qD
d0ZtGXlIvUZ/SNVMB/mn2yhhGtq+SYE47MDPr0i9QyTFhZpcjljkDBTLOwylJIDgQW0mEYb2T+GT
KoAychj1j/4PTkmi7zJHL149urbPMfcAdvBzIbrXBuWRpt/0JhHiCAP6pGNHw9OLvlYrpiOMbpoQ
qqN2pGA8HRY4Ronmd/pDFmJqayM//PiEXdXG/16wh04L5v2JXc9byv0oytfaNJSi7VreShZa1mLY
vrwYEc3TE3i9UvbXlC6uEMYaZKqhj5eYIkIwsourUGEToloJlFqLTOeD7lUAQTfuXFCNa2ondbhp
ajt8Tq0n/952tyupAS+BKy8zWLRmECzsYECwaEwC1k6Cn1QI272wDrp6wr09Vx1cSSuMNu1JG4Wh
p2+bTUxZW+Omhu+cr15TJpZFPHyAs8cmCIG927+fkySDJn0yFloVjFcbIc/7e/5UupkluYfI0VTS
jeQrBsCLHrC5bC3z4JqQ+AVc5zCXdZGHNVQ1fqk7G2eYniSF+KuQfnpD75A/vxdBXEZuPqfsunyB
mtvAdKVjd99wuPOn0g/hQ/yH5kHBN6X2fs1AEMvsX/tyTIjoAHXn8SvfvLWRzibO8W1iT3amw2px
8l8TRsW9dV16hWmtrdOmJo4YgBBuQW8bcJRgeNna3alVRJZnY7za11QqkCg83ZnvUuuBN9ubNQwK
2TAp8vuHl0sh3IyK0emgcAesWy+7tyX3BhPVDV8tlEnYAUwH6nIiY9uZq2sXAOyvLNTBOtywX7zl
kH+Uj11vPzMS3pAN6nwGvxlc6NSrAuvaZKNRsK8QZLxH1/xyZGy6a3d9AL/3SuKjCRVNWRd3Ldkc
ck9TD225gvIacADho722vwgh9saFBVfSyAU9z0NX+tfzmMZHdAOOu4ob89RgEuHbk6NcZ8UXXTni
1Yq5dMlKHNFf004otjdPixPXIIYlp7BUXMd4n1VNBPgqcyqnWJFBqY5Nyc8N1GSGlcckdoaqmvZG
QRqt/x4wPjkLwJaia1QYisa1Fv8ifUaGUzLY1UXvp1f5BUvXPoVrG9dY8qyZ6zwuinlTS8aJqdvh
nOAWhDCFoUE5zdYiEWPOgDs/wq52gATuvukBRBMsiL8xvvJya/AfknxG0lJAq4Xr/Axkjuf4e9vn
kzleXKz1ODmIbTJt8TKJ70E1srd/KIBE38Dw6ReFkPA/l1qPSIztAE9I6XTAIccSzE2F7lrLEGyN
h4qbF710BrZLdBAcGK3JPbyKm/NXvwLWy5fR1gRMo8GuOXWxAbhO9U3j/aALXdqifWizX+Cy3k69
BOoZxkKMb+0qIw3OE+6DHoLfA6Z/3+CNTZo5usUHeexp0JPdm1MfuECs53XxZstNrrUuQ27tHh0E
tTSxmUFIWVGs7KpuIuwivYxexxJy5haAxiQhxQkgkqiFUXUdmF2326S+PqdVkE8fW1z3b8lYt/qq
FxbJIA8L/k9A5rERvJz8Na4YINbbA4ugtqWUWH2eKtTxOYgMvJXFD/FYnfu4v/KitGUs12Liv1AQ
YjKhGh3ZSk3qqDFhotzNO2hHv4zTvcnBlJLlsYh1zA8yAh6whY4kVBPH6wGiXsJAbd8gqkhGhh4y
AJTagBwCVm4/lsO0blv13LEpsLJLBJUih7ztS3CFXaNl4XqOxF3cltxpB/JQkh4I+JNYzwOsJ2Fh
KhS9OB+F8QYhhc/tjb38JkRwO/0piMc0mEqgfNF+DQ7Upa9l9abfUqsMyd7lp9sq98Z9c19tuDeH
e3VPOFJboXR9oMjc0YxHWVUY5WYVVyFgJPMXNKBJpzZLFm9blf8PBz6jREz33ZoWHeV/DXFDrq8+
logDrs6wuqZ8XD4OeBRY8goaLasVv14onI9uDyh/ocqpleqqr5B4m9m5vOjWtXIEswTsfcb+ZcgB
q6D/SxffIk7991wKFbz/BxgnmBRXln61VQTIwCXdY07zRdIEjcUB2RW0lisJ5BjEFNfD0Kw33Hou
3elgMegmewpjwiCdfvOZZjOyaJV8BzERMu5fpvanANCT2/veR1tNwCH3raYN77UTCNOXp5VTBxGN
TJBCLYpnprNdr/E3rF6JlO4s4xG83T1qLbAQyacXeb0hzoyVoQFoF3f9dXoOqWHRdzIlWHTMR/59
AeuZRaA03P7VzMzBlEpRg7QtjES9wZwdAHHRtWcjPKI5OFwfSyqWt37R8vUJpGJyz0eoNYY08OX1
MuQ63TwTsx2WEppGXcv/ad7A2VxFfYh24zXgfXL9acBaroOnDIFa0vo+EkSE4hjOsBkUsHiOentF
RlKH0XO3NY823mL/rIfsLkNy8vGciOyCVQoypIIN+E99d9iKGVb1HEAdvy9K4ARp01SLpJ3cf8ZJ
eSkaGafQAAIf/HjSeiJJ4wXIuNAwIoYL/ca6rmbp8hqLOfv/e/suQua3oSzAFe+9r5SZBPWGW/6U
+G7PlQzL6NO1bFCqjFsLJcJiZja98NgiCHpcp2nLnXCLTq7rcjQqajLEzxXKQI3iwC3BC94cMjeQ
R7o95J8VPtPjcYZmBHZK0rnWjjCwAx2/xKwa78hUcprbntYymdJqrGYoc97/tSlGq22HWq5T6BEI
KnCFhpgZ2PQlwdp1GdqMtxFkqp/twi6+AaKB8+JndauZD8kHHiMHXNxMuyYgnvQcpHCd2dfid4U4
SpqJGf2z0KvV91N1MSY8ghyejU4Y5mdM9+mYLmk/dG8GN5rAAhmKhP7NFFfxvohuGh53F0d64y8B
M5xwvxJQPOIxiyYhY+eN/bJrFmKP3XP/fpgON5HaFZX5THSQmLGEy7/VYy4Om5Br/PDmTtz55bkq
DwSbKktOzZm9V0UBDqXj8/PzWqU2WFv6HOujnViKGlkmB/sDoTRGUWgAmn05tlypJ5fmuY8SNljf
K4X/3fi3Dwvk6eJXinSJJHCxJtvVGm9q1Nb2+gp2HwPc5MlgQAq+jOcFamtYT2SMwUFqqrG0P6q6
VuoPdj0djlmFq+MQ+aa3SpHC5ABsZft2bLw3/1nkKd2Tw++jNHdD2zKPimxKMSs3Hyw0X5JwQxvU
fsG5XN1OFYA2O8DdrQFyVYA8/+VFLJO/aidjXzevlFigWrmN1c7z+kUK3c7gZ7Kt76mFuS1TXnbq
xmgvWIBTreJBRFkhJYWlVzPqjzOuIyu2Nga0PkwG6weopPyuuboBwGcYldoM8BThLjYCDAqk6NCw
KOGaLyuZpGfIMuFdV8+f2I72t1xaMrPSDJphHvMwBvoid1sI3t7plE6H1EJ+xGO27ouE/FsH+9Bw
ZZFxA0Zkc8CyA22Ph9YbJVqD8pdiLk8HcQsJ8AbKw8dmmYfo1c+HpSxpNfz4YBrqUZlxxi9uQiJU
Z13+qaBT6X+Kd7jc5lbeCrisnbmWNJaOEPav+c1u0znNV8CMwoGVILiocXYjmCjlA7eAzfRPUDXO
XW/IaerZuWysnYdjeE6DpdGkvsq5+Z/MTTCcarI4kt/W7xY5kcmCyEmMZgHOv8uGcYcTa906RXqA
oZ1S6Qj1NnuaMSJwSdlC61tN9sFudVKMSk7R35bnMSlsPfGZwBIg/5oOUV9Ii3W7rvaRyv5KDO5h
gqyHJ6JSaKAwKJ/I6zWLOEcqzgm3zWcBKARk1Xn1CrCLzVE5WI7oFIBIdZXL2DSyMk0WJ+3uqxxJ
YJgrO5KwLTM2NXbOgnyD9GlefQ7jJ9VJ/ci4XFkxkMOicFFCyoYQqWBfEhsqY+rPa9+T1H+8q7oS
Xizfsj5t3mn8LZqqCP4xcG8+xJcMACBdomosO799YZazPq+VgDkO4rGz8FBtgbN24Os074bg9LGp
vDNT4sSUhMP7Shx/JRSrGonU6nT4DWgiMZQOzVjp+p+Xu6HrnMfkTPZNs9LpZjTUJ2mpUFrLDRDy
GpH7ZCaCqrnxKIMnqivZcTnATGPnUbNtvtdZCEHqmlDkCOgqzAaysKxni5DGMtrI2p7NaevPcr/u
tFHdYqsFbolPrBnT+t30WqRBt4HwgQbEcMyiqzIklwzPhnDAkyT6vR9t7UG2bJEM2D0rLuVPRdFe
O93vg+gN990Hh2PXVPLOBOsF5ZxeNAhFmP1Xa0FTim+0xKv39qt+hUk9FX6Kp0/pTIfXPbpG1M+1
XOPPT0/wlsx76uBDh2ZiPIQppxyCAN/A7OMuupNKr4WywTz8UPqGwfWkn99y5tuX415uSys5j7bO
dthFbKYJrSwoCcaFuV+Ax8lt9gyybnOXMV+qX+mPEoQwvwnaeSApLuPgV5Hn+7ohFybSL9C98StF
1PThKiJQL9QJCXhsIgS0oi7frW9cSEcplfsnK3QuiY2SF8A9g3n2Con6baX9zCvDwYAxcI6Yza5h
nLAM0I26CKkAkv9IBjFOUz/VjKjtiIzTDmVyURHaStjMsFDQkvg7AlLMMpwPVSdxTy/c3oAmqirC
O74p8wZBHyeCI5frEMaLxjXgKor5hHmx8nZdP6VgNlRH677dyLKWtPDs3BmIVK3+/0+eVg6s4StJ
ov09X/N9eBdrxv6B8sZyZGYui0Mu025ITEPLmjgw8mRvQ447qQPAyKNd2LxlEpPi5X9D4wUkMS9c
eWtGCN0nH5AhNUCwl+XY7qIF2+s8KnynF37JPuR7AEJqO2GwrvRVpSqlSrvd302YOVsEImuwBBFN
Y+jKnJuIZ8+dhaa9FxlUM3T/m/ikjt+I9zjUzHeufALk/d6xFB99jjLq2IkSoBRo29+G5C7tsc91
JZsp1pzBLBTpf6tVV3tYJ6hgcRUefaeGdY1mzYO/cjGczQYKC9s7HLEvijxdbTwHOikPETjw5p8c
6KJtKcN3ScHLXHZCL7trA/cDOvfQWzfzt8+hpH0NlswYOxzYxjYdT0V2LtpCJmc25ZUXr7r2Gkqh
Vk6wxjxpOm6Z8o56EMC3rDmmNU0cNArEIFUD7RcK/ej/nMcHKsF/kB37LXqs/jVy5QFLgK0Wga3H
DrbtGFMF28eo7Gj/NPHyfEaa9vcNaHzZgOnP9eZdvJZAUUMKS3xCAOzifhoy7v5pm6cLXQ3IHXyr
OkYHeOF6NF4Zq6DexgziQqKjWLuprgv2M/Ewbch2hdqcYFZ4hS36t2q3FLqinuDFR+e/kTmEBNNj
VARxJUqONWO8fT8xDlAoW+RkU2cD41fM3bZGA/JWp6MLIWdMu3nAz3kOyQAaoI1U/fAWIFO0VWw0
BQFEkTnuZK4/6IqKvgZk/CAIebH4Mw10viBU/n/Nk+KpotfVZcQTRXuhlt291yadwHoGb2Do+Qw7
v8TDjYvYKWYpqcUwoqCWUdkc7oAUtsiWngJbMiV4gllNFQ9p5g4CL8F/oq8tjkiEszwFKbfDt0b+
mMyrUiD2vhhG4xxhxfd/EnGb0cGvnhPOFKUBMbYhHK+WGFem8Td4nwLRF6dkFxLIpDlJhRe+SNy2
lY+fPeZLpIJfdvtE9RYz2BZiVhl/EUMUgiZFH6akx1xuuousQyaezhKuCq4bvxIc8m+JqxPxsuQC
/zamAzbtabSALOWgEahw32qn1XyZETs0JbZ/u+CXwrfnts1ABCCIwlwd26j8UEPj92fS5jLekYvT
8QzrQxECvDzK/UI8IHQ70qCEWL1Y4hf6pGNUS8lCMBo2ClrHNM3Wi401YGPd0QYVhBuCqKDnIvmT
fsjLPOabuiPLzKYr5ebUQLJ6+kxnve0aD/NXEK1iMyv+zy+6VjLVJhPVBENs6IoyXNPTeVRexKjd
bvYwIDD3V20XiGnOeVN05e6gjxQJ5Qj9+MHL+bpwNTg/8zvAN4B2qA3tAwKvspQ4sHGrQAh0y4+L
3DgZfouRGe8GJJ5gzg96s4vQu8diZKOs2yCYbOyRLNJqOlr5ccDNcRtFUZzYHHwAu49eDrY2CgC2
zFIFKxBbIZhSUXx/df0KL1XPeWoDDo48XLKQ7Cv4qYTiFDcXWYWhcgNGL36+uDKoNmvt1V1XXwu3
Z5Fj/m/71tlw4CCUNEDNzw6KFkofcRcDuJJ02bsdS4Mv7VdKIKpgjQ3SdwxkZFhLB76NqSqWk2io
oHFxzF5SkPXVMW749Z8iJdxkG/6v+ChrqB3Sv0OcNlJLiyjd5itrdY/eIrb9oEcm2+3ihos5zIj6
kTcAXRkK8w4jr8N58/d5sl3bnKvncaFreQVGiB5A9cM4mfcuN0pwx1jEUSi4Drwbh3z2J2hadpHn
55bXnLpCdhnKxI/8N+mA5qvzE0RrzwlA3jWJT8MexB9m4bjxNiQW/9silVoL7aZwymoEcse3/l2i
DCJ3tlAkpUkXYG0DYi3h+zZq6xP9JKs9UeG4VAmC4u6LkVYzMopD2lvX3OgkwFhGVetWILinwzwk
jENqlGbBp6oWcbaLZyOg1q24Xv3CLgOJAdxCy0gZWkE5j4N3MdGn9SSBPYCbG/WrJpUaBw2h+BFm
6mJ8c86KV8qld7/4DjVQ4tKUoHtOLIouGdybAKGGKmyad8JBgn7TA+oz6DgBrOxOdsvQw0uxSGsK
f+r/tbdicccsHjZlwMidjcl5PSP8m5j2MxDC7u2FleqU/pdjN2vZZpdoOOsUJIA7zFLyQp4d/R4s
9+BJg6EgOWRyh3PVXg1d/umJr6E76fpQZ1TTCuMtXUM5sDZd1+s2Z0J52j+NYdP8+l2aIhvkoip7
OPhHNoUbBDv/lrzB8dsU+stmLYg359ydUFbdjF1ypRMsTLk2wncL3p8KHydam4204ORlUsIaXq1e
NiwnCJO4p3JT3ftceytDoWubXUldjVVnU0l5EOQv3fS4szv/FfD3TnNR1JPKO29PD0mFjbvX436D
6shuvH9RB1Y0BzTyQ3yWOTQ47O9nbG1TLP/F+nbvP6UXkcUjeDAY0IWpSqbdyVKUZxll0Tu0Q4Mq
ZeolgnK3fO8P+X1pJSYG9Xj8l8WYxqOL93UKagtG4pZ2Q3FCIEklp48HFz5MPml2x4J9rdYEo7je
cF0JPMZN1wZ3/voPR/9O18iaTLEc8KNWR+1YYh+TJDhMzpKU7HtmzbiL4QjtduU9VVuXp4ze0FBU
FZ12scnLa5tFOmq1lNr+UAPBGECohS4dyiUin2+W4XwT3wvH6/pV+rbSySZZ/F/HVx4vY6d6pQca
uOqZpONiH0lK/2UVZYchlPUn+uCiSvraQ+OheKx7znwbAVNBJV602EUWYer3ngEO3lj4iWYG3p/V
rE27UrCWX7JRM9Li06HyJpQpUKIIMxZjyBSU3nd+J5TP7Ml6J+yixUIb9+13oHY/4xUqf8YTyli3
n3HsBayyFcgmOVR5VE3F9C1k/hrZo7GMF2jEDcA7heb+F+pqnmG7xly70FQIRFZFGOK3X/1dPDBB
egFmW+58O1gHPatUkK63Yips5oViOwl9RTFG0wz1cgHNtqIx8FCnx8nAs41/RIcvO3TJLBciw9JA
9Jg6AfHZcvd4pDbso7ENJFZCMZg9XOG1MWf97OOW4jHg0BNIMEYYYWts1HBK9pVOLhJhF3iz21bh
0XNHljbZEL1sr5/y2chgWjlwuQeapk7hBNKeMsKGsNfGpOooqOTuos6Pm4t2cRY26Q4GAWTNQ093
xjxPnWXUZBmDI2IV4NgKIZ/u8bHA5+XfQItXrWyNnjIdUV9lkxeFbxqP9C7AKVBec6tryCJy4SZR
ljCC6eCVjVH9B4mwAjyG6covAb+ZxOeUukKfD5Lj6CWsbCQIfnr09M2CLlhoRQXo+cgvsexTcBHh
sVJUiDmhGtKyZL71Cejj6v0+/Q499rAXulrmnA9+CDTEYJB3cxGKXV4gfbSLPOg6J40BxCEq0SWs
N6LG/2jCBDzeff+uoYx/HQaIHD/D8/xO1tIagsCMh7inVNAKWq+Y+tKF/ekqHeCDnMnH+MLjHwTU
IS037Z5/qi+OAm+pWJRBPLlTW23y3R9nFbAD6c3szTP4BoVrbChfCYudc7Yxe2rF8+O9jI/A93hx
U5PEDNmpzs0ZsAweCoBTbW1O2Ng8QtGO9V2FZvZkBQB0B5P3LLHqP+U9QoiGY98Liph+hb2fpfek
bHsckvGr+0v2TsR8jSERGeZUjrGgh/MCYsMJVULn6Iw2qyriGEfw0mv7EGEKlSBEWB9HY4u3FALq
z64upequfwbwws9fwH9Emdvktg4kiQKdLZTXhO2GJUFqoZThYJ4m9NDcXPHto09pEpWgcJsqoAg9
szQeqScgZwXnYoasjnRV7i0VftC2MeyyfCdnqrVpZXNZOsorv8kbkGWmYjSS3Tm7fXpGX8r66ybr
VO/0atdz0XGB5ceRF8esP2GEA+J7oHfZVwyqMfNi8AQTgszm57I9Q0JcJPW0jzrlNveAh38iyu3X
8e8wvMGzoR5IBV485POzsqyexoV0xl4TdxtJKTN4gxafPownY8OKLgtIflBSGRrnvq5mcLRYyjhN
EvlIC4rLokz2OzWAboH7L/470FLCuW6D/wWg0YsIhNzFi33Sza/zFEGA2Tje+pX7CHSzPxG69ksY
/biniqf7TH7hlwzzudSMFFLaxotEpYsmCN4s0JTrSnRYswQ6RjqAjWhchLc3hRM7Mbe+u/zEYkug
dFyOm8u/dj6J9xhRqe/t/tCa0tmuKwd9Liw6NcWh6MCPp4NoxcgU4WODV/kMtV1Y531W7zsSUa72
4GTtN6jZW4k56sWPkMeJQd/3zEORmgkd4ofMC4ItAXUDm/oO2sYW4IjvhiE2EZieJ7bkdX40JrkV
RXbiJe/LUid0ZjByAR92uAB11mreMksu1/DDFMR7NQgVzEyWDEQ1TO42PukUh1sRM4r1m5xLgrEI
rFPuultuDFOHdOy+8LA23W+B5bNE7gtYIRQYRo7bhQ6P4pFK4UN73E4jPc4p8TzZbmRJ2dFmFyLM
60oNtkaqOYUhY5FmgDqOUviNPSdAxRQUIGs4YT+VoRa1fwydBRrr84UYxV+wXX9eW73jDrdH7cld
scgrF/Ws+TgFqWKJJsAoZO1Hlf/OzxL20rA7uwkJbmcmRKJ0iyifpUI9H9CrVv6HoMsDGaY0qMTq
Oj3Z9arJNwmbx02cm2z0O7wgZTHIS+1+gqvq/hobpDoqyJ2EM2Ea/Gd+D3FU9bw74Nfp/ibl9lv6
5DCjjCPBrJ26WRp+SdsG8brzSitR6ZmXbT99Xd7VCs8dikpfIrwLqTEt9C0q7Afs/tYYl+/cysMJ
Eb2WZsf0hO3KN8+gXRW95awuNTMGrggTzOj3o8bSpiQateGCrhIA9rEKvto/fgmHuTKSsN6C0V57
hnDfRFdEryVy3uQ2C0fEktoAchfl46juhchFTv6J9SnnVODhqrzaCIgNVIEa+NpYQGzG77/mqHb8
78haqnSQ3aBryyAcSMlxMxqIDEfLGybD54Hhd8TV5VphS702IApSFKqWgp7rFsm7CfK7NkVQIzCw
VH1jqx3M9sOi93g5g/+REI6cCMdWZEJS5dbpFLtIY9nt/yp3BHR20/NhecdL1nEH7i4T3X5S6mH8
BwNH5faeTVQZjnJydloOhLfuIPV98aVQBVt0cfpDhL+ev7ICA0zVLYUkixUXuKlkNGmPUaH+pSiy
3X0e4hjywzomO6atro/qAJGzWIEsiJsc3dkc6qm8Ycc+CVHFvTdvjUVxlgNrotuCZZcTOHWgUTto
mdp11Ulpe72ngrl12tqbpOWitg6fEBVxxwMmDYkV6c7asOeZi5WkpfbdPHFhCtBuy2N7kibTsRdf
WxCRMbFmx/gkbTVX+qdXPwxdNwzqSd19gaIyHWCu5NxUa3JitKzx5OcxpmejiS9oT7hVgFxY5K+l
ZbqRWy+NmN3MYjdwC76mz8I4qINy4WBAjr0bx3jeCu/DOi2SGC7p5tDhoWk7BRDlSzRbr9elG7wR
uipdwQ+0F5eBK/A4kSqdqVCDTslDRDVuqD6LGFA98hsFF1O6phYNDRLgps1rZUmRifn5p5OX+WyT
z06CsMRrN6GCLQYMBDRAUAN1hA6QSf16sTDyshRkayns0wWX3N153bnVsKkPgzq5a/J7+pOfCyym
pqUb8dP7uCvpdimXf+dGACcNa0WUaLhXYhNZ6KQeuDtvKTsEbF01f8AC/XNzg7va18dgJvR39ogk
VysUsR9TyB/M8Cd2yc4yw35jNQINOhwY2IyYcWlBxBgm+K37ZL25C1GIM5PWAZoEKijimHf0VO/4
tzEu1GOJAtWEu3ron37DSyV7E834jxVF5B3R6t779SXw7mycuX+5/NaLZuP8clLEFjF1ZkPTEpGS
bpt+fpIM61AwqjG+OmYrVHlJPykqOO/FzWrA83bdIjkC5Z7b8QYC8SVUnCU4QZlidnxm3+W+9qm9
ja844g241NXTRcBW8iYVzVEinPwIgRWYsq5H4uj+9zw3HpZiosF8gRXykOibrHU2ioreo+u7n0Ss
fQ4EMF12ak0fQsiR/+wVUvbuzd5o7WQrMTreLAK6KF2ONCaO+jqwwQHdTbo+cN2LViaNVyRA8de2
KGDyudhA6BWLRXAVpVXAta2WvWRnDygpNyY8WFgA+iarv1W/CFwqMMQ1BSJhn6nFox2qvPqhD7SD
HhJawJEVUVPYSBoShLbrc3JjlQi2M86pX5edOUJRjpZL+0ARPv65wKnj6J+M1b5RGY7oribitjrF
uAQ3G2ncIeawu+/JX2S0zy7py/odyMvEF/QNltGosAUX1xNPkT5uaEWPzgPuSAZAzTH71eGQc/aw
Ih/2bPSYirXNzGWIAO6HnxjpNaCEGLpZTTXhx84qmjPuM9Q0pGzl0wylLoDOZadTQgIngtNf1tjf
ZuQWva3iiDHs/zJR/njyWnU5XkWZLHHVPXyimvDtpd41dbIo4JfwVPAp1Ye8QVOuxRz8oYa23go4
spXfwYe8C1hgPSZjX0KKkAhpd2nxRvpPA1z1IEKdzZ5eJR2WLyJEClna/ajMWowOw2/qwdxIoapd
Yb2qbcpvPRFJfoviltPLiW+V+JtRCH2W2UUrj9ddoLx5PhHPF0DY7o5O8fjHRtEN5maKMdqOJTTQ
vkuV92OUpmIFuJDnDiMXmX+wyMRzG74sWaccMw4Urt1l0gLRaUP/vRr7z2c1McjkQXdtSHIlu3WK
YD3kAyeK5EAgsaP8XAm5gngDZYrsp7tJVbJ8ANJikiyKY0c0gTINBX+ZeNNBu8J+Ow6CUugCU4U7
i45Lw6MTBgUtKHerWPWw0dZlja5ELZ6owWQh0Y50RNESmTqHKfg1iCtyDyLqDtngMKFJsbFaLYFq
VDjKRposJSzuLgGSXfCAauYb821CznZ4d4A21Q9EWcIsyy5IYhHs/X9E7pwODBCSBjdisQ3QHwgV
MPg6JPE5fFVBJAYpMLHLjJJ4t36Hs0aHs8ojjKnb9lJ/zQspvxKaQEVqBsI2BFnBQIgQX16n8J45
hhaeMgUgAXS/BH2s6J7Mozpu266f8LatGB6q3TlFAENrW2Z4rnlobaazQZNVvMjJYmqOhO/IF9jV
0FW4OnRrgbJOFHDIE30eA+E656YpkFTFxi1fqQz7gCPKx1vJsZKpboQIXoicUabG1CVJr4JdL+VY
O3xzLwu8odM/Rtj1KxDfFtvylZYXkDxs16hy1fcmwbe38JlZ86DT/sAA5fBdaPCtREtFGDxC5mFw
pOW9iPJvUlbNbwWlRqjNlvl/dXgwn3bgtAXryYM+NJTFRDEljvyjuoHtHVkhvR2+GaeC8dm4I9WA
Vkjs2deyt0mpD+vxQ950nsQI4m+uDqr0/qVeBqW8a9Snu6Mxre/FvOR7PbfoYJXXI+UmO/1oZ6g+
0WD/ZYA2v/7xL8UaRn7JyFgsQ/0RRBHjpXafhOQD/u6IBegpkeD5X4KqFZZrx3CW9TZs1hcEOuID
fL2kmJtK8xzSUEv9KuE750Jq2FXk9aHncxKe5FSvMiRj10EHK0kZKMTAImGAZPArKIctlg0rRrC0
qGsKTaJI6m5zW8x4Mrx0sDqACdGZD0Y+hSsw90NoAQs0OLLJF6i/65j4mSCWwlVHZjJTVBHe6Vpm
mUgA/ZsMdsRjXW8QFLkg7xKzUAYcwFs3IwotodD+DpV8hRep5TInySwahkilX501fgDDtCVG6yAi
fS7awVmgyCNw3DDm5ujVLEC97Pqsle556/mSl2vkSvDkjqX0/ss5ecJmSh6G+zlhGCm7gC1av32X
OT15mqT+4PQ1Gz3xJtJznjJXuMLjX4uZqR96kSyZecPqSf6Z09m+UtyPugXVQ5rNDkULYF8H1Dk1
2wdbuzuYyc5/7Jh4o4/8tfDEFd2ckVIrZFbfx1700cBcsfcIvKMIFuu9FBAcIs0OOGXKNqnV5BqS
JRPFN7vmsqAroF1AWp4cNZQTLQhOh+EEpbUAJQKa/MWiUh93kP+7S9Yj4p/CnH2AkY3e01RDdSj0
duTdU50J/q1goyOgF8ZG67h7UakuL+QVk8Cks48QggVcZefcZJ4DwjQaX3pupBQnBZFqZRLcMEvj
MuX02tS9ZNO0m6Ty8Vazt+E/ISoRYXAXgyWA/vxD14/V18Sr6AAn/a6z8zXvSJIEB1/sjuMFQQeb
maiAk8ose33ICs03sLLkVvEp05HffAN/vrmrRjA4vqGCBbFVeoeMjvaWVHtTMAKGoov7ktGFog5y
7QZlIkdKnPYpIfYtUojNySkudAQ9pHboORrxyj0YkpfUEklokYCfHllKf3jTVD7XRSt09nxUi0r2
So8yCNjGZMC6eMtFTGFan2QQkIpviwDG4y9pL/nBrAs7/i2pAKooi8zyMFww2FvQqqIP8uqV+otF
tgV5TJ7sJ6D/EmAxNbuyPm54TlpVe4MSXX/SGCahVhbj28cM5bCoaPKRdYkTm6vD4PLtW6TzfddH
vjQmqFEGhm9OG8vLCAok3grduq+QlPylt8H4rC5RE99Dm20BXxLnBhjkvP8s96wWWkKrJs7ei/CS
fxU6eqZ79W7ABmfKmwcZyLPekwzvTqTqRitoKs7ImA5eggIpshoSx2TU2G59fBsTIs+fM6vhRweP
XhQ3pWZFXgHRNoNFn6tdJvs1YhY6BXfut0phATLEKpEqNcc4oN35cGRqlA22QDfyFe9mu8Zw6zMs
RAZug6enJOjpbnvoro8FRJ6qq3r1bdmf9hpyFZZgtihSnJF2bZS6LbzGYyjro8gD9f25I7urW4pk
9p1jm+IlgTrDZeMPWEeaw1mPlP2kOgO10deqJip0h/yLzhZA1NE3C8pJIOYE0YjUTj2duDXzIud0
JjNDBTy14mSRFJBA3Wgx3hy3ftNa+GZmSEo9roxzPzLDgOCiUUWtJ0tRH9n/2o407P2KR0qZ+3X6
UevAmzYsx9yCyXQgex4OnGCz0pngGTZlN88KApTaiVPrrfXvq6nfv5tVkaRQs6CoUCFvXVJ26rYL
6XDP3df6m1OMGsr5Ir/5VOHxIz8ipSmKF+zHr7fWjtWJzuYeAWzZQrQXw0t1DKCEz0uKwAdFBz57
NVI7Tm9c7x5CyeLpRRuytt/Y1o3OTVffTzHy/t/7wbDbVQGMPDpxpXit8X4uoff0UNlkrqLfvw9Q
x836AZKV+53+Sr9lHe21zggdHJ2ETuhswAVNnbx6DBfgWX+D4izbNnj0+UP/vmnxWawGOkwaWU6E
uWxtgWVV72vz3okWH6ioTVPsfQNLZrfzgZg8NFQIYY5W1ngP6wkEfw1IHNvFf+Nk/KcNUGwDtunA
78F0AuN/XFuopnu9p8ZWYunvidoOXprEjU8G1ecIbjIaXf3tykZPCbTndALLHAJuhCYipP2CfXbL
fMW9lEttOeXhb5oNNqp+T4FgTpaCcrXOKu8cP1rrLVZye48iUvMVDSv+VXyj97krm7rNAPhLmrLI
ejw6Tlyl5PS5rFAh1jW/iiHR/mGSEocPWSILGtmRP3jGzfXz91eahi9dz7/2xYVar0asdw/xMlFR
KR1TOXNeRTDCcK8bMtzbI4L91SnlJJxRaUeQdxnd2kMM0m8K80YOt8Kw5CtCzYWxsDZqILUWHue5
qHyzaDLuHy0OV2X72Vnc9yW2WCSFgXyHy5rqZOXh9/k4HYJsj1LZy5YmqkzVIfIp01UfScTwAgFR
JvOE1HS/T9kfKGFOZx2Zs5DbzhHWJyakIs+rtnd2JJj3IXY2qRW/iYC76kMkYSjFmwLmGWsZriBW
yoUvOUUVW9UjFbzfqox4PgvGe591njAQtu1MtfQNCExMmKP/NrWyiC9Laj2JoLQ3XB0uuviF+/u4
GjIZ79iEJO7yXu/rLQJGefRX3ciPC6JuUO6NYT3eqvEIGrrR02EQOgRXaudBeKZy0mk4nppP+s6d
lq1PDQNAoJeToBnRgOg+QT48caRC/iVKq/8tQpHb50Xpy0hmhnllBj6FR33UVwYhvCKj/GLIUvfE
YJQlK841xBNmCn7it8akMOiUykNGpZjWpDKI6z7B229r+LPxwRtyac63qP0Jj4yECxBGdKsONWa7
DsEGtt7p+7EROGZpFY81mupCIGUDsbRNhikj8u8RXNTYuKm1iSX4T8PVTeBgM6WlbSXJc/3olCRV
kyZS9qWcbrJCx1/37BZEoqMWLvpMWflueD1jAg6gwNrRLFUHL9S54q+PW/FSOlDsEdxaHvhShMqD
3sl4xYNCHqF9XkJ16sTqaBWWtyUpjbIrstEMi0i6pxbZT/cXpIEsQqlTHHs7QOgMoFvf9ReufPCs
TlWUljRemfOoVrJ1iNN9Wjna5DqqKB5eHiV9R1ojP123Jv4vpyLW6XvY8tmNaKIY5ELXJPvCK/3R
V1z4djm1JO2DCRtEmF1A0H6uoXChcFdbZwa72fTwLNeVopSOcejrPgSTEWJ4obf5WHPAu7pjuC/0
HkkuctAxnc5y9xqzAC5BibyX23zJKqX0ucWu5/7GhrdmvzapPM4m52KiSWVJBNbhhLHlTIgj5ihX
NxnDIIfZOSLUopwDV9ZZeq8cpwfQLsgTZ1chfcNH2fJM3ndAEYO/X5xRnnDB/Mh4gw0Tdxz7rAUI
QPCdxY8IRIetK+ymbJ+h/0Rz8hGz/WP3hphPO1mEtXOotvyDSmynhfh3fDHrb1qE40Q68z6BFbK5
D9h+wPDbydx1nK9J44QmiePU4yshGxTJqY7O8otmIa22WVIWwJ93Vfms01XsM/aCY/Lbk5nTmvX+
vaMGzXOi2YkKt/ptbND0KWMfFHj7d3u9WkkqhCXrPJJKn/nz3O9ZL+NWP0HF+6x4tz1DCrp0BEkj
g2Xf6oZ9L2ksCklv6lKPGcQIuIZqUmCVzk2lWPpj7qTpNnnxp/UGLntTxVO/QjF9q/1ZiLnc3sSj
pcFb9jNe1dz9jhD5tOg2FGlOm6A4cZeiox4Qzm/QgfmEZaGUP+cIdrQ5BK/SdlQQ4AmUII7WzhsN
gFkGWPi0f3wkf7kRlCMCHZfmpfKJSvNBY21xdFdlzdE15XPEMaj8qu/PBdyT8v6GPGawqZMoU9/b
hmeN94wCR1k9uNfZw7QumZq2MS+MlbM2/os6j7XDvx7JvquK6GhqReijCloP3+uS4rYKVroMyF1m
a54AMt5JZ3ifSh7/VmZ5nmszTvmoMsP8Tsz5ExdTSAxiWneMphQugvDROtd00QRhJjwjoDAjpkEe
vk7N9PcVvnPyVsPsy/ieRxRgbrWkisRw3+f5CuIWFtDoPdwrt0+k0XISKVxTjD+0qionakCxEOlX
ZPKTgJUNE3rNMK1himsbAojJqUHhI2Q1jCap33XZ346wV1mDqbcVR3AXJvyTA/osBQT+gkH5uOPo
CPAdT3VI57GZBuLyT4PjhsOJhgiviZ3xiN664dtdiFu2UdQuQyLMG/QxTCVwGc+fUrkDNZaRUAnL
yRW/bO9p8u+AkpgNsnXwkJ4r46oU9G9+0xpcSjDatt3Vfo/yR5XSWY/rDTZuOiSFlkjeN2k3jyn0
5ngeV9OSG/6eHDxjsnLo25b/682t7dV3QZ2gbx4tc91yrNMb3SzwkhTMY7WrJB0FosIGHGnVA4sY
/29tXhOrxsISvfmCJ83mg5WkPlPhiqgLa4rGvXDrWdCowBWZK6HlHfosMkf9qL2Tz+APAJji1ngD
ar81DjnEDTYG67dx/Zcwkr7rY2us5neAaUD1peJqQWnxik0mccqjbbvD+hVcAK1IS/UmvIaV35lN
gEJCY//76dH+0goqOXOzofwLd1hoiC4xxZ34bC1e7LoITuqdEzmIZ7HSNWGp593yUS4joAI0SJ7j
5WDj4Q3huQBc3e6DQM9Kvj4EQ3Vw3QfilG6G5pjEjEXvsOcwq1YPAR6JKu8yTbfb1bN2Wpr1sU6M
7ebdcE3ApKLw1h6JMrJiKf7QKElqDsmrJmyuurDv9/fSpjXa/XUMGq/Q++YkTqJA9Q1CYMAErsch
VMWR/Uj5lJo5LBOangd5+gJFjWy5mc1JKdVPip0zDkGsNw9xh5WgsX8yDCnHNh9ZIZlrNRp7szp2
1kdizGmDNGR8AvJEdSuxdm6aq8AiWXnzttDNn5coV83/Km7DZu7LH08M88LRGZxBuATvBIqGgls+
K2C6S9HICcPW+p0nnxRRA7A5b6n5bagIScjXCnMHL5+IFWaLsngTQliA+ejsuOjVEcSqk1+YyAua
IoXsOl+SwrdQacxwhdeHszPUiVeO8Aokw/rTiKO1hDdNB86bP563myW8z7tKI8QgBCJEoZf5HBtd
tudJyl0Lqp0QnW9AaubJlQMucvkLbbvHjSV+MDZ6pxlHgFFF9IYyTPFkfmWh4vP/f5d7gyNrtFXh
R9EgaQCV0hawEN3CYdb8R7pDCFOg0tx9cXYv8AZtGEEM+Xb5dn7ktf722hg45rNkApGgS36rJnI+
bKpRd0y9guA9b69Gsyyd4KomYwHHzIhfpRkI6vt48AKpufSOHroDNYEeOW8VHgPaJdZ2fc/yyawk
QZJr+UnfB8wOo7LUqlqjAzBU+ylmsD2D5Fagu8Fbc6GrwHhZFVyeStTxfTzaWYW0JLoPT+rvBCMH
q9Z7rhmQ1PKgPGoDfOQTk0jktKKW/m5F8LZRHhNPon/9B0BfaStHWPQqn8bsQfZiViBXdid7XHoC
H4DZ/AEmnjvzjZClOrPdXKVwwZiyvQIhreDWnzkgbkvVNGmGBuMdG87xLZoTVPIXsF/gcvuxFVs6
O9LlPA7GdFlzdWsU+1tS7SSFhxaZWesGm+78Ji/Ak4EFDUy8I7K5gXgUNhVZBOEXIrLUtBaV/dtZ
WaPenIcS+v7KytnaLLCrSdphL4sN6N74As1nouvk66FOyUSbWygyPgMoOPLLov1RxgWgpOEzVJkE
63ExEntZa8POsV3sM2IQAYZRPzw+Ffxrou5CYmfn5EFte32PENGk/wBO7FYmhwT8KirZJESGVbh5
K85Zk8EMbLw9U72uREvwzfr4JTFM+W0IeTiROAiS62XyKe6G/AfX5WMvjsf0i176W7x1YzflVSsG
p72rQ+AOidRJq7H23WmEaSe+sR6sMXt/31y27cjU8XwF1IGt7qQn9aXsYJc0s8mtNsuRbBZWSTFs
tUYYkC86FjNq9xWhE41xvmA0nhEZ3LYp7Tk2hHx+DytVYB+EZ2DjNbFWqTv052zVpwonxHEmm9Lq
JsuBCTaGrK+bbGP8yedRukzzHucPuJiCt1p9qJUQfpds+KZnX4eNajmhmlptheF+gCMTwPd7nGqD
q32CWqYOYJbECEBiqsVYzztddwG/fVSEP9/XtsGWMwFhsaJd+ftFx345G3gYE47SHgk0cslFAnZn
zb/airyJpwnsKtvdpO+mMIH2mSmWF1+VssdI0SgHDUsAYhql0sN4VrQSGEZKKqcrs7BnlNmQf1D2
F0qLddKWRC0R/1MnwllA1Ic+o2n2tantmsq1GAqCFogbdtiqinboI09kS9cm+B0dlptkwBIFZiFG
F2CscgjYTMVakkXCug6BFPSBY+aHyxDYoaX57Q+RwNvb4UN73mR/2odYYmw7JNQpdHT12Jhgu/lQ
kJwpao0F0aPcuA5iN/okcyz3xCKf+HUNccd6fNNbvU/rav7Z+tlw9mVqdcDitV3hP1No9wBVVR+r
e3gYN94snX0bWJafBRov9T7gBIt9HeMbdgHjJdRuzhdxseWRauGCniaTnND2Bv2LbK4AiSmxgXtm
h818k/58PkdridXe3dSkqY3S9F3aKLcccZ1SleQXHWct3Sh9u3abaw9IaHVnXMeOzxIGWtnC9GuQ
Eg89guQzCE04TukXawKqeY7b9pqRHJ8v7h+IGVxkv4+7E/8P78qbT6fynEfaHElwl//rYpXB6Z72
9THrEkx52V0dwlzx1IWE80zs0Q8v9dXo9Oj6WJ3GY7QM5n/3yDyBv0BLny1bAkRAFqMQOKxjyKSQ
+EDEmyznBDZMPpJ4ar7N2Sff0z9sj5SCGR3nwroBJTWRHREUX2wmhBB9FYoaysPXZNMfOY8FEQrz
0rJtOnxzzuyqPmH5tEhw4zGajgBVDIMy61jKR40CUhDSE7JEf3iTz37twde7XtNaahcaamnXVYwQ
bu4sOcWPF+RVI2CZtAjkVfwtOtjM9D795PozqzmHcYrHZIsohdZPmOlPIEmBm2IJ0Vr7ovlBvr0M
yZ7YXvyA7l8o8RAPR3HYwoYBRTZm7m/MZyIYdr24al+2aoQCFgJHx6+gOlsuYGaA6nmeTaGim+Ie
Ekqr5lxJBOuUJpykhngRKxurmB+msBRS17Ys4i93IPIzFhnYhRCygezgLMjg4RPeya4yVuSURsRR
CzVdYBr3tVIvtVxUi3A27lCJvr69QQZ6XpLkcI/KGHP9Kn3e+YhUAhYIZp0lh3cWV++x5eNqTH/d
58WnaBOxqjTxRFKsZIonydcDU4CYBQlWNQsVX6mL+k14v7F4IlA3S2hyUav3/0xgd7ZD2v6I4E8A
RDMIUDA+fzDdK09r6yPzL/tU1In/iLf6j3yVrC55wzkeIsYG3fkKItLfo4kThKxNFfRWaRmRtxtI
7dK2ob1QZsiSXDDCwfj8acSC8k9Eji5MwPpKHBhm0whC9TtkEVSQ77p615KZFW0Da+INhmWJxzpm
/MA0Zr3O8uy6oYvCwDFKSX/4Xt+HXm10e575M9wU1kxBAf3OlshJYVZ63HQjsMTzcKIYOh3w/L86
UCFOaq2iTAD5oKlZza73DwmjQrWYMjQINTCh6E5pOZcHL3owHbmtodyo14TMTMmkbJ3ycjx8W4j7
W6keBvwBM78lpnDYDlHGLA5Tw/p5UkrfBz0DFzK7oHAWRaYozZHuPcfc8Ng9eklWD2kT4rQy6+GU
amYYwhQDD5GwXow6kfZMMKtEHVXhsDLBJxbSxgqY8rqoaMJGPixXZAB4f0R25VttoBLI1FJXtMmp
oAdknZ8Zdq41vSvPhedbepvpPSOkX3Q6YmAs0fwzfd1ER483YJi1mXHPbCByT2S9NgamvvEJDl3/
/Z2L99WdpQvaEF4J2irCXCLwi3v5fqDPo3HY0uhy2hu2T+EsM+cEaHl4hFy9kXtVAa+TCicPXs0B
2KjCkH4anNzGx1FrrkN0LtwTf6aZAdtT61dNaTrLiOZxG4cTy+qd1Jc3Rs7zLJH2t3q/nsHiWobq
0hJM/DBqshAlNzMnMWvZmePPzVIzKNBGxCheaNt6KeBKmffHakA7i+DLQnNOoKAWtvTIPjgeC0wW
5kPl+MbsYHPrxNmHo0kgIGCYUwVfjotlIVbsJ5CC/TCQZaUaGRX6aQjsx/6w9qCvNg9A4Ahl5QPa
Cgsin4rz5dtCBNrzShqn26w894PT/p8nbOJQgecBW41gBLojj/JExBgp47Q34L6awsMHzZgrIhXz
OZ7lCoXgfhU3D7a08TKn0Lj1Zuwb2Om1rwtqfZ2UygKPOEkZ9hUbGCrg+A8+ipb28j/Tfvn+3mFN
2JmBP82Pu3Q1Iwb9NnKWewr3Eirk2EqC17QK+Pz15uZHxMrGHfkJImdAZb497+MWAu0K054Em8f9
xDPbvrpKGRuORuwoRDJ07uyUzegWuu5W6oPiIvKGai3Z7Of0AHtMLSOVoAJXUdTQmwfvsoxvHPmQ
e25NT5x1L+8sKk+r2Nyzpc8dZVbWXppTTEYtSznAo0aZFoNs7xJEKEEtY8h1tmecKuBsLHhi1XHY
Z6AWL/UD3VgLrSK15bOur9Sww0kRWiuCHhw/FWgiY1De3bLAtKWzFnb/mDfA1YkbG0I+aAmBnpjR
lr0XUoORkxcn/fgpL3u0pN/biAo0ApeGDie5YYI7pksWNewjiKuYPSNH7JstlXTxYun3A20quTEL
rBgDzDwVyeFeYaH50YU/vMLLS8RvzlZceRagXTQmrKzufwjaFTveiDpGoGIiSGpav9WCZsBH6weP
fqcf+YpCdpqfUapvqtUFNGubCh4ydHclg6ffUBvpCvDGHt41W4Qyd+fX5tckLeBAjaM1VqEq5kC0
q3uX7JGyfMeb3sB+YQCHVLZaszAWS4DOYwt/JAsl17+Z49St+bM3LvBgOsY9CzahSJqRNQz6dEcc
FiHpohfXffreofpgw05NG95qz2GoSHkEs3tpdiWO3dH6nqgr8lFcEwAwFJxpEbWCYeBamMzlSAIj
Ym6jNZ8qzKtNhFJRAQ2lZNs4ev1z6E4JDJ4gpoPMOxVLhB3sfC+L2fdB3O9CSqZNFaUoAaAIV+C0
7pgjjz6qZ9N+eJDJKx+Bujn8G1BXVU6h/cc/VOKcoCVs+TiQ35NuHHNBjkgx89mOXCHnSoBWC5Hh
IFH8PcRPO4E1klfte+ZG2TyD0jUgCT+nWnXS75yNQpkq0sNOj/g4mbI8bsOpHZv4Tn6g5Wo+41kN
+CZ0lU1VYqpWH1yb65kjKdS/8vmTQJ6VEcZEMS7kTEgpreBAuyJ+oqyjW62UPppzaNB6cyFX+Xcl
lfZNoJjtcMM8dZY7Pp/fqACSTxdS4zAYA8GFETiyeFDIxK+nzf7ja4uWY6SdWnA4F2g6lJnm4K8C
puow0WgI2R22hjqC38yr2NFRrhwJ0/BdxEI+HOxLaD4phwL6fk84AUmhR49cH6BU6Xc5SRtt3ecN
I9r3pyRjRm3COMcOp8s/kglBeqlV+NwqwU7vBPr6U2cbZiE/OciQ53c+sLLFD5xcpbUxvj3BW1v9
d87yDnv/euTotytIQrjwoj5hAhnQY4ccdfu/rFx0pQDFr3pw/SvuR7pCt+PS4oQEz4W6LHuqENua
8Tl4/lpW6qQpe/JsRnzJGghfCLPSlbOoJ1scfs1OFS3ceZJQL6U4DWUJSVEgwYItD7yyAeGjYu4Q
7i7yDek9atSbXc1x5K8ypq2ZZq4mxJrxRVJmiXtP+eUO6PDDA5FByivQByn6MnV0CFsoxRpQ/pzo
nKqsS52g04G3xVyzq7tR2383371ug1g1Yyf/txTpr1lV6WUtFMDGFg9zPTmSKZsZmjSc96+Mzhfd
MgvEzZKIdhz7OKZJChl+xNFQDtyE1ATqMAQXXIXwMBWTHFtL1Q//i+rlwMAzfAqyS65iUnsT09Aw
j7Le3piHq28b4mmNbTuZ4idkADmctA15mtdKB315/R+0HxK+I1sh43TAcwtG2BApQqrwXNIYEfCZ
ULZkCNvxFeJ8XMr3XSZBEadWQt9sTm1tCEmI1IMpODi4JpJNNvuOPbr6zhF1nsCYGClEhPNDHwkQ
80N3CmnBJY8hDBj8tOvB2V/NVWdNPP0M4xllvAq/muuKMfsOUbI9Auoe/1TGT4bup0+LUCbo7h+z
mzaoMwKT8LpWvUZMZjihfAfAA+NKiet+dlQ/j0JORkFHXbGcZ8SoQVCLhbhcewZNpbR24mHT6QjD
Tad4oAZYPz/aeqeZup9mjRNg+4sWb1CCY6d7HqspvTLGY3Cz2dMOIZxUbg7aiOHJtDKhvTjQhGtp
LYNvqTyHY8J5vP6rjc2BNULqopLYk/beGE+NoLqAPRn1L01mLa9tjJPqN+idjQbLd0TZgNNVocjl
7lNRTtPOyBD5XfScsoTJsmcN3R1FeUbZTgcJD9mqVbV9Q/Lp/9FbJJ2nK2oar3uJlcI9F639uBPq
ynIUpaOhjeYY3CikfdzyOFdCAAHEMVaKA9M5UZWK1+5b1fN4QnVUKK4pFPpmaz2ecvgQB+D8GRWy
whz3PBiCOWl1YNwYVeRhDIBhZaejson7Ey74lpSMH4jyAi9UHUOxwFdMEM4DgVs6WeHnBQtD2Wfj
OznFOhcBN7FngHhlYp32+b3Q/1btU0hhHUA5w9vOVTylMy84sj0YSUJNtxVZtvEdhDGu1srFnmK2
brl9JSq++UKK3gPYRBQSvTqjUzpyY9AIQNrzGQf2HEs/SaLDVnoVJ2Zlmv+wxW5k0kxWxX5utg3y
OTgksBk5Isr48L642vNKEz29Dj1P4d91lr5Oo4nLDP5d8J5xnyJluwozuGjp45+6A9Fm2kYiiqBg
rSXFeK4qdurtnYkebrptA7w3pVxhYAMASoTqHtOThjb8QyyN2MxKR8PMZmQVs7SSd60hvDsnqlqx
BOKDi+rHZzcveewDSLR30wLdkwUrzJkFZRNQWx82g2wZGEofP308LFcKqHRNgSvYdx6hySiC2ZGP
SUM5vE1/HSo7VplEqb8eQRbzYA/cBe/t8NpF1VpPFzRJa6rQ7CciRhqO4c5GFmiZcPxwGJO/Df7w
jLxVFWZRQaZRnpYW3UD8f+q+95EAeyLpDg0NZ2uaUbEPDqOa6eciv4ROBEh7MmuVFQnDaJIPop+9
BB/Ce6anmtgDmyciOCwYyDDyKHU+9LZiErwk7dbf4IiYNrXGCA63i3JbQHcOm4VfPV5H/CemIesl
u3R7b5w9T7QnFBIpmMyhzyNgoQw7wc6IKs+2axDu+IfZcdwmmF7YRYTs1BMNYnAw3FLNiKRVomGG
eKVVJwjZN2VMFIgOAHmux8KE4xRlD7G0xrMMaTYFRDZNHByB8EykI0705OacUbkKQSLjRKph+lZw
naieCotpSOGNP+asaLLl+fcXZ+gdzMZFelM9ixkykKW6nraxt40t557z46jZVN7BM9j0FGsRTQ86
SfXQR2I37rc6TZJUDUA7XGk00wlcloSkBSFhtvQ4kEJONjW6dssajI/rYLbHl25qtRMA9OHOt0kO
Tl1SrMGytJ4AfFG3hHaDUnIR462PK5YphWdpUEwOY8WPrn9lqRTrVBE1SqFdrdgdztJa+cV6YdUl
Sx9gy8Fynb3iLg4xVndtZ96GHB3KDUgB/iBRyvGTtfchk307wLHplRJYazeW6n2UShVTh/BsDRtu
n8QE2AxXy0VLot20aX/0yYWo5CE8rUvWXRtyBLHSXm/acDq9NswAfv5MfIwtA6pDaHvbDtZtfZDr
Uu08RmHyp+CxBZfFegak8BZNZJ8p0U1dV7NxFyxmkTUhAPDFmM+nTpr1cN1sbMcuvVZLuTkeoDLo
HgqRe3TLTrQu6eSiZr1utBj6vqkbqslxW9O7fdJ/BfvdAjayg/ukPxGEzRWHtfEl5yEadXIH2jxa
dqdIq5hODoyAFosrNvVA2pPnzpEnJZl+or2BviEQLvXC7NK3q5S9m/JxKUfqyaYhx5PF49+93OMF
SSHEpTJV91JnnAH/5XD3DJQpcNZJK2wFwvgbQ9fpMopZNR6yy2mxWGVSuGaJ00swJZexq4UPDgWe
U5nl1rNrubtriZk1n8kYjq+IenYzWoZCg9WcWFKZrizC1FB5CbDav/AGVw8yYn46HTDkGE9nozNk
m+sWKNIByyVFifNz1EEG8k8SanIgYZDIKiEUcA5l2jmKlED1oRx5tPepG1RCUC+IE5+em7HT1FDx
U2O7wuHwYaCNjlD0C+HiO/EHS1ynvqL2ZOFrd9iT1sgCCJWtJhdcm4UOyn4BNEkj+0tSdplmRQyw
jAYled0nYTJy4w/rBOoaG4H3W+Mpir2LHEXJxE/ZQ+YzwDn0kbbckYgi/mTjCkXOUGvTB6IiseY7
/vMhCdaHe0AvbBiETvkY1wSQNRZLG7jzMRREcF/P6VmRtFeEyCK3YGLp6Io+3FdSYqzpoGPZOA13
qzP3tjWKBRmb906tQjq4i2XcefWK0P3kUtYEqm968/Rx42BKYg2055oqGEXxIDLqml4I4F490WZr
W4ZJB25Q9k6yQTA3trl3r9j3IQ8wylgqDXNgPJZpFqz5omtAmlDwNIjg/04ZYzAkj+AEjLGCJlGp
eLpe11xJfiiz0IW8xJIoBpC2eeCTHi7qngs+tLzLHEGolE0pNYuib8nxPIQLf0O/UH7dSqUp15xN
7QQkZyH5nXZSGcWV9Jn8AjBQ1IoczWpdKqoK2fwhQ17LhJ0FAIEzxULA8yXkjQBmv5vQH0eigIvB
28j1k6N6cDhM1AqeU2iQCJJMjP8dSEdmm++lOF/LYpTmesrC6P2J/Rc2NyuhUoQox1hUlPIHQhhZ
EsVlS3p9V7KSPXi1770hLIe3BuXqGKvww8lOtfr5UROqsTWsya2QVXFldpS5JnkGGwPdZD6zz/A+
oX0TdZCz5J27askSxc0DNfxqNYEOXmP/3tz9dJbRu6bFGMGn4iD7BAWK2+RPEYd6QhaJhVqlF7VV
0Qb3FfPI+zGCgLt1UQyoThP7wuKALBPX0ZhnIyEjrb6o6atX/VwfKNOBfeEbxKabHHTZPpJZNsLr
aFUK9kNvdoIyi7wJivfIS71n5HN/3xjBHhc7aydIC413iov0w9j1mp+l0lGzBfyTC1Wg6S5pv5Rn
ZITERzaz2JRv3rr5UvSqjc+mors9ymFQnvhyZswBLww25T3y2hvfBw0MZ1RmTUJaAb1rqkJqxa+d
juDW2o/uWmmrRRlb/R2Qpo4BzP6fpNI1lX5jyd9iswV5cKJg5K2RlLwV7bPp78ImscyOALp3p96g
K/mFLmDTNOJixYYgt8zLeUvYl7dv2ybhub2xMKGq9uF/LmINlBrrsCHM0RqiepmG7TceKbdYEh0C
9ZtBH7gdAnJNo2sZ6sBt/h/3LmA9O3oAU9J3rpl9ghFA0wX8IqKICw+RS9TO/q+/YMKVda4ea7Na
NewqwcF9150JX4iVf2tuRaOKiio26GU3fJUiKlHP4ooIVxQSfuEUvXUW64NIN9q2G60mPFCpVOHk
UMwTJx7FIB0anc9GEERUDA10GhC/Vz1O/FVU0wAKWCQVP7/DKhUnhRb2msrpdcfvqAhYccH6RW9E
I0ciL/Rv4opDwN8iAGsGyv453l7nw0kIK1dh9vrYCZ4X0BbRpWR50csQ+WEHVDxnLqVjNLJKf7Wy
5e29GE4T+//78JMmjFtw9UANv7VS1dWz1gpZEYz4Aq1s7jnoKm9d4kmTzZKlAnjHH+PEDhiEH91I
N/OckhxcZ1k7bsmc9C3ZStYg7gbhhQFifCaI1YiQMbnWfnt7X79aI0gyYR6o5fvReHdW3b7sCU2w
vUFolBm6W+MzRvQtIblsLO9IijL+4J81YsLV8u0MmQvt+F3BPX96od8woq78NZJRdmWx6vs/rR+v
rwfCc346WHOmULrorbJvrIgdVcibdgxNjUw1z9yT99Y4R+efGMFDUsW8+VGlQA/33NlQtnlzuJIC
O1GLdKemWLCCbJzS+3GdqpR2ynnHC89cGE41tUvxv7fA2mUdXolQzwDOFcqDzAP/qBwwiAaLgHOp
jTw+ZXYe4ndsyeJ8mkmxhy8oXy8vMwHg4CPY1zziREovU1DZ07Oud4FHxy2KtoLyPYl14qrSJWrW
xwC74kWGa5dO6uc+VV55z/ZheiASN4WtYfc2KVFu9g1N74XwZPSHNVNMmcaHEV71Bv8BQfiKmAsu
+e+Z3N/8ZkwhvzaBWLSnxDOtM1EAk2jYQxjLZBJs0lz6mTxbsYCZlFal8xt++dWMeDEhGPKEEhCd
oOksNH615wHuF8mm6zCtq0Vwr2U+GnXayeKBw2Z5u7EFW27KSwbk/VX9gP5u1/v06P52Mxgn69wT
MJfSxHbeBrF/DHF/9w6OP9LXjdebIbZoSFXdz5FdZTVtJsvNY8RTGolRXEiH3+Jcq2y4yyqR13SJ
mbE7qPhzPwpWpTQvhyxT68Igug7N9sasGAyYC9LVgYmI8/Q0SsR5+F3P6fcxMKYSk/HIgo80nFGV
SxVpjJ8UEVGWzcnTuqEyv3ccwOSecAPiTbLWWA4NO/uSXx7Vnhs661yTz6BIvwrTElivU3CEP3tz
3/Xm5wb8TE8AWfgbRad0zkAPHK+C31bSdMUAvz8y7FkFzafUOo1e5uaBqXD/jArIxJhboNfAfHbp
eUidGVCoWoynl+ehNBT2sTimt/x8oclWEvrKtz3USxvR228R4cOIGf3Wb0ARmzcr+TD8sSmR60sq
VsWwK75XedG/fweCScmmgTTheIpGRlPsZP/UZk8TxataYPyC4hxtLatnzqZmpPT+rUaioUFRB7yE
xDuKDrpQh74i4dahbwvCGanEClZVnojiWMV09k8UTUDzsa/qaqZgDjqv7PY8YsFNBi2lK8ovlK56
ItWh7gzw+xpWgG2NEsLiBINd2u4hGXrWi/7qTpBRIf7IdNyCuZ+n5KkmjlLyEUwRMG6/wFKe8/7m
AaOLCe/zVzDRtOAtBU0KGDq/3s9ySuS8umpHS/P32bX9hn4AjMcY53HiCqdUn8CqZVbolrzYHlhn
ZFhTmWV3CQCeg/x1dZS4LTDKQldj8gBGaTabRiVLURAVtCBLpDSTmnc4w5EM1RRcM3YBMMgBc7gv
suDxjz6vS6SjIpezGOKP4sOjJF6sMUea3Ug4pdMM9QCVInqBnPKF685XxRSNbtU+GPpnozrH9+6h
IPsZlf5HJ2vmSnsrV1681ATFYHRKDafyxOYXODiDlI5n1Xpw7Ex1bdEkofDdB9w9gcyZ05Ak4ghq
G7b/lPfDV18LxwjTYsdFw38NVOnhaHBovETYEP2JUbS+g5nT9KJn7CrQK42f9GCHZpIQ26Xncwb5
2g1ieskk8BK8kA9OXBdRkMfWioXhzaiv3wDASeF2bZB5vq535XPg51nKg2ky6C1pkJZOU52IWVJi
Cqb7E3GhaW9wRBLQltYm1j/lhtB5mnwwYcdaUAQ6+E7BtI2jf0BPAQAcD0YerivA3aM7PYK3pJqa
dM21ZiLRCLTFt3YeO6medsbPt2SgQTzT6tYqUcXzmsxPUxcgCsNttr3l+uEh8GaXJJ5sgkFmryoR
aVVlHrhwwtSHwwa6qSm/8AihA3yeURgkJWb/8Jd4Cps/uVURqcFgIgbcB8F3eNFIFWEPqhQrPg4T
wWaG7VdsuQfeSS6MQO2XqLvTWS5pG75HZVaxXn/7Y4I6wSMno2OdbGLvTjdRZAh+d5EtDkhurLv2
E6cw10ErCGvNwklPsJUKtjLURjmkdA7VJqbjpGByU8e1GBhL4b5VGUm8SzFM1XviKsUxJEnLTy+m
Rx4Krg0ytGVu8G0VgJoLbudOu7+fK4KdEOwETpZFwfJHxAh5n5hUggpEObWVqZCJf3rsniQ5FF9C
SBJ/WVBHlDZnUy7s6r+62KEZcsk/PRbGcbzWE+q0WP5xbQsPc3lCN5MaETN0566uc6cfj9j4qeE5
5rkq6/V7AAl8TT9FkkMk2efcN+PGcGaxctXfiTlCylerJPxk+0o15HeSpeqCxUY+hTLiQh60/qLU
PSYbaUCzZC27No/pi7ANwD6tXN3A1XLfzzjHfVLfvIFy84/vwGJgXayTT+0DXn3ic+csra/kP346
NH07WWPgevdynM5UXWI4oJA2HUwGD2X2xaR5W/ENsyPqLAWqFQmfp7mbqOlkzxRtt/1BJfZzuVo7
X8U5WMR/37RDDVur1bQbFxQCQIx7/HuBgh3W6EydAJtevGP0zckX8j5ReLX1ejiQ4SP5SRmib6Vb
gpiRt0eRZl15s+9wqe/6bhRNBhAw7XPdGFYL24qXJ2kozZzqzxJIgOCQuQHFQJn3MK/FRagz4FWj
asime4Ro+hCh0Py9xwSjp5o9dxh/7cDk+tWjJuZGM1rNAvwWW/L7mNTb13Jss7rJv9uDIPCkWe0W
mD0/pQhgRRnaiBefCtP2VqhUS44ProTDPLek0NuU0hH5Qd7LsU2OlKnWLNvzxUO0XTOyNnfq/2qb
SYQXglcx43gKGd7TKHwfs1o+nuBFHryFyno8O8UUzcbg98qsKENU1XnMX1JP6NeezdtZpErF3Qzb
R2ZPLl97mEGir52X/n+sWiab5FAMRRH/437jDKWYAY8pHb051ot0JNoA/cdhjQV9mGAD+xl0qY7Y
l2wl5Ar1y2MYAB8CFbXiTDfHL2sVTNNWVNaiDs4glAARnhPHptSZgQsczRrttDy44GdkDVuv692n
FxFQh85WQHMJ/HBpC+8QQTXqo1bs1oTm0lUViL6ojZkSRVa/VplIXyCjOjtR9X76dtCDIq8CFpMN
a63dKELFZxHVhOFGx15TGZ/BrkX7eansi+VLv1PAniK1WlorKBBxSpgK/wKtRA6im5LaDB1h0oRO
YRnRhJf1Sls1fUb4y91/j0j4uKCH8ANRz7JQavJauFKgjYzQt0y4Zb8FPW1ldusy3Z+hLh6hAyzB
QhGpwgz9LHXCbH7/SQFAnf0DH9zBhJCVpe83+9txuay/U29VOFr+yuhnv36kbkllbMwCHsA9s7IL
xfCAUiMDlo0cgT+kdgunA4j0tjHXXOs+6MlxgZoa+ynaz1p8W8XNf22ocDH1hLlsjnNvWY+44om3
GF3lUM9JyjIrPG/V0fQcqIRb3BtDymcfOZMUSGydCI2+W3tC988PzKc/j1kMv1zcbstTsJYuaKXC
6lVODDd7s84KBsvqo0+VHu2skCL4SX2cFN3oBEuox2hoIqYF70/scEI+WAO2TqYr+vNyhZzhfNGF
0M7PTsC5rPc0CRTCRki0G9qhc1PiETSrZUqa82Phy1YbhAbOW17235jXcSWcwFZZQ7+Ct9h/Qd1W
/epC6kElmP1wnNktb/FBkrMk+fbToSwZw5wa0zVb05JuISDLSfJKbp99XEiRwQ3NrVyjzR1jtTLL
mCCp0FPnSRrdEGPo3hcpWl/4sIN+vvgqvkiQrIDw2MKHUBesFiZf4qZWUpa8yUsir0miwXHAjdb1
mYxpx3MCjIj+0dlTWktDaQRj/m0ZeS2B5UR6MgsRrtWXYqTKfua9f7f8V5EBKR8UbmXJ01sk9HaI
jwVF+0H8qsaUP3z3bWiEzTXEjeYCQ4ebKXc694oL5109Nzac77iPdciwChxhtF3XLiubr5ki8/Fv
Qx+pFyXCgYy6C+cTNgaAqmmB5kHi2TQz1TFI2xWEAzqsMEBNbCb+kOmIgzAsBtfzl3+RYNGA8kK4
rnDH92pssVSlnODK+BhSCZroc9MYwoH23XhBWaDN+XzyrXr9Pj6SViP9Pcqp1F1MqNJ9PLX95Ex7
tpJCRHaJOtx6xrWcwiQWScm5iAuQQuMV6nnn16QS1u/uoiA4cgUHkb1SwhncuJvo6Gnz44wTcvL1
StbFYqXnJilW8j7ZCUpFhcAiWhwyF2IO2PQHw5f4JNRBzM5F2SbNztk7BnNZjB5EFJMl6XmZvd9b
GjHYl+efoVMYpICFjdClNPfngv+P53eXzAM1M3CH3eihFBg6gsPe1F+5slLw/muaJrSz5O3q9aRv
PVDKqs4oLec7W7XGi4lxCZZO2mBNfsfTKn2orzdofFPB+G5uZc9CpDOSyhbEX1u4Ewr2+ShFKbt0
WCFozBs3sJL5lNhYv9h9Vj5vu1wF41yaZaKIPv2x+A9GfaM6tTa2V3pLv/wo8+GHrjlWfUt/FjCA
M/f/h+djnbYOOHIrKjQLy36FG8rJIgaLQWSh4qjGsl3800zLTDSlXF36RQ91l7rKce/8pHAJD1M4
TKph1gJNYGlpXsWt81FA84/nqUBT3Td5oc2YvM8KwfP88GhVl++UfjMak37ymiMxHzcEDTHpRDz1
MVUMwLvl7s7wzl88MvecuA4JRb7KmzaBlosGib+SWjl8FnGablnVE4bBmoT8LkrD9sct9jgzfnqO
1mGSM3HX4Jj1UtNUkqqJ9Qp4G3+J28iMB4lBwd1j12cNma7XkEzjOAYEQOXigicx0/pZR2ir543h
Qni+NOTyjYnV9Z/cmW2YusHojXRs9BOjXioBlyjRoi5xZVy/8cTdKQR22xuZ+ubC7zuDPtZl22QH
8AHUz9G+7J+5+w2Xy2bzuL1HdKsdzJk9woKWSPzihVgILP6JkARys6jhFu6/po7rZtXOaH+J2CKx
+Pu+Ck8gFgVOm2XgQaHFRmbQC5DtodffPXUOWx4YRrT8syWbT+R3QLUJm9su3fojMkHfsd4+/yqj
4zSOv2FFB2Njhavc0GIkPZMorRv0vpsJtDQXFLB83dZoqHUvwFaWSfI3ReToyXsG90mnDZyNDztK
CE4/5kJAsSl6acVOAe5TDn/na8feBZC2aSMDrds1xeLQFwAppFm2BqiKrvsd0/vDkyJopv5z5IXv
cI8+TrVONlfNPVlfImeoCefx9RHQyZfFyh/e4Y3Zeyn4ii8Chuz3ZwkSwfrhfGwRKw9D8EL+3eR2
avpIaKz6l9cjcdKMmUuse5OtAx9HW6nNaV7S5h0nBlQ00rwIIPSzxBuWPvad2DU7oLtJkIjBSZ/s
zjvXt5YEhU/SZGbw/OHbUTegBo6iMePetd1Xyxth2WnOmXZ7oQ1VcuG1Z9l3S3Lmb9Rvj+pr45wY
FKMoJAVtESIwP/Ja7JH1SfQ8DQ2iunr2nl1mNLA5sdJcDWdtNbk+ZEAGfBgBkVwvBGDn+xQ4sxIX
2m3LIQvqqiX7fart31BHg9i2NbHIg1hA/SZyDSqT+r6yFT3ahcPx1jGX/nxptjXr1PQ+WPx0A3Y8
1Knyy9AGZjorlAjnPB+T0RpFqgbtfGIpTAOX/IbpfojrffEEtBuJw5jRm/rMQBxP1eZzVl2BUJma
yKSoD4inCTdW5DsOb665tQR96tykqE6Z0TYSjLGTl5BXapZKWGHueYe/dJnf0dfwkWc+dhPwDwQW
2H1ifHZ3/d44XTdCWCTo9xKBxYdzwzcHPNMf7paed6q+5NhEtBApIz2YE2uh6pcQjoB77ug2cqty
D72tW/kAmU8sL3OsckUeuoekwQGDLCD8i8wGsm07i348Hg6ulf+aaevo9piiJtKn+O2s1Z4kyQfu
jdVa3hY4yVBkD5qkTCHklD12u4rTGPlSQJJVzN+WX9UwRIeaMylJ4GSU6ESfHp9BR99ifcg0YKsN
cAdBMmJdxMfkhrh0WxchZCw4MfBSyh+pwQ5/tqbrPS8cHwHZpuaF3yWIByEyvxigYn5dqjg/6I9h
gg5jjilXnPjmSdoc/kho8fvP9IuYDvZ3qUZoE6Oj/who6reCrs4DawavqUVarzmG0qXGE8evjDoJ
xzUNWakmKzHOilyhmeDoAsdiXY1z2+OfHDBBtRGo28oL1GfX4D6FF5Wpw9oiVbHH2nhQbClHYNj3
nfxJq6HeoNMQCEfDf9Jv3VH3KKpMxNOPhdMqY30cEhUhtUWRZ8XdIYvChajaLJXXdk9S5E2NpIjW
jCehOlShgNuDpoM+M+6dNeEuPI04FZ7N1AHXU3aWlPnmPZ/FLEqRLPpZkwPzEQfDeiLdvk3r2Sq3
OQfMwOyjaH+8GsGzXHW2AyMxLNmYeJKdU3Z4d0kyGsf4DkD4x6lt4uKncyT1gOgKzMnHelF0qakW
g6ooSGWgLRzu0nXw62XSGGIJ9X1BCISmXVhkktcQdYXD+RIr3hl91hpUais4zbvxEGIxaazWsxPs
FmLhs9tjs/xbqGfFXCpxv6GZBrZHAPGlXr3+Mm1oTgPT87u09AyaJQza/q0fr0x8+/4cEDdSKF+0
+7XdXpjx1gd+vFFlySNfcbSS0QZykZbeXlp6MjfZQMQkwneMqi+kAXYu7ceg2/67Su/u5CptsydZ
ypxefkEjSyAr4ogaX70FRpJs5c2W5X8WMT511L8nOX0l87lF4gV4JIvlvkWjBI9+zMqvIPIXetIq
crYIH4QnKckk3yVzW/0jN6gF7+b6JnfE3Laups2pIyfnHNycjZHFk8XcMLeRtE0OMps/HfxxnbG8
h/Fcn2RORacVpFS2I6mInJk1Mq2ePQUASyor/Jb3A+mrsuDmNf4kBVGlXVAXU0qJzJcDaVhOBfWe
Iv3xYO+MwJIZ470GGMbytGnqGnMAJ0GGkUfCAmayjvyWxK6YFTRIM1N+HNkLRDGohVp3ZXjBoJf+
MrTUDqi2V0Lb3IsipKBb8OcoA0OZjw0HTMn5k+09QPf8S20JbZf/Lfc1yLlYFtTtLZpNuV4ZZ1ox
6oET2BeYmmPr/TjkR7U2xLT8WpXS+BXNBixqn4kqY4Fjwl7YgzlLMtkdz80XSMn/OYgZKIkpg4wJ
uo83NE+tFWinloM7zHY3zMuon3ApdQuc+I/whtuOO+V4vo+s07yTvK0Jlbipc+o+udl3YvYShXBc
M0qUD8I2C2Mill2INUHJeZzPx6QnqHxow0SSotQNmKE+HfxipxBSBusCj8Y7+optFrFbI/G6Q/ff
G2UPCVwR0NRbiNuJiUoZYj6NWHinuxv7sJ7/rI6A2tL+cwzrr1MYHB/jsHUWjzf6DiusSdCk9VTd
38663AB8jR7MEkbV/L7ZIZVDTqoY7nYrynpSByhLGujrq0jHfqCxGh8+c1aawMwhhVnfrnJS4Ka2
aDj2di+Kcsei3Bhrim5QkjbArHQLXKWdR1fgd1yWZ0vSPZVEHPQ418cwnBcVrFkZsJ1fZgQXEStR
NGtqFvwtFZupL6beh4OANjcGii/yogS8EitxZFPNy3LWf24Nn1pGLWtUi7DWeaPAEkeycKizdckX
sMgBJT0ngRNK5QCMnM2O9B2GmJSNJJLCox5S2IElezk624rn2Ikz7IhSzaMks/C4/jGctre5FVte
buBVG2W1nTSgBfQtemiBgq5kvCEMAmfU/vtRBwzLlhcOzcADUjsDsUcxC46o42ZcQ6PKd6j7Ihfb
6mQuKZ2LVDbKyWdovflL1IZKv2cQtjJgFR/n/6zJ8PsnFCAa+iBkqMKzyAQJOXPs/KpEIyi3Gik0
+fhzUT/JgWaZIjEqxIKKRq0enyPMlaMB6k3ZhmkTbh0aqVwr6N4l1dan1cgdvZjUkUSXKIrqZNS1
x5iF80Acpkv4H2Ouc8zY7cx27manvinGTNvx8UqNbzzkBJZEfkDb+Q3r4YaV0wCPgkwLwmeiZ5LI
lE8NiyougIarekyAv7Pqq/steWV77AGrB8Qb86ZT5Rov4O1vkfULAoz3tYROZlxX86H5tiCgfLFF
nRF/E9R7hcil4adjA3vK7ex/Jjg/XfJHjT5+pB3IvSXb91UMMJ9THMIZsk1U5H2005Pu12qnFs/2
UqqXjAis+Gb6+jSlGSFSJK5mSDaZw9LwKqavY1pKUhpVymKAlL2+pJQ0NBwnPloLJYfOj4RUv5/b
il94XzOKsfa0LraibMo/OuoA6nQ1twbZkkb42CcdUGUxNUEN6ct+H78ge6pbM+T0N7B+Aznyc09/
njYz5ATq1g4lXlVViTn0n6GGNOMesO3PQ25llwV4+kqsMXTxxTNcAIlVTDuI+bngKutk/IvDcNCJ
twozYKtoBqOfC9aHCJr236HjEjARn+4rR/hdyncRK/Yp1Nfg3tNt9ROzXx79pxEHdOzZNwbQlB4C
vD/oQul9/HPdAuvwXo4YF97CBJY9Q0g6V/RFUByy/uN8oMwJVMCquXiSbPRaNErNFqV5NSh6AOqu
lW6g0E+8/Bw3oqISGdtMhwEY4B75wUShH7IjEmJa0o7t9Y6GKstYXLLn4XGVpfEIt0lf+FynDQV5
h45ZPbRh4Iq1h+lu3gNSoQwx8MikxZhA1iEW89ok1UwOMK6U6Wnw/w8Ld0lnovTTJDzn5l6wZdqY
OOpveWOZz18ZK0p/JbslSGukIyxuLmA++4JRvy2brRxzsKn+GrPxKyG+/Xk/ScRth9JbRXFX6aVJ
3YlnT7wmM+PhgO4yETGx8YW7yQoPWEbofbYtbC3DnneXkKmD8ZqEhOaeLkP7vdjkABmsWBpGr+ps
KVoRkb8QB6rh9ZtP6hIM4MBSE3KjKPcZT1NKl5SvLEmxAeJHo+bWqNvw/Ca7nXqpywjc0QS9pRnx
M7z6LD8N/RmU+OAnKt8y+hWw7Psr/jogzrdRif91fbbGA03+Qr02KII0IWlmzitRTvMOxhdCY04p
vYTQuXtt2myxbDBAtAJApsCaXDd94wAsdGp0muwGfF/mGGk3J1Vn04fDGYyYpYUhHwru5LuOq/aV
vy6XSzN+XsYuOjUQKXpax5F1CIX1SzqEUPZsICSljlRYxtek5bIhHOOeWDiZInqjIBKoI0ynt9zp
E/XmxHP5xgubgzrvzqa1zK8X7F3Yny6gmnJplTjT10HrKqpi0V+xi0lj2sggHUlVpNzxW0WxoaDf
Sqi+XOVppbc4MOwpgYvUbTKc5ou4maCrbafsjqdWt64CqAt6PbJlnW//4LKeogafCjRDOF+PYVWt
IaV7lzdL/+tJMbDepsJTT6pkfHjXT8xMSgAFA6X6XJPgE8Dfp9E/DDKJghgsC/tAL9ZEkdIz50EE
PkZzAVnE6Y+PorbamCrT/ZaAsefUYNhiASQqUw9l8khwEMuxHFRQAKC/drgtfILTLDZZQ2GKadVJ
oL681IfdvwWPY0pJJCpRxu8VHli0oMcAO9TKm3u0MlsyEWtd3mi+ZvdVhEunHN6cG4euVnmnfnh/
jZW0y7V2kfGHyctHuNOVk9kc0wOzbZLMFNqfP9QkIKNng0DuoO5pMoYA/ZpaoD2g/oAoNmGCAZtd
BuSMSPssUBDwl9SH5BwH09HIaZmwj7H/7iACk04TlAUXwAlBegJKNtyiAbU+ujJ1ac4Dd47Skh/U
S7DaHz7Z478zywQB5e9jOMUHgBUglSCh51+Q0LQzEP6zt5MIekgsfdiaRCWvd3N5aGOBFZS1QNdV
XwZTIOxtMb2pK6iaT0QCcdUriyKF78xiCsBEW3M/a7N0wzLUU2uT8ixsV8E5JeaU1rIQV5fl7hE3
1+02bUaD9BHJINqDmv8zLSYN1dEh14HnI6jwrfn5e3d6Li0q5W7oUvV1lqEVO0dXYQ/750qJTNDf
dSAn8FMQmTjTyCD9pe76YOhoHF1ay3/INZ8DglGLnU2SlPsR5+UdA0sSwzr9ZvV6lEdcNsFeismo
uiBb6Y6jOW/uyr5pZbmXgTW8VjAkSt1ArxbDGJGshZKmOc9IaDDlmDAqycU4EqJWvux/w4KCq6Zq
XeE2r4VxZfLWqPXjtuFh08x4k/UWKFaazgYmVj82292WthMtdvv+kpBxWae+7gnosOaRgiYeTBE4
Hr+eI2xg4x99TUlLxC26q/xtvZely1Xo6cJm7DtpjBQX+6vqbWA1KEC/He0X5Ct6tBH3LCdW3l/X
9K3xBluulTfK3RumZ9804K2CDxozWdBgDo3Q/POOtB8szH8AEXnz1lWKiqj3lYZdfnKVXkJFJ8M5
rGZKmzFoS5MF1yZ02U2aWBdNS179HcUpI/o02nBQH1MZFuNKt7fRwQGCp6RIQTT5U1sTF/kqM2ye
rRsnVubejaZlKacpgPFFpvkF0k6iGiuOTCCNzPMnq1GFhUDlqyAvvYQQ5wQNysVEDNjqZjxZgxyM
BIs4fkUaru+csW6YDaY91hnRvwpOuAFs+spI80f31wKvfbw93CyDjfc05A5FXRw5jmKilHiKOC/b
we2yl6Wkqz8rvdC+fIpAJnZL97e6lgRl2KqkIEbGd1isGekVOgFAuOA6En38eg6HpLw/Ec+3QvqG
2eKV6v0DE73vOsbiDqbYLct6vS7G+J4+xcN38Vx8Nzh3FAR5CX0+XcYb4T1Ef0rni2WhMN0pYmgL
y+OjPa6En/L7Aqz+jc4E/ssD4mzBiviF1FmQWblsgtE1uY9i7YgWpisz/7Fgz5XCxede2Buv27ZJ
jjayQZYMewmLfwiVeyZbnAZEwxeZAWEPT0ccjNGwsHYu2dhNG4Y579kAr7CR6inBPBhUwZKQcOzY
IoZoLKpD7UOUBOtlzOJJxOgMNO7nIFEgkK/Nm6m73ZSAjQ/ELnV0T17bAmn4+3qldnepiHIHP1YV
qcv8A+aBMGvtNb54KvElZV5dFVWgeY4pIGAg51tWCvw90rCIEFrVjqO1+vMa+JK6+rP/tJjjL6qF
JYmPH72HR/sHW0ADXwqzmLB/BW/Plex13mdliQwogl7K7D8s3ZuRGGaWysq3iUqpi5mdwgQVcztP
JUs8S5eDggsw1D0BcekHATbSN/inbiSN8xiGKHnjiP2p8a7tmVUcNwv/Gmd8sGgtlkd/KohzKNFX
/Evi9i9DJSI1xTF6WJ++bn/4FdhVLaKXJ9NG3l70K3DD8pilRCHU2h+mwn2rslkVl7HxJ/uVmyG9
BS/zj+/CK9a3xbPeVols8J9mHikAILhMNOrhzG8iYn+JRFSIZ7fSwNvSLSa1zVmH92lszgbHwG//
xgwW3AMGiGaoWUHJdVtdWb6Upucciz2v6IKrF9QRW7v8/IUSnKAqb89bbvthlKczGWcdpckJPcmI
JG9/lK13ZHLz/lIE0oRzPkgYAd6Na0jhSZSN/8EAh3qazFz0onOfcKH03hfri4Php7Yo/cnqFqCx
i3MB5YoO6tRtTD/vRnELed/yWma1bj5fGsIcq4mnanNdsjNpLw2JJzAxkrZMLZ4BcxrEYV4HYsUd
BloB7OMrhBXBWM6OlkGb+Q7IE5KC25n7fuuORT5NDg+2HSV7LO0KV6/ocO0DSX/hOkR9ElNG2Q1T
IOpIjRweTs0UxWjaeuM45yWkOzd+iYoRszT7FwIwCMwWpPByIxB3AifePjA/WsDfO18cMM/pmKBg
TN1jE2R6iJCN8GCdwQ8uzhWes8llyD4m2MICEC4ABUNh6p7sx2yRf/GkyNWjA9BF7ZecnXOcMssB
bEtI5+ORqLVzvVRZ2jhP7hds2H7E6QPEyUUufg2Dqvb2Kyrm2emfQW0Kkg6ELUCMcUa67FJDRwfR
eCZnF14GUtNy0eyP4kjuoz63X5ybi2osi0hFU3GJuD7vDv5moKGwIeR+GArBAKlwQ/uCYnGM4rRa
gcSXuJLvoXz58A78z8axDQkxBvqwVQ1HnQ5SR09UdmKIu1KQ2mCeplfyV48JOBu7BUGz2dyt5OR0
9+8ylKMiH2dAJiZKP6cdWQcYNyi53NwCJJnCmIlhsx1pjI5OWTY1c3Se1/9qmjinwllF+fLv2wT8
+mjTzr/pkBN+P4U/OJISzQ1piBN7E2ZMZihvCTAi0sImjGlbatVYWySFPT17KqZVLFSBHONKXeZj
FVZE7Sz3hX+mdpUeH3czc1w64y8zHYmzNVdiTvBb8OxjaYBWCp2bGCGNBAkBpxprpK8asIeu44zz
tTMwYbw0HIDlnllApjYpROrZubrrnf/sUM0eAmHirDmnI8CfLgk1qcxxBgeIpEaP7GOviDqBkwO3
99InrPozH68LI2Vh8S94RuBsYDavfMwSOlJ4jTIURWwQXjBY5H/jrIgAz7JD41TnKIGBbMEABLRp
9fbAyahfENc8jKrZsPMrjYr0UhjMsD/u3mEX7ED/zqB+hEmfzmm0+odhbA6uTn7wFNMO6/ueSan+
Qw70o6M+vKY3+21Goo2jc9zBiPftUUFXsiMx2SNiqQn34zMU3MeecXwmCEDoCbKxXc5jPLaW219d
8Zw1zEOtL+aWwXDV9W+3EeXimuD0aMpyajdPtDINQVOgj1ows7fCvgIponYXBUp3hEpD0JBuG1I8
Kt2Z1hB7pArHbjxXXI3Q07z0vo40ZN8uq4EAjyaWKxrWJR6yz7xF7R0PbYi5KPWYAV0bEl0axRwQ
PhNX2d5ZVqht6CFpA677XSccjbZrqAozkWtiVNQu1VG7XsIAiBNJAxEF/QHwuQhJvDS8wRqbG0Kw
21CHfx2zgHTz6Waqd1jLJGDeG2bHcDVlPv6UB8qpEP6s84mNhZlT18rRXCXTP8hAksCPsnETPP73
2tM3Pu+XoW3ubKmRxFRKI4wd2mnR+623nXZX806/rzEnGl7LMnGMc3fjEppF9+i9MjBPCLAU7ai8
kj94o4bdV8t4iCyOHkeBtz3kYDxJjXprb/TUMXZKVtcWf9HNKLDt+sVf9ZKXTKXJqpZjnd1ZqBWx
mexJ6APdyUYUVyjKzzQyU/pgSW5fiXtn2UTH7WOG0z5Xm1jTw0ishmnjRzgIirWOAQ4SSawRSzIl
+kGIn+GT0y01WMBc2z8L2MvsaqWayUDw0zU0l7vkls9EOSfOKaik9NCuw4DGReGRsk35LbPkB8KV
KMKrlt+efHskG62dptJxLkjp4tks4kvrDHfr7tRgJtmC1ktOvLYy9TDr7J9F7C4eVPB3o9aLSvjk
d4Qyz/6jwaocvZqLvRk/8rrZYgdeZQsaFYvrqf2n2Vs2IuD2h8aPLRpD+ldY63zH/sjqQ6lwQ0Xu
5Zkokmjw/INoLw77P0VK5of7Y2IDOF70tZRy+W5+YhZgrsrYhk3cE+IC7FIKES5f9axZtN2OPNNw
4ruslK7eC3UcaE6DmvmVoM+3n5KsGS8TchXMDz90Pq8z75N601ySNHbF3bAaxNals7kzAV9p8y9X
RD1sV2FVNp0r3koUcm6VOGUu8ptGOKRQezZaxfA943vzXdoOXmFEbr3wIgsGAIK31ytwE4nnyIdI
hwdYVjNQT22y1pvd7Gk9StTvAkScS2X38wof2zRDgzLO5Fx5chM0GBuowrFL6K2CSW0j0xnGfS18
6sRB0CFdd2STDIjIP7vBW2aG+VF0w6X1A5k1XxC9YHVrqjs8+Lmz5Nktm61hg0nyV7a9FDLxh78D
YUvE7ADFRpxnVS1gJvhU/xZ8bSfN/fODOvRdbJGqdgPNllfXCIO1gRxlTSKp127qvF0eFsWob+P0
4CjhBgtVS0m1dFIV0+/ysf7nyWwWWh9zxc/JLIxR8L9thvQuPu1ZdMIUbRJPQ3/PnvB61JcUNQ2e
yQtBmjeu5SDKD1lU0yOpSPjb7AXNGnxrFGik6TfuRZ+MIR/86Jw7gaVIfyrjM5gfktBsjB61b8fT
3gkM2/NUPSnc4fZb1FEZLXQu6vieQRyIkpHq8QEP3h3HsbZyYaoU3cK8I1PCo7a/hxRPREWgyyJI
sd1EJ1YlFIm+mlezXAGM77aSrZO/I954my1TFNO2BfgrtcO2r5+jJrKq011TQcIia53+FLhxMhCw
2W935k754Rra8A3l6+nQS5ZbTS5alSUNkJwSPxfZNxr3OWc2ILwDZ4kOK+RCtHV8xkQuSAi8mB91
gMrxb91OJitX2kj+xFbxKJOQrhLVekBt74WPLSGFw1YBDP5tNSbgBVCg9V5huTg88kJOq8K19CWZ
EXnniwCwbNMGNydYkO5iKSjNTL9qDLvSG88ZR55Oq9/szCyeeqIO0pvi+ZJN+mrqJSPDgqAtTeDr
7mdQeYG6W1ie5cSsoRZmPmhZEL24pMfcwGANhaXH1nFZ0YEtqu90/1CBpAJO9baFYsJCCoqHeKo8
K3ycnquOqpggTn4uQzZNMZg2Jv6KO7vALAa8r2ADdRqVVPO8rvyAcRkRDtTwCiwHfZUipmjhzrOn
mahDCJ9nNBeo1G/7iV+S95G84JtkWpWUtgaSbKPOHaoHGwXfwmVVYgigfSd/8IysbIps88C1XvI9
J2Oc7drPp12jZ9AdoKpBe/kR114Jf7QbIQMsPuFhXqw3ts+Y9Rr/MQf3omEuPAxI88Tr77SWKb8X
DskRJ8wt08Sf9dmVmptZhVsda3Sg1t+vyKpOWFRV3BM/FT80LQWPk8hs2kIlNvAPaXAAHcufXydm
WQT6o3Oinrqvsbktn7IRPYJse8YfjOMORi9p2v1t+IL0r/mRrSUHFDOW7eImOE3v2gopfCXjwR6Y
l9HWjOb3guzr/A8+sREeNyJYyPdUOlrggnfWETe7LQ0h2dfxBylWqJ9jP88FmbdodkvtbAXeBpRy
BUP7Uwub9tfrhRISjQXPml4AF6XGaDsQ0XhqV8YZZQBcmE47xGMGPE8xn558XpiA7DiS1Idpt6pF
+zpY2/kTjStNlHGEpuZabgQC2Om6Xdb0Aa1zlV5pldxQCjQ4vwsV2SmkWectg9LLcHA2jAw7QHyl
PWER5/gREt0XYTee0WjQTUy9Sv6qwUXrnz39Hn3pZjBvRR4ysGIOrd+UxCGonFG02K95pZw7lAOW
YpUv8Wp739EfuPuLvq0yH+usBwOEtTzwD0YyiTNpv+7Wx5Fhfz3fqVxwNF61pmA8cniylEIrC6OL
LNeVFif3zHX6cbsvNL/1EqDy1ZAWU9ekKNhZLAgjViykqozQqxYP1Uhgp/QgSRd/3Dp4kPdFTS0d
5cxpN5GQlyNKIossQjYIsxm54wsdLtTmuCeZbQVN6JAKRFaOY1oXtuB1ApumqvJ8IWM3ND+OVb2h
OdiTXNQsF/aFoLZVqye22vzC2rAQ0IEpnDP2dUNrzE4fumXoDwI3xXxkLzjakHj9lBKwWQ1vassO
e4ULLg1Hx4uU+oLd4qDM7dxwVMBAG5qSo5U6DJZKi6GDYCpyyVmZ89wa9TUQL2+AC0Xm2UMCdJS7
BL2UXF4siFeFMFAZ1UtxXVjba2roZFKxqN49IsOBmlc09b4L7N6mM7APMKsB688PcLoJuPutvf+T
+hUX535ZEDpSbZYtdoUpBnbB8Kfe2F5L/n9XIOq7WRQpT4I6NSEm9AvReU+ZVuKRRTz0v3DWSSLl
Mhc7eF9UgowRcntaM4AAaG0Jqtj96q1as1LTYStJSBZ8d2GHZ+rfeW0WRGZRMRzBjDWkjIJiDjd4
jrVUfUOkmDcK8iqWS5ucW+ArUraGsoGj8qj9Fs22Jb2prU1j78FIkW6xdikNjazizR4k5cULo0zY
aVrbuhO2ZDCp0BlDa+f4CLItJBNowMWfX3l/tGl4b+6n+tMO0d9gXgEESbaCbbCZkYIwkiiYzkpL
yA+sEJ6uK29HUOTI4bXlQWMrI8w0+ECnoX2dgaTdl7uSKQyySX4QomiNtfRayoX3DBlHk1YdzMo6
/kY2UooxZ+lGPGpmSOby9FIIUS5sm2uWKJadi5mdsHcH/AyZe1LMZ5mCG0bL4RbaGwV+g+EHgfWE
XFoblFN8ydg5XvJ4VPqsCnOLCBxdqycgB7AmlizAySbW+wopxCgIPwaj8tEGVVeeyxFaylh2B6nI
U9lfkqHv8PviSHAMi1cAAhjnmJ1SUtgEtym7DSydQIy1gZxCqibOUFL1WiMgg9OYH3qTG5PfQE9F
anI7cdQcLJFa/3YbuoMV81fZc/gTj194klgRKr6mVVhOwJ34a5xHfkiH1XzxfNE7oyDQiFhoGNmM
Wp+Cp2d5qKI7XO6qyF0D6zOQqlhwx7OlPuY5KOYyx8lFunusJQ/gRdMatvGhTnWuuFG2ijxXMkaD
JyXOkb/i3W5/EPXgn79X9pNJkvQety5G7QB6FSFbevEN7dDqLevA+4VcAsa8M0aAtCJAiNMLPgAU
bEgPQbv80V24CYCfq51ab8yEtaoePxqaIPUhF8RQMeFnLo+Z+5e6T8jUokqb8jdhqHm7zjl6fbt2
m+uNg8MrtMlkVYoo6daC5//BWG2yi4xgpiDRO+Duiqf8UiBckF9GZNMtd5uHFoMlM345GkUAke0w
YgOFnImNJ1A+kEtbXDFi+Uj1VjFVLGAy/3oLAV6koecJpN7ZjLTO56y9jf6aLaL9CCmX3Q09yHSc
NS3gRMLiU1BPFNHuTZcWTUCcZea7J7oC6MU0sGDZ3vhFDugcMwrrKVM0ADY9y+MRfaHqcFfS3hZY
7jX2M/s2QwtUPUcwtzMBAzIgU0y92eZ2/pJUAKKqk4yNb88I3GMZEN+CqQmfqT3ruj5Hk7J1kv8s
3CjKivMchymOSN/FlsdEtZVBpjIcc2oD7pIUBBiwEUHoX3wMFO1AwGo2kFADyvdUvcgzmuNhZm0l
NscaaSxHcjQRiws9Os0EyGXohwCfT2U9Y9I9uikIulKmaedr7gTO0+ISe/2v07u/TNaNaCWipyxz
upZXYl4C9o2LEdbpYwb5UWdwd0r+IyEGkN1y6gpXOKchXmBOPEM741ZjpdYwgFkUXNmQDsBH3X/F
FFGlySI9cBzzUvwVoBjePCrcb//tFR1vzD7inugJEmecSl7SKs9lhbEd4gZ0dR6yNdi5GqZtMCjf
ZBSy68MqbtLAww6+KXiceM2Vmyfv941qnFGGA7tADMO+VTehwP+m1RZk3NFApojEdUpNeutgLHGr
SfVDfjr/kxzEjTicLw7acgnxmQQiESnb9iE87LMay+G4SdJjbMLnxBjuU/4KQKpnl6wmfS6VwelS
QIcGmVbjVsR8pNOYT3vn16ddnImkHw2cN3VagQ0nsKfNNCAplss81f3IraYSvCnNTaKKdOYggSFE
v2gnLmDbyQBE7vdjn8i9x+FFqiQE13rawXTH54o0zXvp/zATuy58rTY3YyjsmRVMTmHrdRgoNClC
Kt7LHz8eEwPC8QhvEurgLE/ha6H4AKmc2vi+75pdZrkMEnKFpCuCBviYM84GNVzrRbht3MCN0F8g
eYTVq5ihpINuUi37E8c5Ss8BFGj+siicAwI/MOC0nuplJ29C53Z4h+hMUf77T7eEzE3D8kj9IuUp
U5vFHDgfwOQFB4kltgPGRwzZ0T/iLAcLSX34q/IzHacEJpYrPXfwCCfUA+etuRbEGpenXRdZFSTZ
OHMhaKFwWwG32CNMwFJhJeZnA9uteStmTZi/DxtLUmKsZbOiVjRbQIJH4D72o21I4B3hJoXVpGsr
TxDkLzPBX4jhq3Gn6OPSqlaqTlxhsGLaiqOlL1mseYAeBF7wjX1W5HlOMemUx/ZH6b1UyjEkX59V
0pXABI3THk9iLadlFVDLnvC//EQArCjNGhfhg5rYzn4o0R7nxeu2zuTggAEj9Xn3two//whTY9Xy
xCtxem7gP61klqNPQ+AWEThpjZdEYJaWmHpJvbX9JALgPitcbEckx/l4KDva9fAOaUZIlpzY9DEs
SKtTRnDUmCroI6eVZaT36+xCvvxgNU4IUJoa20gpSinKDzLdEBiGUdxMnCg3cPjHe03Q6KB2QLUV
iHUdY2PpoEAeoiQWEbeXsvxjEEvcCPMF4RiwYKG1viwoA+euH+zcYEYmxFz85g9nre4jZoC6NXuG
t7ypwh0f76QcIifA3KBXxrz/AjTaZ7DaydaFp75YZ620lNUxJufsYnmly5XbpVBKAduL2v0XOiO8
U5rtH22A39VcV2d1QDb9oN31OhZ9Ul3+mvwbKh1YWtNpcTPQtE44zk3liIyctmmlJmPYp+g3Fest
Mx93fppzmV+Dipha2NRJJTWydO29lG1Vhhj2saihCBrUeRIhej/yx2JM5WDlYPl8G0geV0vPgIF1
bIzBQfWJZg/l+IDvG4WGwBvCwYid4B7rsnub0DWSFgW1ETKolfHC7P1yPr+SMSRidj3E4aUE35N8
cmgxJe7HF+N3EpqtE7mCGQzhqJhckYu/eX8QJO5xXsdhrNFrRht/4g3oEgiFmpXEvShTrTtqY7Dk
Goa86Go+KiBPQ/W2IvwokeSSEdoGVNMOYz25Hdt+pOQ9KOBhZDWLDWZhkdu+yF7lJ0Mx0aSYDDTx
VUO7m/RJVsDMpNRkFHk2Ff3IK32x/19AhencG26pjWPJzMQHjvlllm90dsvm6NjNJw1YCdR24Dcf
bH1T7MKeqj4znvVOKUD8v1ZmjkFuL5vGnUoIzvUSCQZLh+B8HCeucAxDGJbZLaJ4c/OgibYqWt0i
64xpVTto3GYdIZKSZb4ZFQA5uy+c0PVattCXkE3Al69KNLvxSWpofkp6ZJR6U5c66euQaoom6Vfn
8Yuwqy+8Yc8S7Z3s9La7p/HZsMF/sXb49qU5uHqhxb1RPPCFIkaXRudkcABkauWERTf89+wh9EoY
ues5lg04Mn/8B2yqQszgSFt/HjeSUa4+kAdCxp5m53GM5Mlp98xuVgfv0z0zOqsFz9FIkH7liVXe
BpjQ4MRX2oCOCN+e6rLUlNAjuluOwP/ZY+4i0zQzkebAP3FUQzEES0Bp6KSR3JNF3KDKf7WjtDOS
2tmZx6h5R2xv4eFYzNqaTQY0OUbDNTHa5psL2USpFcjlYeH54V5OhnK+LMD83mMq3DmbG6cVlxhc
wwQ7fu2wolw4xLTbp8LHyulHMmYHorkUpt1Yq/4uemqI7oxNhLeD2Bohbjl/9+0yVpFOhNXSTXCf
3su6/LIJ+pNfNnL8QrQ6za3q8ZF08DsDO3XiCAnW2VK/SG3tUehe6tMat61DK85PyLOCrhVjXlQZ
Hxv44Up4FQhOdhqBG3wbqj1TUOD8zRRoF8bRYJttZnNj9izQdp24uvbTTjPYII/vDzWxUJwoE5uC
0NVFDD/h9zARJo7tRz0DS+olhgK2FV9tf3SR8Vws7YYJ7LbB1w8/6utQKAo9FSpnd4OwyE5n2MC8
yjpATMSqarFRlJfvzO8UHG/9siH3VLq4IM+3K398GB1mtsGOH5VRfCfw81ljoNsrdqojg+TsTBrA
ADjTw51S7Vsi0Gwc6BzTuHL4BI4dGJItr0DwW+HK12Uz0rE1o+hjcFQVa8Jq3WaOwywEq6XqJFkF
wDiIvw7EXlkGTVh6qj0Kemc0rsuuP324nBNkgxcqwOfO18C9c3KR+DTpFF4bEslk85j8Q+SsN/le
ga+1sp9lmI4ZzvjgH9qTgTk8PXunDuRK1Gp3NkatFLixMEIIcLwJe8536OsoW2CPalQGiU3jzr6/
Z5maAz34F1cuU2O+/trxqw6u+4Apyk/9r4HM2fAVM5hLKlCViA+wQr7dCLesp90zvTnD6OU6kIYa
SLbxDiSS5WtrliMmLbwL5fmu92eMnnAk3SkE8jXajVYarDYj4utb8AOT+HxZPwMD8turJoIZFiQI
F51UGoVa1TmfI7cLTa11nKnHFa/rNJhUsdsrbv0dNV1ZPtmRLJcjH4p7rzFNwpGBKEdS4NKIwNKy
11T6O5QNGSz0lvR7pbqtNzFTJyqStBR936YGh8bgsxO3Wyqc/tXQNaX6ijrmSCHB7wFbURm1+l7x
yd9jkQoubYVOxkU1u3Q1WZKEu3EmPJq9NB1Z5RnWyaJzls9ekd9Z8+BV6UDrBMS63G9XsZPmnYim
/iXGIb1oCBYHwvBBYbwaBME9H//MShq9OYMSOltzHR54f1WDl/D2SztscMKsv2FJyxFB1NYWHuMM
DMvNVNs5WlDOS0q+V1YvQyEJM7Z9Dts+3QGMNx+JJuuPtNl03kwk48VVi3PxrHGLAZUGt7umVneY
X8uELpWWR8VeNDRG/4qh0FWiUrPt1oJKWLcdzj1ZCJu8KWeUK6BkZ/Y48HE28h4mo7NP2h4ncuSa
o1BVudlLQJx469vQAUQxcnOs3ql3PCVH6wa7Ctb9+35JFjQwKfPYMaa/Qfg8Lc6WYoojCJ+FlgsH
Yhx3qv+lvbS8kRDV3Ku0XD8YhzdcLdBV/TovS4mr2mRS2EXYH1+uByDZ67PGSmbUNmOceEeINQaH
nJ4xpwTXCKl7h7B4EEiRX3pWPdL41d1WfxztvX+C4cPuflv89ldvjkyYM9qPN+9JEiKmIo8GHOBl
K8ak50UWBIRfW2bFnLGRLosJLVdcEgB6Q8KWwKKZ3lSBhvlBIhbspcBBiQqmJPRkZypVVswTcXVX
p4IjkE0Nk0JLEc0D1QiX2IH9S5EHTJwxiINfbC8YT9zqnR7WUsZPo92rQ71YIeeLHOL/0cxKgIya
JJvQ0QKneqKWm/NYVBrlf6pA0+UqbwB6o9Yo5waO+mxz+u09HIuAAEPUwPuDLO7PZ2PxgLuBMqds
3c2EsU7OImqgeZV71m6245tsTdsZsbKwGIy3LGttnZf/qsxRb6Hzu0/bPr0IzIAU8BmXGK2AZvzV
TmeMlcuec9Nm1p0lG4mhLBvFjVtHRTy9KOeu9nVXtwvStxdRVCFgxLPEIajN6tDQnhWQnOzBt00t
n/PTjS2kcJA9AdyHab16zUYj07wWX8TUICJ+n9aaZ0bzN7+F5uECPwkB1nL7XfX1grLiQKi9S5qB
uItEd51wSf5RCBbHL3YIGRt8LjQrelyv4zfvz2tZX7TeS8lTYf4Run2bhFMKPkY/QMryBQEoe/c/
tGcxca5wib/buRfK2X3eaOOX0BDEIpLusZggCTYzhWBGNJBh/9XXIv9qPTc9rlMEZxd0modGRCG7
FCjmyxuSSTK33Vc2KQh5Cl0p9JJzSqpRNRlHQfA82ZUcFssQg4Vjh84L3X/kv0C74yqi2HAn4FGK
M4UDctukwJZz1QS7oKCFjdvcgCxQbfr01TwCEQIMW8+slfEY1+IWjbMozTSs5240xcL5vSH6asQP
6IDGj8fjCzsC9BPO/ezMbinkJdURTifS6rvRUi1JSOpKUC5Q2x1nQX6Rb79XaPr8xxQTdLquLtWG
IdA8eET2r4+7Lgy1BcUz2pIpKnau62etNo/3Z5n7UNXbwQkxCYpY90RHreF2P28un0HcDIeON2hE
lbHUYPb0BUxsdRtp58xcBIhfR1xQ6f1q9a0aLAuxf7tOrwVkli357DBUs71KvX0Bb+KjxO3ql9hx
lJFXJJo3etFod9uzb7SMKepXUbwepjCU49ioyVxugvA8mId6oxlHLgnckOCF9lHs7QZf1N/8omKK
3D5fBTkpuY59hpKcYKnCIuUWcWV0JQ/57KKe+FNLKQzSuFwAsDdtFaDIH0HfHvFd0xQfIWUltPPq
M0Wk7kiWUEXrQrTGBpqBMoFlSGEJRBdtow0KSipkEPK4CrJ4FYngOJ6bCIsL0+kCfg1bjbf1Bn2x
9bOVK6e0guIOVeJ8bOpWij8a3NU/04Xum1u76oCQDLgR+41LD440OZejNHgjN/CTRabz1ExasrBm
ASCWYHiyQ4/lHnaXz44PaRpKgwuvFaFsnHzY4ENfDiYomFqlTQMrLQ6hckrjnezCMZmsSo3xSjzG
jsZkqG9Jowi/qv0WyKgm+15e4rDi1BtiHIufPWdMZQ+4kFQJIX3FoKBwbQ7bD0sjATdUhoCk8JFn
fgNBBDp1wz403t8239SM8jEwJYEeMeX8XgRUH381JUKFvw0LR4ag0fZ385BU/qzVAWcDSbLzvNyW
bwVGFT1oRfvuk7MAXRv7C3Uap0/1ySBzYf1Jh6A8USP13sZqxTqJ+L6WgH+YJ3jk6DeHuFO2kwmB
pG0vS+PGINWr8ZEbCNUJkGZqvDOqDE9OP88vSwoThGb/+p/38IGhTAfc8tkoQBotHAQQEn0xTK8o
a/zl9MrWzZdSxrC41vzx8PVMo0D/jiyFGbvk5gejuyWT19i0jt+nY1CNbRcATCyAfrQg/38qG4Xy
hwikxDQ0k5HQEu9vfe1Jz4sWpMBB+r5bqJ1/JJJLp9rHzq7m/LuthETbjN1rkOrB2X2yPaGnkKBJ
VS+rGfcnb31lnjIRgJ/aXd7z1S9rA89zMXBQQXQXrX064aCOWyKS6L6onc+SJ2ggP8roYSZ6881R
PV3sSpI5Nj3QwgmASilLWitPAxMq0z5Y3MDQnXYg0jaPOfnZdShok1qkB6OiK+ch3n/LoYDDpTc9
rmZ+AmAr8fhg9zmOy+ftGk2QVHEs4zTtREAYyuAP4xm+ukI9Z7lkkbvEke3pk4ZXCYyDydSUzVub
r2PnRnjuMguCR7kcmkh+6QIonhSkY4bQxZe0A6lgzgztE93k5mrJc9dNYyLastzYkwz4WvgnRl2W
lg92IwPG+7IoFRoXAV5dh3VdrIvMqmlM9PUS4ODa/QdqSJ3uRFsSY1AHe5j1mklRTPWeYpB59Nog
1ZFQK8QZpaDbPZAD0Mzk9yb7tYwNMysPiWm/eCBfMRlzwQp15AB/aJ2yADX4MCzZHoqJJ2B0GSPU
4jDnpgdTdmODipAhYEygLnt6/RX6FY3jVRMhFwGMnqZuXDREablIMRvNdA3oWcAxou/lUmP1R5WC
Z7ub+Bmq7r836tKciBCXXddMgtx8j+lOkpbLiyvTtjIZ6bWE2p95Vcv00fOOyOsbJ9Bd8bl28Ru6
3SO++3XzCKZaPK4r17Ri67GKqCTC35gWLOameoo75pedzvjeFLMiM0U37cuzETZyXONMK2yF3htv
dYoTOiBh12BvF00e90krZ7wUD8AYr+OLBhmTWM6MSqZVY3GZQcsVwart7rDuqhA/TTw9wPFdwWCo
7uMVAO1itCUHSRM/vublyrESJ2Kq1i7ZXZrQvfPy8QFXtBhSsR7p5UFSxiTFXWmYgeCDCw4mWu9R
TKxSweTNBMgHTg25+TgURl/LAdM0TKE9utl1tnrvkne3iS+g6NBEM+Nkql9jB6+BHoFcATmaIneZ
/dJr+OhfzvuGx92/OiP2L9q1lGOwFlVxRRiZr281bdyJRssZJHDNkKPfG8A58fYiC5menIvMaBZG
sUxxbC+fVxt1Yyy8PCpHVeTttT4oL7en768RpBKDCtzoxFHHLFmkSVbRP1RAJquTivMPZyT6Jigy
1+H6neCD+uHvfMn617Fle6AHmc9vUGB0kCJkl5Z7MJc8hcfiHQ1O1i3pOvctuNwR6r0w7BBWE07N
/TAVo/kt/O3ZNSE4ESoCqJK4t5dWSyKuwyfHMGgwnKieSAKEvLdEQZzLh4tjtPultZIX2KMJqbUI
h8EZ3wF5mWwniUkOJhFP1RK+Rku/Els0SV0nIWjU+xoP5HaQ7RP7gtOKsxYQ10yZVfW9qHdfniGW
SCpT9/ym97/IKf2cbWs61WDMcuFlq72WOJM3PJjuPITZmxhlplscr9Qe7AJMvYlqKcYRSqPzHJax
9o31w847zrwytCN3T4KH0HIdpFRZkj+tek78R6NN/+Y76dBco8B0se63VVHh+pslwOIxZJuXXRd3
9EBpHsS/p4817xanhVRK2ApUE4XOKs6aYNxH9i9VdQDNoPwRYUjJBTTWtVRIFCYandrgJf6/N2c+
LTNk3F3bHXh2bIVt3r0fW6/OgCX7k9pFuntYTbF8A59MZcranJPQxyjV8JCSqSsnHGWNZE/fPE+r
FJ3b7kZ3m20M6WdYcPFHiTN/HmX62EmLh3zB4ipoisf8Wk6EVZrnr81FZ6khTfQluTvQjxQQ3djF
W7JyEkRhWrZIU1eInXU6+86Oe/UzGGX6CMvEc4Kxp7upEqsy6ZmKEaUdFcS9G3cjL1i0nFYv8kOx
juQBeNMc7vGYVNDcuacpaV/qY6YkuEVKsZV2RqvSK1+p29XmklW82pZuwqLexWLvJ0k2+VBv0Kjv
GSzNpWkyTpTj7NROKvuCLPqI7nm/bTrPdCUcBAhIZb6/8icf8EPohCcOtw2G9NoAuxzF/eDktyi7
3bmD0Dgr7pHsfdYx7oGYApltng21iUuobeUZ5TD2sbRSFI50yjzEyhyXo+VpBQC22yngg+JY4xbf
a5FXWb3UthgUFO3Icaknea1764aLmOm6iIewASbVSjhreHcOTiunZXevDt5wv3EEndAsXede2NOa
q97kdb7NYQ2uTSdAr/0Z/h75dxmxGrPjKXrC+0fY6WHpGoQRYq6TtEPUt8L9vs93BBwNk/Ml/Tp/
EkYwD777bJMRylmPB2/G6BRZLsJk03GIQ42m0MaPGoL2TJ2ZaxOoUTKHrxrpGjKrTp3V/k3aYJyW
4JlvmnqiqaKDOj+S4C1aoL2ge3y/vfqq6vm5jbDgKvV1UmlypqxmB8zAuBJHCg0P2uXWtotXAfsk
uxN+YSx52lFWu/eKJr6ssDXOOQogVYViPlmHM7N4vNe1mDpGoTAYtanSzSlR/UEvJyqIx7cIFAXK
oTfrFrowjJG2paAjPaJ4hdfiaXu7+valZkNqDMxK9m/55FMrpkcMm2xVnbFUtgXUUkoV4Q/RhvM+
5odX4nAPDEx53WJBggpCz4hH75F31dZMbT5KNdbRGeciQXnLmQLXpdfCnHvZKjGcqOSodgSNgxka
MMLlTkXJMJzr8RXi4OpNVpa7JCPGXSznWH7CEmywWOTkPK4SewzBEwBXLX8UdirYVg/LiU2EAYSt
xYmIm/tsH/rkyIcS64akaOqmdJ4ZgVtsTqYAHhg6aTyGUK/QZ5Ol5ZGcyj/k/W2OXUIV6QwHJ36r
pmTBVEVJLuaeliXfKpXtCQz22Yb4eSbTnM8b/K6xZyXz29wiGW27JE2ZSAZBFkbxbQ/vBwoTbFUj
ZykvuphpGAtcR+yYNLYVhdDqlNYQmuCxikYecofnX45vsGn6/FWrbdm2Yi/jcxmlNTtqkPoXE5at
BlcqTHXe7YggaCV3beQDudmE6amD3WSZL+ENJRUCZSzBx6nU0leOeMWiG6hjP88W9soCfaOFaXL/
KfiOiXMPKQHUgoP8dLzXJcsca0ygz/tC/XpRj61/ms/oiKwLB3P7HhdhfNjjZTqPE68ML7SGP8g9
SbaK3o4ayqyfqise6yBa62DyIC4sua2Lae9Q5LQPMuvbIDA7P5zGPE4+w0TYgmAlSo/Zl9Yv7LkZ
IPBCdCnyIgO2uXgkyzyQcZ7AQVEIsY9w8NXB/Sh/KCauuxdsZkeVlIzpTmef2wCTdY2x0UsHMvoA
QLPBt+i4P8orWOSU3iEMpHc/xZEOIsmIw/gk6jakE/0zv/jJdrnXLPEhXuz3lIfiQFdg3Z6a1Km/
oz1WVNYJ9wf1wI1SPJ2IVt2VHchmee0Q6S7wVJsA+/7rFpeT4yjFeqDEZke93oIG+pyN65362MtZ
rIc50L5mnszbXqg0cHpHdvqO+PMGBvTcqkJfgm7KL9/TwYzNZDWJeZfb8spTA4PFhR3eaaUCONuA
h29rG7gxSoStZgWflmlaWWaYbzQqIH2p81+2HNs1WnWBBwDvVuSDQ5wMjtIbswCO2aeyjLG8aVpA
qiM/YYyfD5FqFap5db/Mx9zqIQpczg9UaBYOsJB2TH5UXBJyVQlmLX4EtD/IgHn5cMISpa+HBCbm
2FEfOkVeRzRInpj4AQaVpa1PhDu+2wLA5gqmMyE8x4LsU1l2x/AXLTkiiTZ4ttcQgqOPv0Rx38gB
NMcdqSr5YW/zdPAp6FWII+hjF0TtXxm4ERgipLcZ1ggFamAmvYkBlti96Uxl3cEGDVlOK9PxbYgJ
4mPBTzJ2XqoRvXood33e6HaL04KVK5NkDHDEWJqMnGCp6E/DER9TIRAjNXdB+MYokQ6sBBC1exE+
ZIG159cjqbCaWqCVpfdZDqk4/coQ2x4jc1j5gS6w53aZ725VLjPVAh0tee+mNtCneEd5CC6GeRn7
RGqdFPQUkD+qmiLbY3GDixYjnn9K767ZPdwEPKWld06qLHbaWVnL1vaa4IDJr0il17lElUkGsiQT
M0YzZUrN7qinGEti5LD+J/QsBrrsCuQ2rYWzL56DQEEQr+ybh54QgPmPVm/mDpo5xbcXmS1+8p4o
zor3ep/BYKxqBoyYCKkommNKtnPqedxfAsrqqz81ZYnkWGRJ5M/cLsDWdMKj3/t3j8sY5g7BvMsy
xd9TDX517N1zkY/uR5cQ07Qegxn7VZkGgUeJQROF974mS5ONO9lviNRda3t8aM+d5vFOtQazjJfU
ekgGKdbZEcxVpCEAw0VEIkfP+feLinKYDHY5lCJuMfsmi/YKkzT0xlgSO3wFLsgqic59+WPKZl2I
3jgMtbSghMHziU+DzSZv53eG7fUzpzDuQ7fJ/+HvgFy40OWaXhEJvy2nOC1G9kpyB0V4wb8fMYs+
TwlHXEuWp1mxbTnn2SmPPhYDvjYV5PnciYqfrbRV0W87+6lJluboAEJyBX7mFV4xC6dESttoz0AB
P3+ABk9uRuVD/9iu3x+56r9nmj+6P16sr7Q1xdUGfW0XT57VOuH0q0vjvM9rk2gIL69kdHaUxSr6
nJ5BENtm4bQBibiE/kQ3SdZ+u+Cn+jwUcaDCLEzI7cqN+hmHi7/TiqYi8FzPSRH7eS4G3tbowHLJ
M4WpaGIgvo2zBY1Q0VTJmdp9kuJvwsi2bSKen2qkGhTKFLTJT5HWrcnrBwOGcr12niEkjUNP5wT3
zPrLGJZU7dNTBU12KSZDLgWXd8cRDTzWmPYLZtALjkR6hDLw/6/7eQtYYHqU8iJ/7/A+oZuHdPyo
WSRxFU03TByy/1j5I76J50fomSdI/5/ZdP4p6FWTaVzn7tGtyTNM2VPv6p1jo6ozzQrCQ+ubJdjM
vwSOpf07pDl6Y1Q+j5fJK2T/oAAJK3Nbesi4cX8JqOp3Lj582KxjoJyYKmJbPXAbl5umPA7AWtas
npXp4q1YqN8XXVBi0xLpM5NO0vs9QEzgFGT16Nzdvxd+GqwsyXDjcz9MU9ixuQS4gH30OAm5+xD1
CXkEsWnvHfHq43H8hAeNNv+QM7N9sHyyzahV/KzqI4BIcXv/z8RoBQkdb0hlgT20xaCGLOkRWLrR
AlmRGaMlPtZJJeQXbWHv4cVvWucw8o/3SPwf0KVus9QiE1JAyiq1GVjwE4vaASweajwczvprb3rM
usPQFuu4XNGPFMKEX21LUkZ62nbaF0G+kmWO+5W1RcWYCFP9IVtDDgcC3cgyrDZFs7t1HYZzTa0F
G1Z/B7yJF3RHwPLYKlgBJAYZxqW582ezrr7SGCX3KFTvQCoTE5q4v6M7zXvRWVSC8ZdsXZ7kWfXP
ARy5kJKxQhdO1k3GG5OmHPS4wNj3sb/x0a0k4NosN3lY83sr/Js7ajLjlmeXZESMFs+W9KJvscvr
Ft2e7YhFJmV38CDZvhRd1tuj8/5GjLEFl03OiPJ1XciXFjb29ODQtuawB2y4j6QIflRxrotGNSOY
lKIoocYySrEZhQ5GGyvBcEIf9y7mbXALCw3w2botdg7lwKffAV1lkh08GSsf+DCuf1g57XCUFE7b
k4H/XfdkkFu3REw9ZDIomNSUwuPl46C4lIdMWs61PHhAy9ACC+skM2gMlFLAnOqfq/oVm/7bEJQl
4UxXxaTrZKikvHqdpLNGaA9V7+Ph44YQfWUNj3mVinqLrzmqb0mkeFrnq8JiuIvGnpdhunRI+f9j
YJCKf91wEFtep3BiCAKDkQAcuTdeKQcAC9DKc+NvA9fBhAIFiTzP+KgKSfucV4QYdFvhkTXY4ieD
BTFFcy0TBbsVUOuXs4bsdygf+ko+E851heoqA6254CFBzJdWGGWhjhZLAUVaH+ysION6CPmUO+1w
8oJQjKicWOjwdkzXXr7VCeqltto4DUiRw5IGh1rlcn3V0tsvjv3WJtE03uoStuUZzilCBLTx6PFm
4hrvhG2RF8cLQ2E3jCRK1/BIbFsX/H10NqB0EX/5lqYzv5eAQrJO/sAIH3TpEhT6JLjb+sANDYtg
gzdvlOqlHGDZ+DO+VqU1R29snF/0eLYvVFnwoG4124KLnouNYFAQZAB/1BVpamLyZ9r5Zbbhf7Zm
trclS2n6hS8VGLJKCEshNxqHA7K6sb/w8wTQbEVI/b7YJ2Ay1LLJAaAEvpakbCSZrYXnbxFhcVYn
BxacI5PINpS/WB8FyWuPxQqT/oHKkyezJfcdJi6LcgHQV1WWQqvJoKOtLoWHKQ/9/lM5ZumTNDim
eTStjYlqlfS+U7arZcoumqmGwFZVXWDYEwxB9Xw5xN/EladlQ0ib5v9b+dhZXfsCYUKymOvfwdfb
yqQGY5MGlU0TTRedq1F2A9uO997C8HzaNKBFaL7A2y9z50feCnYsVkw8KxAXIFh6UJhN+erX+KnW
XLBsdHJJDRco3AfwluhlQgmOxPW1xdXDgjniMPMIlKeiAGGQa9DtrEjZh2NAkhCRQWY/wjyJZqrS
E2UuPFSqYGcUhDw4u81KCr03jqpwTH8abyGxiAuLl6USZj8vlTZJN3fWtmKfnN8UY/vYmfU9fEHN
q15Snv1Ao4HwfBwTDM0pKNjzBC1hVe7WLrkd4V2/Yi1iHh0itAbzR0i+PATf/zcDEPuJv7IC0mOI
ZHqJ9NFMVN5+RsbpK5IzVM3IIDmrFIfFwDCHXvoibVjaaTjs7Q/RjHj1Juutlh0QK4Zm6y7kEGwY
20UJgL23cOlkOMKmxh6xhVbKakKPM+HRHN3tcmPTis+0AoAfLfObG+uDJtFy54jiK0gOUpzC6GCw
A16D5ze6YPJFQxAUW+AK1+oJWXTDfekR7Ea8deLpxyPA2ErqqurQeTQog7YLacYLo8bXxHRwoM8/
tn6ofFkuSHiuAb76sWIelVK8Z4+oGloJTCyApfNauB6RrpnX3CSgxXp/akwhESy0kkdtJKgMtHFm
MODuc3htJpyac9+0AVqryMV3qG7TLAb2oeNGudVb2295WigCxiJ0IxSmIY4DjHgD3bherRjUhxGG
cB1DaafrQQJhiwJSilffcdlzGOgtpX5vR01RnWoqR9jERySdmLfgAO0SbQ3OnRIylTwVHrBX0AZt
ydAoHTuP0uJA3tui9AcqZ39N38z4qcL+4w6d7taAU8kxtxw0+XU4hegCW1vGq/InYgYhzGo1eikd
4qGqd5kS06Y+p1MJIC390lQpE/L5mB2YDyGKoqKbrLVdoMHWUOdZHs8ZVXyR0+vrwwQ2AulUdmYk
eWZQh+LFNavU4X1NFSb+tZVwSLzVjF3UL0+b5PtIpENGw3j/V3DnVWFYxZGglzIrw0po6V/tnuw1
NeiIOVIHntONP/HHj/7U+8ZE7G1Z0CiTp15IfRHAP0n7dnfWo5SiJnI5dBmDl3u1sHIpQQOQX3JF
kNZiHPSHDiQR2J6hVd33LEptDZfC6xMopSX+mMSo+xa4+psnQkJLsZrVDxckP4YOACWtcqX3tYxF
bo3bPk0MDk+MPZrB0oHiVdFxLr3Ny0YUmwm3xA1yDHjJn5Ov3+0rkeDsreyUMT/nfwShu8pRhJHC
ee3OPX28+VI+C+5HzSCwx1EW02yvd9o2wKRFBXaYfDd0CN143gZ3MVnFd2T5tvjsQWYT3m17gwei
z70PMmvdtgg+NE0w8QRl03FDN52gF0P0uSdfZGWUmOJvpi7cQGSiN8sq9f5SycxQx0igY1L78hpy
mRlbJNTKHFFJOPhMwWDXdRFEbo+JLuue6F+52brjo2kbwJam91zdBnJdIb/4pW/b8sXv7s636v5D
zNwAvv1xMZqExzuCzsTFMvi/xuSfnSiP1aCDptb8kGvVp+vNyhixmW5jpg57vWj5FqNo3Vb2Bhrz
WIqLJJvmGaUltUEgdrB5ZWLZquiV2LerVI8iB6qpWuevls7Nylh3lRcz0zh9u+9an0rQT5E1Xxve
mXS4jWdLYqPqZLe8C0WFaFQfnqD5DgiH4Uka/NGJfT2NYCXv6B92wzZdHcDqA8bSxCRq2HCKr4DU
DcVL8bUrCj+DD4OmEgFxE6kJAuDZV7OJbjDoa+fQ2EOugEPWXh6o+97HsSci3ZN+MURZEKZxJwo4
5c8FTHn7CQgHzcZyfZHx/LU8EbH16GzOcWWniGUx23sPiU7wkhHikoaadBwmZ0B5bKnOPHavxtjV
QXACo0DIUB8UeOpk349jVA7ztSbdciY63Z8dm5MHB5DCjSh+W6Ka/N4GH6dLYdd1BboSymc0/aZk
yfDnchUvAHlTnUsqf4olNffdxDCoZ83jbOkBBGnb/dk/T2BQ8tkaCv5sUF6ZFT6X41pTATvxyBDl
6rovWd9rdCpLe6+U4VnQsLP2vPzD+EPwCaZ/xW1RI9F7RyqF3jJ+Ifm7ak9UU7AKg3EREALtIcEy
Lbpb5tGFbd6mzusLvIIA20GCjFFylrSFaTcsxV17Tom688HFA/USesiugTKb/swFob2tk41oMqba
Gh0eJTuz0dO9eQ8bmkoi2zO9xuGjCcV0YJpDGBYcBkD09XdJjVgEyatvCsMoDmYZOPW7WvVCUHjk
GNu8OfCSZLwgVWMwm9c7lucHbeMteIIpMon69RdVu2r/YGrdo3L1Ruo1KAELqrAQi6PLRxn0TaEs
rHez/tXfdaF7iBex3l87SUbQh9kSxq3KvlPCTk3V68Q2LlqAAsr8l3oFwG93UoM6NoPxMxAKg2we
DySQfwTnjT1/heew06sJvOwPcA8gd+YXqucDpwXuYbwMZDK2DFdhobjLCrAREMNnP830p6jFn3G4
6miuNlmKtvR4iBNXnRQkPUpWh5T2mRHqxuaF+oBBoCJZe4LNlzFjPCA+H5RyF+3jq/xN2cH3nA9T
jY+iJ4JRq9H0V13xdvuBkIQmaYYTVCGzL9vUhbMQov/hEMMpD8ldufdzA5/62UtfWXG6/g0S7aQ8
K3IP1tMkDzGbEMvC1VHEnmDFx0GpaOIVjJ7brpUO7+Qzi3Rrkqho2y6brJyOxP4sDr/zY2GEzduu
kXUj+uuDjasGppOihzO2MsCmhiLLmN544jAOZAnlVsnvuYPtKBd+pyqTtosZbGnYvmaaB4bw+q5f
VgvlQsX94hLYFgDD4wtTdd22g+VLq8dQvzfVMve5LLQ/KlNcdPccU3DBAo6TwF1IJ+d34ztvtveM
/38KvPirnx+A9yeNOtOCJIpt8TRxuKDbQeBjOzdoisOQ6jxZk5k4DqKhG9NQ1wKEJQSMp8RYN2w1
KI67CWXZOgooWh/e7FxfcgdSTAKqEaGRFgdNYpKZzlC+L9+sAEVELISr8kvtoF+/HXL46luFShC9
0iZjFAQzH4PZ46wGnHuHJ8DKqOnK3qKkPD0IpLyQ8Nk285IWF7EYsQAT+nd3u1Am71+gJ25dCskX
sCFavL9ydORdetqjZ+WzH9z9ufW2VvJUhVXhsOSNAoH4OwGrSxAhhRdL8OMuQl89Jw1SJ4tcoTxS
zrn8bzGIIMg0x7eHHe/LycnTItrj5L0FjU8aG0MmWqL+yNo9zegIIo5Pi9WzIfKNCIwh55l8ZQ6K
+8pa8uiDcQ99vo6FnDfubaFyzIH3ZRZRDxeMVHBLvaqIRgwLp0ImJBo2VLKfbnTbg9pPHV7U0xaJ
Pgkt4O94Bso30rGtRCSbSpEA4I5zHaXcgAoDRXE+4a9FEuyFFO9ZXDuOnNwq7HZxwcU939hDHZi/
Y5ZwCixhV6U7xLFmkfnbms6IUzMe57JAKP9Hg2P7z6DsyeWI8NneA6Hem1C2rab59Ajuft4SNHtI
izCWVlWbNGlVReak6Acjp5X0GQWDGBTfcgxm5uT2EQ9cfICs77iKjsWZmvfk6VR72B/NDLUOtN1Z
Wu7N+MxWgaKtq1/963rodVGNTSmUv/QwYOCOxDb1mBWgmlzrGefuKyFbJqsBYbXaYVM2mxnA1NJy
W2X46DnDFzwNsisfVi/cLD9DnmQ1r7gluHl+G0L4Vq08JADcTiMlKeLX8z/dBASAmZU0x1cCbnFK
erS5MNVK3BMTGbxgf3KllDpiBFIHhKxf8+RFPPtgbwujoVmjoMVS0+6c8p/wa95/39GVVE+65ZXm
+mxMkLLPN8ISat3Qd6Utn0zpjx8flsFr60nLplberP+Wt/2PcWXd6jcbGns0YArcGnhVrmRfNUVR
yMMAUz4tXKxvIEvyGik+smWTtBMi5nXG5eJxb1G322/Sbpvp6lodbuRNkJnxuytOvuT1Can2Hx4c
+bgetImmmi7Je61hhKBpkrqM/liVV3S6FF1HbeBxXA1mg3J5FTmumx+1lQ0+a0aLbrMtwSlRgaEa
mnR0/ftxGi1LtxXrM37jyLO748l6SE31jHQPVtuU0bq3q5IBWi9MddLGic04q/si+u0JqaS/+a6X
YXM37Jw/PI5OoQVkQBH2jSmSNio6FlMZbPwmMoZGbdimlzRCLQH1FA/BqhVwEJO3PP+30/Qovz9/
E0v3Z4l23nCfI39KX8eLh6kdG+iwZ+7n3ZXkIlLJNsqa/uAAWtGlmFKfSJWmJ6foJNpooAYAsTUY
haJGSkY0vLoLVs0zBmGySaloWVVlCJk0otnU6P9JN6SH5oTn3XKKi0P8oX58HG3k+0QEOFuC/biX
0ZiNBhpDjGtgdj9yd1SMqtr0UwzQGvQv/9e5AXtZXdMziAj2/z4zpyqMWu8/SKRWrDdAlPcyXyfl
xr5dqrIBYqRbtldfJJ3yfS+xIfceguuI5z6dzxDIQ6Tu8ZCywDn/CULtUESi1A3YBqxdmAJR7E2M
g/J38pA6h1tnprJzjFqRi1QATkJ5QiyprjYN6zdXmqd1B6uq3J/uBPwvhSd6KGWdOhCJUAAIFoO9
Gu62EFqbMwYftf5/vkvEnyx/HE8jOY24KSJsIUEAqIaCOhx2o9Gct2nPH3mlNCX1rzC5//sjgzVg
50NrJkk74mrM73RlTMUFX9Ovi00QRl8I19e2j6tdoH/Y41ozt3cvm1wX+X9ohg3Ofz1L+2uPbGGk
lXce3x/VLHEyxD6J/OHMfuh/FtVrrOCkhY8FveookZ6+Oxm0V4k1zlOyjNc0ZsZFZB06lPqtPEuK
sxs1eR1x6SmnFoNeQuzkTHMRm+hGsEOzc01lXfVqqculO4B9lr3U9NiMUXO9kS7u0zQh4MclOe8d
Z4e4Vs3UcvyqhZVGHszfXTf1hARxeAQjQuIbSsmxMGi3SylIue6jXa7qjrZwRrV+XgmPR07Rva9t
VoIVlg6WYKeGkobItRaOKRAHPPiu0DIQgqZVUY1QmQmiNOwdMpX+tuBSs4DLJlk3xZ6pQgHWqWk7
Ru+EE0ALd9y0tFOQUUmh9G+HrcWMzpJmgE03hCgzSOBYCaPYs0D1NrC4dzFBcy3BvhZJKIgr5yDM
WGckFj7YxNxiM2T2jbPAxmkjDSnlylG4o/z8RhGV6FB7hOYYkZ/OSkHkQUi04YOhTTHgBjRQnomn
npw0CBq2VXxZrGBenqBn2KVEmLRCElXmP10ncc2G5xnn1NlK8RN8ERP4wxgi/zUEAR621PE4ykVu
fdArkBZrKX62AFj8iqJf+6dx+4aFb+BstCUy7X0cA1DYq+ciul2TwyGu/FF+TxlnZ5vhx1p3Iz9x
Uc1vFgZwYwskqvBm3TUwTL8jVRsmNawcYwzNKKGvz1b7T7yJjhWo3LLWJA32n2HkbU7bH2OsBYNX
HBOAmNxya55wnCiPA7u6v80RN6YRZpaaEt7MxyjZZO7cZ253obM18334N5nYCk/MqQA02tewhdX5
pM1OStJugj5BOOzXX9WiFyyLdbs2c+p41AZ1F2rcvgOk7vfZWzQJUV4af5DOy7zbQfkUVOlRtQeu
H/pINC+CYA7vNjosHhvbD8fZ9YoZOMjBt2CPumJhOPnJngqxfDNBvg9N+kz0IJN17Nm3p8Utmmmw
wSFQP2KrtKTRCEHouVR65rni9jgIMuHW1Sn82bHwzwqJv/sq7UwM+p3LQj3OuoGIBqxgvqgQ6Lgh
5j3ymxSu2cuMmf+HK/MTf37uYVieUk8zl4zETsXhsf3aumR80pjLWEfdiaiM6l8+hv9XOkDz1JDd
Wd30a35SJ7M3t1EcfeZxuD3NBiRF1P1Viu8M0o0jES0XOreGOvmqseb5byOVPonG/9a/Z0M4IJ8h
/e76rvOtanTPow0xmohjJWw3BzGmuW/RMdvOuhIfMfpgHtdpVKR9zpQLW7YOODPEnfpcWihET2+i
cNQWCV1wY4GAHYgapNDKesNtZAGHknI0FXGE6pqCffO1yixY6bQxQgFDbA7XyDsH2hp1aXxB7Wn6
ADRtwQLnZ8NRU3qQ5rY9BWSHVM21xHTAcXDcKcGVnzsrgUtVesyrysXsb3SMuHkeAwx48KApKCK5
rqizbO23eCsVB/6uFILxU4ANAw4Wehd8y3nhE7/RgtE96u82tEjzIHPh1A+gTr8Gv1TzEH/PSgpI
9kkOjRXgLCKSh8aU6gEwy1vgN7GTfT4mr+CttnfNH3JPpi+H65Ay4UDsH+b3EpOEYYQm6fdKD2Bh
6prFzClt6vE/Mjcf79iggekvN5URN8AJRaL0j42Xr750g8Ix1tIjb49Nvr0um5Vq7p65yFDc3+my
oepx9uWdPr9uloFrD8VjRZmSBMb1XHNgG0rPOfh/klUO6DB09PdkrZ+YEETacqrA+LIlv56cKK7c
9Sb3m4Bki4/hDxW11OHiKsiZHPIwjrWH/29b0zEiwqQflmz9vG+w9kTQSfpBW1F3xS2ohaFQggFX
OnYklL2SqAmhrpHKaeE+jAJm4l/JGtokKd2qZibQfv1QDU28ayXShDTVA7wj4u+251f5GwA8+xD/
jTrf9y8MydeVSReV7BWyn7kis1MMdnKqoLpo/6jGaTsiWEdgS27x3qopN6OfV8srjahn3XnikQgd
V/+AtwlB401wIr2N0TueZ6Jf13zUFDxI7bJxvM3qRyV0sLCEbs2pOKlpuqStwkR05xkTBpr21nJx
DM7wASe+uoBB4RGYil28BTV8mR4ZB9qmVrTPZghRDWXxsFWwNGZLth3TKBHyLK9CdOZFiVTGRit7
r8XaDN8itGftRhEO0D5NSWEXFnHlGCycWM789ZDnnG33CuaAGFF+6mEyWjCCpuQmcVgj6o7BHN6Z
v4WK757oo+p3YclK4iDpy4jIreDdOFdxIIt6QMxk30Kf9/rf3uZ9fyqwKjXupt03O14baQouGhIN
rghktOW+r9vxaE3toNE0pl1vVGw88TZ+z7ovdCE3TiLihu9R3QaMdxtexhTn+1Ralzh+FyaP+z7+
x0+LnhaiZ9nlUzF2Mek32zLQHhtbhWNM8MnV+9f49ZSSReWKN9Hd55hQAR89C0GBkf0GFrOHasVJ
gv52EajtR9P+tVUFowUkO9t1tfud310AU59HTh/Xgylfkyz5uEDnYKfC9le/CquBmhqevfgbb8zu
tL009XzWotLl+7QoVzvow3bZwg2cc+N4mJAA9TZ27ffasHJl3+b7z20OA4WOuU2hWv4CUVAJbC+X
syx1cwf4wx8taJw1ZafViukpLkJGCH/Wskdpffb2ulQ7QEtgg2dRq4I84UtPX25e1Dt2JrhoOfMF
yy3fBytgpJUiFCAw5Eh2ylHKoul3vilqXrg0glbe0J0BCOJ0/tPMsPiMttHloQ4lw4iRlzVOxCVX
VVx7Lb6JUesfQif1nnVFg4BRbMHQs5fzYGOBO5DiyozmsDwbCIaPJ0ET/LbYpDeHiYujJOWkgDP6
nCTxNQE8deyYFmPM+bvRLgKpJUZVnnSbUKuBGY7SOgjK4xZhmekLLx801+bIYDNraXn1GEansjqJ
XGzzpklSH+A2apYs81BQjkCHC7iau81i25lvfHso581FzKtGTDyGhb2YN3JOLpD9TNEvoo+eUcwC
ZcWXRYEm8IYXqFep4otk094Ol6qhMD23nuK6tYbL6Vt8lyPgTAgJnRexX5Miy8oLxXRy+qWt87jf
79K10S8AwExhXgkj3WQJU5mYenNgjzZuf3x5+Dp2aBQ7bGUPyZ8102cDxgLmUaAMP+jAOZUTZDjd
0+e3Q0gqWPAQceePRSXPDXNgfEn45a4YAULfn9hThWce5FC8Il+oxFTlIOdowcFajnvBgKb+XQx7
qUqz5hVCBBU5PYl1jmw9AC9ZQAyy8us71Kg8lpU+pp2Z2Vl/IwrZumipgIbtAn1OEqlq+ZVSyIqv
LgPY6clBhDRZlfcIa+J6PDg8r7r5BxGT0+KjyudzrDFNJJVn+EhEfrier3/XKKZXUqXztvrVn5wY
nwf1JLVJpnNloLUV+0obp0P4JbGS5CPRsJoti3JVoUP+pEzwezaPrFczjET9MdiCAw2gRKxLubfW
y+LLyk/u0TUWhkjvfP68yQuE9pgMRkgJdGaoXx6s4CTUcXkXC6lNaBTY3UL1/N6Ltj33hVRoV4gB
2lNOM1XE9AV1w/teM1C2uPfKqGv76Ldgdm9bXGkSrnTXo+7BIjuY3ZNeuKtQ9HGff8a+0Ct2xDc4
WS5ZpfgSUjHVsNziKVfHYspGjcDnoN/AdUrdEypwjSDiYDWZJDWlgoAogBRoLWGZNXb7TO5HJWfb
U92hjg509Jwx938ow3SR4K72akd0m0D89s2CxkinrCYkAamL3Qz5WLr0YjXjh4+Uos0ozakqkjj+
mfFsJKfmZn5AMdtVFNaORqiIX7Xcy8QIVApZcgzADOFV5SJlkhk6aYsVpUMoLnab0+oMkz1lwIYP
hSTLlxN5X9ubYHrC9ll4ErjMxPbF/4IsLYLDoTyF/H0ceP8GYQNBDBhRiWi2LLsv0zInso3Fk1ci
JAcg9LKaeLXhhL/19O/eeGGhVE2PqWnUr7R7nAY6SKSPz+rJzTvhaYgtqh7cCDbCR/c/uZBKcedz
9o7Ob+2WnpiDQkhjEemX1X2ps44+S02pXdioCdLotPJglAGeOEEcqLBzxUBHoLtV0mTUHd2s6c45
ZCIRe6QrSXzOnbGOJ+oQ+zNTkzxGXSh2AbBXCXvEWm3xDzwrh9hqIV2G270oE08sgQoeTLEnvTra
L5jw7KdLQDvyMlr5Vgc0FE8W/HfT6b7oBzl9ufl9r3g7BWrsOw5eImiqzd5guGURieIh1ksQrF8I
BXmRt/cUpvIEll6Ope/ctwM9YjE8ZDsLjRp1OkPl/Q7tg2DM/Zm4X/4pTr4RhS1pNwliANYKzAC3
r0bXrsf5zfUprc1YSWXUTYIZC3GBYcb5q4TjFImLSYgVkiPBHNNZhcGF2dgoP0nO6oryStOm9eEs
PWw2AtGu1adt4Z7yNB0SwMUe9++JNH9Q42jUB878niR1DO7nTy9vdxU6ukhY8e5gczN+aE/nWHmj
G+p8ZQh2gUm+cStrF/OaChhi4+GhY0VLS3dcVI6z09HtUYh4IV94mQFlT11svI3TCJT5A1XkXPSn
cbNl6IBq+wj23UDy8dX0uFD+qhTXdR8SFR82KpttD3/Y2jI2s8ELgBEydeAu+AKmpkhkTIpLP8Xb
sgPir6SSGUXtDL/lhp4mz5DJ7Yr+wXTvAhgzB54PtJZY2V89Dds3b0wo+FR7DOVGhWCAOsPUyhVZ
iAy85N2MMyY57LmVZ/NetTt3JH/3W46nkjvlK440VAzbL+f6NTQWxdwnywiw9mnl0GEhNBM+Zleg
w9kq2WRO+AzyHpNN19APkH5a00iS/EN7Q0hzT8j2i7DBDFEv1aOzelfwWSKtor4HFzGCnQVps2UC
W7mZa48hvbawdTEVFnPMVMbG6eCTRgfmdmsVyNfl+DTRhkq8MCWDyTT4AHfiuwNaUrNx6irlnc8M
ojjHQIu1ijJQbP19X9wDmiC1n2BgXqKr++mw/5rNoTDJYINuQhPCT0Vr9RuCpmHmtqWHvvb72ahm
dqkiQyEsLTZ58EchLyi5mn6TRjFOy/ATdypnKeinEc8jkYgmHK5ABfsequ5p0DUU1UQM0HrVYBVQ
GfsYD1EeNT+F2XjAsyIKJ7oJjabhLsol5nz1o9UB4J32qrbS1Cjg1LVx5MZK4HZZf7nHCJ2+SXYG
GhOigF40c/rHAINA8gitpkU5pIg/LIHRlSwKypaG7cbKzD5edOiWFzey344iEKqOqRcOmSD6Y3+R
cVP5R404LqTSfxWy/uCtxvetnJWJQF6eixVn2nwCVQ1MyaLiLegPuE9zSW8/Pww4ma/XnVZwFKrL
op1h2hHDQf26WvZV3Oq/E7rXY4RsDzhgqSalxot0IJmbDawX5M0g++4adI0/atMOsMHbPD7f6z81
WBk1IhO9NzbWKwtIYYcEU3fM4siXM6LYDiqRmVbVfN5gx4YV55M97Z8QJLLzqHJAEiNpo4cAXK/z
vHoo4OoqsdvzhsOX/xyuMu6IUAukoz7JHExwtV08AF0XalcmCylnhURR6WXpLV3ezpEaTsxKn8Nm
TOC0kPcRE+rbdKKrYGiwozxDHmkOvxYEM49g4vHlW/bwZLx2hxI0MWJqtKlIvjLFPp8wkl+xz+rc
JIZnRX7mkCLRPOgs852x7YSfvGhdMSMChDks/2QFqPPVKkgvUy5QUJR1YnLWF9nxfIgIkvmFc0+f
GsNTM9tnSdQLCKznkJ0bw3eZ37mVMpKK6fMQW6XX+gC2HJEasyYbyr6VcXHX8nU5tuSJE7TcNLez
QaSpB//rPLePHP42fL/SAky/2Y+PHAT17bi/CY2nPALz6g8+CV2UyQw2E3L539VuuyPaZ5+/aTev
OhKEu4jQ9tu6i4y6Oi/vBycbyXSWPEXVneShECMNqdNDpDiBl9clTYHe+nkO0sG/+E7QZJR3SBqR
kNtR0xXfuG61TV7G1V9133HcNZxYjeRscEnbtGUNJWJMQF5arC757Kd/SV5YJ03PckMd3Sv7KoUr
Y6E8FmoPhoDYeuCO/1KlQqdDryz1Bp10Fyj+rS16n6r3hrsxsXZDF0fY+PuOjT2P6gzQ16FgM2g6
IQ4gD8RjxhN/W2bYh4RG3/FJhkK9vtwfV0GgScvjSCdpgqXn6A8lJu3ZBGXir2vOPvoyORe2gkWe
mb8jd2oGAXUnjaTEXfO8Z4BP4UNK7lMUohpVQiYOh6EFCIoJns8DaU79zz43/d61qnoEe+43KvX3
W503n9eN4NhRnl4N6rWpUP2M4/oJN2BdoEcxALFmSz0e62dSFjoUGGW1sFRYoghgw/2qeY2cd5Dv
Qz5aNP6JSQgtoRRek6Va9PanvH9uiKmynQY5p+IJoleB+U5z39P9sW5eS0eeyKd4ArLYDN+XwLG/
A1gBBvZJbx5UeLlSJZHUV2VVSOSHyWysOCxlt3me01xgnQBfJ/71uzEsFHYILFKibZtMOqjmJUFN
e97GUV92CdQL8H/VE8vvJWyIWxfg8dQoOKmMO8nWtM05nX7KXDc9UNMhCBHMasnguqGAHXUMIhkM
MHR8Wa0yQqliMUoe9pi6y2K960c94JyNF1OtDHtIz9IMTL0V+uEsVEgmNZ5edddqeWYzhFWpq+HS
DamKRJvnJabLVtyasWFahDKkv4zqQRvQB/WTkTe99wEWVEVRjh+wPAblf1GDICUbcq0xEv+iEuzT
HU0+riqXE92TE8MMO5g7HrSJnIVDgszjmv2IwGYqpMpLFDUmVb9Qjs+K8R03jPkxu5VDyMZiaK4k
ShnpkakVGajaExSlZnN3LhCdiZECPfQa6FkWbV41JXff3CC1pBTtvsz6wpahE9W9dMc3xsvLY8zI
X37QTLgR10d8wUo6y1SG+K5Z9lTJt2u8TfW5YniqsB2QKJuT0SVf6YAZqcR8u4JxpSMdN9Gj08Aw
a6dUV1kjjUokIo5B4Lz+Qjr+asuicvNAnAf5JJ7himmf5aW7XX/nJ4Z5a/RBmtCZwLKNFhPcvv3W
TFIZi2IwKzPPpOKGtlyKM5qUQ8RB578DI49HyfT4zSarYYexkv3NlsxAtvwl5DFcc+C9hi1GE1gr
xk6ryDr3TOf2Z9+CVXYwNViphoLDeQedCYNcWw1MKuxtO1nucD+QbeoLVQvLxPsOw9csKmqbnHda
J6rPensE0FqVkXYTyW5XK3LBfHsNBpNoY2MCJ+FZKah6qCkyzze5CcnKaC9rTjCvcy0C/QL+d63q
/HsZ9b3H/uWoVns3pN31PKve0oMzPmbC673Cqhidn/JN5rb5YPhf/ejsWl+6T7UYp2cbhdv0QlaS
/PwsNjGsx5rliPF/akEE7Q+YyU2GaRU/o7T55AHByuKKL+yE+IEhuzeq8gLp/NquSE3rMo3t+2Ha
IbXjyHNgwQMRRKESDeCnPRVTUOjMb3V3xmoAAnaSEufsKF0Eap/Qme9QDIb8fhx2VkN55Uv6E2uu
fkxTyDcIPDCTDZbpHn03SBuWTJl4kbzXU2/jXfLx7CPqjFxyCKxM5WWgDsh3vqDIlJh+6JuAcRji
J0Fqkc06gHKyjc4dkVLzfNDpo8z/PVQNKO7zqN/j7h883/eI9+hAAeV1hhc++CHWPCQ95UOkkA+g
X1DgZ5OB2t+Hlt/C/NBMPHpQswcPdtaFUB+8wMqoR7OERp7LmYJk75JZKeDHQ8wLY1BKKq3s9LzE
ssHNLaeHq/ohemzB1KyzuX0XbVFZdbH/gSLnACGCfcQcPsp1XLaSY3y72fc7nWsW83ZJirFUsf3j
WIHPp2W3cS416FsfCbfkGZHw83QJeWXgaTLRKCVPRqpon2MuRqjczSayfjjsy0ET1VIe3nBqwnxf
fNRptcgAIhDeHAAG47+dN9nuuExSxZ2yT3nhe3DlYL06hwv8KZ+MPlBFmbQ9LgQxX49a+8Ar0wjN
3afkrvvQt0EVhorJOKEDEMgQkhAHzRq5jiHgdGy92AJjWlWya0MB7S9b4sKEUH6nt3StqF8hDd8d
pIGSxiux3wk96+sQQj+NeUbY93EEBBiAx6i+kfI2xPVinKEz94Vqj6J6FGQwy7dQCL7i933Pffr9
zn9cN6rDREhRUGi+EsTsZ3fUT8l7w8kQBtSluUpRbO/tvKnOKgjBK+W2IBlRMGolNix/nyGRmGjr
WnDw7QzFt0uY1wDo8je588rZKNymsUOF2EEnp9fFOjz9ErhSm7DzyG5nfezS+m+jYu5mvBa7qeRa
gYYLXjoqUHkeB9OhP4C0TrUXVZJRJOKj8TH1e+Vf+SE755IxCzEbm+xMCP+W3G0/bDmf0LJxGvvN
30l+bCGh2m1gTKnzBg3NKyflU4kgBH4O9afopzKykCSH8Cw+XwQdbeDil1NdVQPyfWENnhG1Louu
qBeTkTKKCZoSuVqr1qgbitO9r7bz4uMhWsyuLu9zIqem2WT4lnEGvkEOwSV5mMzhYCoGAI8f6sRw
Gg07ctTsvgCqdN5oKYfdFBsTsCXUYHE7KIBzGPTJmuU8rmpnTlnbJxu6SjATC8MezN6lxQ3A/uCU
YZ6AXjQ7+N7f318WvUPVuRV3emGmpZpYphyCbVbN25wbQQNHmb+EWOpcU6exJ96fJPzTxcSz4BoP
fD9eXV40jWi2GW/VflRpV94Q6A1Og3udU/0C3ncnmYWWfZvZkfl8ZIjle7jLrSnwQX6KT+RAuqd2
FgMgijXYA0LgmW8PC4JfgW1AzDmei9RCEyH3zKBucPpZsibR/OLF1xEfCBGXZEA6xmnGkfeXMx26
ncjJR9VQgVwTmjxL9QdEpxyiYY7ND8qCplVhG+9o1lkqh6jwjmVbzJSRrj3qKLKV0kT/YBcUAU7I
YO7fiwKmn6yCcuC6nKKgMNsCsKK5frrS/+76tU2ypmrt0X2uCaLx28iEpiEpP1h+OLWZatt1Kqq+
3IXv8QdeoHXCBTEbyXDgg2VY5LXYBPnsUC27XsesluORIm7dNqSAJ2oFjK6RxfgGV7XR+ssrvFd8
qJaxxlf7KUi6lS1nBivwC6DHoXt2Pswf4C1vAdYOogLCvp+dd44Rc277J8altSi9KJifwzulYli3
cOjWugpsZDrDf94OiU2MA80TxmraGpg2j+dpEB/cytZj/3nXXXv3gfRz6w7dswgbpP3vmBjXi68s
E3GpeQo/7Lbs2Ae5gcOJhOA00YYFGgwgO12m1EwDutBsK95Kfbt3Ol/eHqzJARvXoCZ+aIBIPW/E
dUPpdj6ohPGl+BLZmuuOjQGIQIs8+XrgSwL140R2OBy1cl8wXG/A7uE+QqnuqzzhIk5+USAL8Pi2
H/rDG6SLH+3/X/CT7SIpwyo0kTkwp0eoaKqMG8s/wh/d9sS4uwmxb8/sQ4sY4BV22foZpOQNt/+1
yrUyVVTrmIEmc6/T+E/oUxeqw4xxNVWJXt1tnUaP8tWQRrnI+epzV6tOwq5a9bnYXq881kxk8pIp
hgQ4AZE9SLLGWIJshVgwaDh9dCbqzICiI0LXt0ofdRkw72gS0GFpDkQLmv4SBylzwLAeuurbeCQd
WrKmm1/OuxudLUHiKCChwy0EE2VguA1rtlpmUSTcbVQmUHHl09IyOJduko8PbknnYelXqb3cxCIl
hHgNl0jnaWHf7rhQGFXqjqBWCx2dzLHRgN76jZM5jyNEoWZZY4lN7/GT4h4kjg2CulFposjO2aLt
GYwu4UJQzjqAz/Z78qiFsrDc0ByEICn1+Snyo8TU/ysx0YQcTEEQLMd5d2ow54nQbHO2Cqjeic4T
DGWp08pV7aUVDouUIX5UE/PpCz6za8rb4KqUlR62AUjB7P1YLYa1SPXHeX2yvcLMdhHq4X/PZ52D
uipdqxbMYvYT0q7/QqBB+ygWkK+KdUSLf4oygQRyxt79EBAtyi9g6MRQnADFLOmgTfVAShi/6xXX
WbNbg/A8J/XJ8VoqorsYOP3eENvK9OHdm4JfbQMG2wNylAZC6lbnJsWgdxha9NZg0O+j6AZcyFGN
cNASU1r3sORbSCF558VPDLjvYBxUoK9wYvlBhRp40CsrfyEm2RmOGcUl9Sr/H4sCx+BAggiDpPsg
D8Ddupa0m/bTS8y3uQpjIDkD93IDrkUiyp67aTPrc7Tq0vJHbrsOnAv1BljUT4Bj/ghs2lXojVCC
l38hihBlwsY3w0HU/WWFbfe1jPz1hDFROMgVFk/rWDltOpA5pb72oFmlF0CWSYHkgiPGI0yUiptp
sadcbKHQT+zY2pFc2r6uQ9gm/4Imt0rVNe+yriq2aTwwKkD1Q74Jirv//47xxRsFu4/6esLG8UcF
tPVRaDCLuwLFwL+JYcIKRDea4onJr7EQm7K8wkeSq0VN4Y3fDTeCqZY4nDFcifO6RmmHwkhnQuOS
3ZS8nFEdROJJmS8b4tuCNOXHdWN+IxJJpUWRBeF/InppjMDt27lXbAKEGZbFEbMLVDWEPd3Azwzw
dGldZt3DGIGDkBcC7r4WcBvZzGGe2WvsMCY5ARX5i2j2fgiqDzxVPfSsF/x9xJyAWbsMxtRnlv3h
c9MD13fmVUJOcIW/XywjDrq7XNL/1adXjWiXTsD4kF3IqQLZNLUj8hrHZpgU/jpCkbQx91KyyusN
VqG6Hn0f0GI8wZ2L6UnfapDLH+i8TyFRUcUKXU07E2jp4PMjUSaWXL1bu/E8uJm9/JCilSKRfCCg
WLFwKUFvXSdo6AOyjAu9rJFGGpDG4ngPw6xKUv/IGOgBdRFXFGD2KxI107GJMHCSNbUG1eVSN7tI
+hNtS0s3eGXG8PXKlDh60gkSw4M4T/fZmZ8EhhN+sb4qjio1wRWFb0dIjccLIt/TE1LZPXY9gtls
99/TEBm1/Kk8E3Mcui+cJunWxjBCZHPeq0twdy80qKdZblhxe0Y4zNdBOygv0YjDP5MzGJPkNwNE
pKJb8IZi4t62BjHwSjH+iN/xIIne5r+2HbvPrS+Om0dvYWKac1gcrLM5+YbwkoWVyctCmOKbLE5z
0I/ZZTPl8GuzZgT3KdzEH0XneJ/TJi7mufB9RuIkoKGZlPY2EDSbzSiOaWKdOzaT+8h5lhLm5d96
fIuE03aKddAc85wbY8W/ceeck3yi2++uE/VTp00TtlNFnzhmp+Rf9bMQYwGAtADRD9TPmANl1QNH
ekBY38TTwxaAQ3ez5i86OFc3J9mFFgzHSOOV77Mer0O8IfumVeUIYtYPNbGUYlvhxcEaHrA6Abqa
Bg/fCiI+Pm9BtF/ndgmz2bdhY2TBqOSOBW2LBIGs6J9ZIoH7K3TYqe8Tcji2/uRJzdierKIhYSUL
0c1QXIL09WOyuGinwDNHJBFSmb5ux+53uPxfLqp1+WwN1+Jja3lKYL/bd7LugeKJQg/gvwC/2frw
Sc4GjDkUjek39kH32WwqRTMHRz6aEQxvLv3IbztCu5SPd0wSofmAAq0WAt88AbQKBkb+pXCcUnUK
6J9bq5vzGHkOlKB7Zma36VUYcv747hJ6RteK3LnT7+Z2qnalhGawDwcykE7fZM6rWVaBHS20koAp
OUeKoaRDNCJkmfEn20sdNmHkjZigKqRQU+WUeBm5528Hbo/4K8kpMnfz8jWAQ0nmvABXZlAgZQQR
v2B5LmwgXqAGNJymxO2P5GzpWrh8NW5yVPA45QDKTXbrzNr0Id1QcFiupTcFiigjTB7PA6WKEouF
Yw73AJTO0kfW4EsX+Gd7Tw21IeUMMOvbzygGRblRsAjwHlnCqU48gMWPOHNZRQ6dNmq6NqzdP/fy
2/wIH2XSZxGxRxpEhJTHvvY4g3hJl49/fE907tV6IE1I8DvDxej4apYWEzcnsch/9hB5rDlEpDwm
plUrMytQuYnpOgdyKuLMLK91iFeJxxf+YcnHhQkcLZbHLfXNblgoXuN3LzGJXLQfndmcCS77Wzs7
tZpKE3ck8f/FuX1OWck0fTp3GGmegUqNiSZerHqEz5XXtzrbIpWTbNXZc8jZ2gqDTLdKgEzDBViV
9lOLMeYMaIqkYDgEJOMt1L3ShMHhMrs/lSaGWcECDKwBlhaNM5cxq7c+4DYRgGILvLTzjBLUb7Y9
4gaoDxMc9mw9a8wvyEvFVCx4U8QiUDkAwkTLPd5GFdKaJ+5ova/4WgVUbZnvJXH6NCPprbl40iOK
KgEEqJre8WeXl8Ptecnt+aOfGpv6ut6iV3TSfjquIyJK7ddk9YhzuJFeMNxx1uHQTXa3vL3D1fnS
jYp5sCV8rK0GlpKLOCEDDAwsWEq0/CbCzn7YkhqD8AD3HxvTsUUG7sx8WhLiIwtpINeNtaXO2Xzv
WoJQFoAX3AVK8VV2p3DQiHFm4YNhFAtpRZYi3c8UQKEa1LDHoAaLN96jpsEg+CGeKxrvOq3AmaLq
11FwZDKDZNSQJonUrFsZr89gmZmjIfyXhFNPE7A7Lr8EkT39RfWomoI1MTZpxuugF2P049+44gGP
ePqMCx8/hbyBX1mUolG/g1Ktq5VtiUUmT+fLimTMsGzUxC5roFAG3pp+5XYsnAVoyLxbw7F3E9j2
60fNTCbQxSRSYJ+tQJMLAmAcWnncv8ZTKLPMpoKF9P8AaiBL1c/OlHed9ocup5Wd7XNvJ8d+9ueD
8lUAXVvSl0Z1/vmpmVesmkFwpu2/TcsFq3FMJGur3A6QPSfKaazB2IE4WQ3IXcyU+bjkps10PGYD
SGu04rGfkJBbwRAd5xh8SgqGJbAVZRBzpZZr+T0h9sLBlsVVt4lfZUwNhUl1Zbqci7dNlTdIOXuc
jmLJs4vR2mPStAAnR9jym85M/gJ8ou0jrYFEP0goPCgLFjtlCG3DiW+V2+RRRnsTy2TnfXPXW7WB
bo6E7r7YB9Li9haGuU35qr5vU/+/wDNV2155sxdsCFeuHhz7lsgk+dRHpr3lBgZnb9k6WLYpEMZx
KMgtzMwmxAL03Gh0QvAvrXEFyjtIP4o42yKRFQVDuW9F6ahYVSLJM+E2IcilkqY7MNZCx4tyDWIH
FZVPQAzUvCvYpyHB4Vg1kJtlle1oc6bIsQc7l/i944srOvjwpAGSmCcYbhk9gvoE5OiPJlODrVAp
J2mGW4ohqutmZ8pjn47x7U2UQXentiroZj7RaVybnN+KViaxkWQqzCFJ+jfREgDyTUE96wZ7VnGa
6wHHy1iKv9I/2LVuZnHKRD8rH9sY9IKeNTFFa5rtcIqxLjEcjpFAgt6ZsrqHp3BI5+SozO4kfTei
F7zRdeYvWamGmwLFv+y/Mmax4C37Ozua4hcf4s+9lKejKC6pCIDtum2c1F+JfjYqczW2doXHs2jF
ANtipVBiJH/vPqJauUitCRu0LYuGBxH3Z3/UEcgwDRn6kGiFkDgOLyFej4MTp1TSwfukA+neqIDu
etFnJ/OJurPl3Dm70FA0jHLb1N2D+bpB9MBgCqoNwyO2M9gh9+UbnAXEoIRrSnWyeATwt/YNupLP
5S5ZX7SbsCV6Tc8Hcjq6q9tp5wUMgMgw9fNO/4naHy4IvlgdODyt8AumiukOd5nu6AFY44kwSx73
oRh/9+tXZNPx8cu9DtfFdfCErvSAoLo94zo0ZItBV6VFwA2XOzKW8TdQtI+HWDWEEiBr0egMkLxD
n79bDqUPC8Kou9nF1qbVoQusWE5vXjOrvYm5PGQnAgofepEtJrHSmSetzaW03484RgX4ArLmztv/
Ac9sxf3+cMIlwuN6h3oRD9NJZsvddSYv+dFDGdnL6zC6SslltMS4VAJgp5t+aY0OM91/H0vXTYY9
+2nC7MnMAw65Tk6OniULoG5tR4eHF84nynhxgWM3bj11cP8GAbisIpnutB/kl4dlrpyHq7pCgdVO
E/RJbPK5JA/5hvbjjACymcpOmgipqYVaWFkBr5DOp65irTIDLpXHV+FaZ73ZyxqdPx691okXLwXD
pfdH6osV4GpeBqgJz4Pbi+erMPqz0l0HbxR/2ATajr2doc0JqGwVuS3TYR/JDPZrzB76V6fJOEtd
+v6eh1bY9+HL9UuHIyIjwQDD+AGDhDFjWJOdnLgTCHRDnZEBqAQFYA+CbTV/vBRa8sHKdiGMN8LJ
NwKJRfzfywHTFCW7+8WfkTWjRHQXjYHPNamcICx+5DyQM5gnodj8LTpOZocVYDSnwEALtMRf5VHQ
Bw4kiwt7XMJl4cSyw04wh8BsuVaGLiiLCtsNizt+POCmVQVMZKgg1Tx/CXtjg9toP4QDOjrmN/S7
9PUNoPhAem8w4g0mjGZYDNEqW+tda1Ymi+q/t6mzDOZt1YIrU2eDWbh22cw6I1CMCe4ru1E6B+Db
43KsT+09WfKfC+z0DfFxViJECCTAMnVJD+FOi3gu0h1JGadZu9VZRIy+mnybzCrSHxmT0aeHbCi8
Alf0yp4w7rxCVxXDr1JYlTGcDka5TcxSCHKxeV7e8bp/fmxY26RfT8ZnKcnN+W5CSo3B9DPQV+gx
8sk9r6Cf1+br1ijU9bcpZktjk0BPHrg2iT0NnUUWxyOZnsLpjCf/wrIdLPzoTL0vk4IaMFwdZhtX
NRjb6jJMQ5H3abYcuwaSYR9Lq+h6B96YIZsnueRwi0Xm1VnARREbQgJyeEGbjI43R+OBRczpyjZd
ypet84Q4hYfycsEtDviTBq4dpWi/aqhMaDiEgC7NjlR76Ksxiqp2ndex15NWpuaWt9edl8UkcsOM
V4UgvhjSRQfoPV4Axe54rKoCQUUYNWdQ/oTawUpF70rDKd9oLUjmdCM3uRDm8dp7GTQh/zWyhREv
Fdc9RiEQI4h9cMQhRbpSPeAbt/LX1lqSlznWD9Wso1xOwLtDYhOD29IxPCkPWrCzv1jxSZ7SJ7PG
EukQJQLr1u+o5XpbHRKG17YMSHzdhqXIbmFS9WadMyXW1IlrcFgJs6APgCmSO2Nh4x/vxTVlvtY1
An7ErMDRZOxNHNtSsRlC0VozL02WJPovQ4p2rAV4vf0NA5RTiX2BcLDy+GcrEVxHe62f2pRwtz4g
0Ej6hD+kFB+1tYcqeqjEktAD7BkUBBbGyqhY+RRDhpEh7+pZEYr40jJXksBrMI9TlvWwqyPQKnls
t8LS9vLaIgQq4rpQykTc0CFfWjukt0/VsKaq8oyZue0b5XglALbYTPDGGZto4tpCkhHFpr4DyRyf
ROhcA9oKvTqg6iUZWgvmtG/uo7JNpoKHiebxtIUpvt4CzR43HnfjUwGJjS4yfstjegBXYXUOZ0Pp
Kn7NmMcCyz/N6t8TR9iW/TVhsdtolAWZWJVi0yXyhxSYTFCovgzZTouCnd5rBYreegvBhtY3gHSH
LKz4FybLPQzdfG+vcqrrnIWVHt3AwT568qVQUo1g/TbA/AGNrJ6wEy/OYuryfQ5hAAmDt26pJM2f
yAnzIoVYYhi/qDzlwE6OkLnujNKWOvmGV0UtZ1N9ncVVyOXKs7e+Z/4EEfxvENE4T5EB8gdleUuM
bnaySRU6gs4pxT9voddDzt9zqXwbxBwSfrJZgWwxvzlqPkWxqJ/fj9dPBjwSOHi8PeHHGbTGUxSZ
1Znaj1EJmf9WdJ6b6bHeLVWRGmpE2CeYa37wEWiNuWBlituRI1mwDEiRmwRS5NOyxZOT9K9aL2Ou
5NKEYW8c1dKAR/dEuUJ94L8Fs0H/jJ4ZEZCcryJL6aNW9oNQl/PscLHwvdRmDGsupXsGpI76qoEm
MiZ+IuCZWAeCQEAeaeG/rCE7VqLQz+PqYEutwLsps51iQgujDcVx/fdjfJQrr+ThWuClXzKKESbU
t7jRi+zLVpIrLUy1TN3APOUkhTdALOymFKpbH9xjSmMXUHBtgKxD7U8mNoQ83TAPrxVStMtr5W+E
Fs/bQJKeOV6QPhmbJwdcp+22g+hVk/mLWf34tBaG1xqCRWagaUqvK0v+/pnS2a5IT6gxlFuMNt2M
/cRtZgxIwnGQ4VCjZ2xe9d1HTIt8LQVXa7Ugoyj7sB/3UW7LR1hOZhS2MujEvIKLlLgmwiy8nCD3
MN1YjG5MYqpLo09KjIPT5abWH+/mXOiMSJK+NLHkZlQI/y1p/sVamItnR6r2Dc8j6NXFV4hDnEBq
DwoqgTzFj2iG1ubJWFO/mGGu+W/pMfGUnCkwsUFWKD0ImvoZo3Pn9/UwhJY6/XCKNu4/wZXN5uS/
4s9dYMrxlEQw4SsmetYw/GfA9w97C9mZPABjbWf1IWKQZDDbBavZrG48gCBXrOmdeCmhhhavasnU
OhRg5/mCXtwp250Vd5Bj8Kl9mjPYlrH5auosVAstHSKS16z+v76P9lPb88uxPqRKj1z8mTC4hK9w
RmS/a4APQR8c22EqbSFoCkCAsPm6d5bSgAQE6tRHXkWhOkiUFis0OobUYAjpZ/kGuSDm9GWSUYW1
CRHG2/b+RW2FtlK8fGW5wm7hAejH0P5Ral14LdnAWefhOEDiqouOxCUNA0xrYb1bjixaEDCX+HT8
ZnmTg11MTqWe6th9EYLSwJqzjy7L1auN5urWxnHpMEDNDuXrvdxgn7IYkE7dQdsGC6Ce+OPUokl9
P2OUbWsYO7JRwpQk4kZ/JdRwaw9gQ8U4uRA5S2v1iQiJYI/bHRXKXAFfH2I1JOLuzdmeJewvLj/3
0GqRzp61F4M2onDWN18UTI44C1zz0YdVTR/kQFO/rhhFBXsYkminZVGUFP1urPStp2kmZfNcpBa7
5FtyOo2+BifLf2LBd2zyLB6QzX/LmvJaLuJTldPsNLB8EU5ZgTZEMqNg4M7svjiBtGQm1kap5VQn
5AD01lt2mp6PJQQI6a6DE3M+xIjurCSdJfY1do80C4TeUTYpxJyodI2Q2peUjv/4myjRmzqC70hW
ZgNackUkSZxTxMbyMANQS5JTfZwIhf1mJRmgE9kPp8SsQLl3DEKv6Fel9Fi4oHQ9ZG3VQp36xQ8H
eV4AfXac8evMK6X1Wvack+WAOsYRaMwU17MYAkvkm9y8Gv+a/Mo94COmODPf2xYa8rD99hbze3GE
QZxOAOxz0xc33BcKSrz9k8v/x5kEUBgjUg4Mm+qxX7WOhvBAhRfqbNxV4a/FG9CabCfkHSJHB1mY
1Cm4O3/h4jIdFkBO/z3DTvX8Jo4LOBlUTXFBNvLPSbvyRbd0TjnAg0MD/vjESlJb1UNVSf5CL309
wPozXw/n6HtAhiRH5s+nhpNWG9+aHFSjU6V26mZJFzWhK7Ln+cyOZZ/J7xCwr6q1OFV2LW6VcG8O
8bKi9qqNU6appk0X2EAfvGrfojGqDha5OelIQhpIcIx8ELI4y9eYxAJIkdnlGbZuSvhZjaNEbvWC
eX/X5zhRBTZqdnqy/1d/QijUNJXsYVc7TxbYcwvDUeA2IPLwU5EQ4erV1Y50SbPK7NHJsMQ79kJN
WrfRJw2iXEscSw0F6fvmwsLffXwY3HPYh3lMcbpv03Xq3RHeB4GrNwed3eC/bEB0A52EgjcL4v2N
PrUt2oYpkGaJvpHcZervLCeXHOppQX1Y97b8kckn+q2cems5XhSiGH42oQ1iQ72b2zizveQb8BQW
re1JMbS70UW/X+IB3bx0qZfEvXvolFRSaNXqZfqhvb3jKd7qrRwOS2novpyEjurbsywZnLxBS2Fe
rTgRWwY84iOrs5EsSbB8kpAf8se58ykli7Fg+lcCKVnpOSXXKhKs91RbTMKMKrhKTpReVmDCgTFk
TJLrWKqTSPNmc7LlfknSKOqjsq7dKK01Myxct3eH/G7fBsT4GzZjQgN90NxPQxoel2e6QrMUQGkZ
U7L9EH5Fhheor8Dx/YoK1LayaivIcpkf2X2AyOIpa+ciMcdyLMnSd4Yee5J0yRGH2KTnvGTfAxLP
pgQlANfI3s3wBMk0PNSw4DIKBg12AjRVk4P762pU/x6V+9oUl6MHXXniMbjpMlKTzzslgjfsmL65
UcyX4lyBfvFID3nQOC3T5YMd1yai37eLom4Uk7FN5RnpXZe2i4ixyjzc/o0hOdd7ZOcUEujOdnc2
cEkG8GojNfhQuhjicxJJZrP8eOaN1TH020AbWiIb7BxAJ0CmX3DLxKgrnMj1cYHqwYhgjnjd7CEw
owBVWbWrq0bW9C9Dves6xLxVBBm6S/0c54gHsN2cShNPubwmDO23JuvPcmvZvWRxsoQ/b67GQ6jg
3MdOXW2vhdnz6Pdnp8XoozRhoMBOS+bOFagUoCnBPKVpXsoqN64E8vtqZhDo8TtCHX0LOytj79cw
GwPzgaMiz3IfSj/1hAXu/D8eyUz3oU5wrLYwghdQESc4YyrpJa+H93GYvpXEwVU1ZaGEq3s37eTU
b3Po0wORLVYPTEVHIRF4PAQMv6bbj6KCXO0r/oFRI/rglcSuRvClpIuh7fYzQQ8fQm5GRF64L3nS
CXKBVZYG4GFfTtXwGBPa8ytPZZ8PLkisQJWY0zSKIwaoP5sGpzNjzKVRoIm60s9vlhanhgK4Ivs6
jeZDubVNXvwuDf9xM+y2jlAN7Zb9/ZOPN4gLYes/F1SkU1yxARgHOqjAWVVGnqBLZFVI72VhB+yp
cC/KbVd9Uy4webv5/s8lw5fNTBgwifm5CYo5giNsy73K2oRHinXuDzavNftuG0SyrUMMooNxyndE
yKGOl93dtbmw1koOa5qM4tkbPfQEkSFmRCFJ02Jd2pH4YPuezyQvitLKBPquesNg5ASGJtJzr5Dv
2v6NkPVMBw6DMIil/vVBsPQ3ovbeD8KCWQgYxlMD9SUsUxTrw5lId3nmZ93u6/sBM1fmJA+KBUci
9jylzXZPsceGbFie/pOqf6Ja3795sHUEHS8l4GA+/ZTzu8frWrH7zQE+VtvmjbuRAd2zhWGweDYX
IJvh3AQwh1OHC6n6NqggrTKMbrV78/xD0aObZvKFWIGxjGA1bPrRzLCM6l0EPFy9LTcOC8pD1hT3
U4kFSVxGO1JAqOh6K8zes120kpE4sdidDM54Lcu+8eDioM5Cd4oLH+rf1yLueeK1qwCzrfiZSqOl
nX+SHG/06tU70s0y6PM4yfbFph+Vz2MBQDwDBUfM6bESpRbwiiuq+/g29KLmqcOq8jVuo/wRa2JB
ruGjcUBenBbDw8RyNIqxqwZuo3W+EAtETV5FIfxz78/4doOTijvYuPz1TEk8zVXcL2qP3k8G39x5
YVUXclXe3vqMWQwUZKy3xRHAASmma7Zm0+XC4A7lCuxNE8ZgS2O+31ges20+dYeKyK5TrgCv5NAc
Ifxe6SxN82YoRP7cXW3d6r/RLGpirrUIzyR5DG3RxaFZD1acrU9RJwQQREX8WWWzOM7uB3hbMU64
kY3fCJwamqH2V5JBIzjOfcyIUI1GaYlmZnSa8a16gR+Ye0C9re8UtlRRw0rMWFyx7vbw+QSpXads
xlujY6StyBOaz6wczwWmQTNHNPDXQqkNvtY2nIhGkqA8Ua01GLbGAX9yD9+q2VOcVkILrvwpnxZU
ezUYqhopDr+zj4EAWj+GQnMetAmg7jgEYO6p8ePbH7lxdWIUOa29PTEtRaanbVMEteCtk0klGd4p
AZ8dW973Ju9Nzww5zeUJ8jnlQ+1QNlMKi3mKfsFrXqm0tmAGL/g1RB8CSyUMVR6mdEriF6WP0/HO
11LWO1RE2WA71E1Lrbt96nBYommhF59hpx0tKpU7P8dmPtsiaEFTaBYab0WfhveTe6pZmd3dZSX8
8gB3rl4R2sw6sPkw4uoKpb++7P4BDiTl+90bewhzCl5575PjNqYzsgOAXcTgip1mqBHDpUP1k20t
r2q1UhAt+SxVzw/fuQQymEoxLWrC6xSo6l07wvr2gZHIpLAy+mZqBMPNXgZ/3gNpwoIvxk1uzRI1
nWJoUh4XgzLYSMzTUg32mMzdDAVlUchBHkFUYWhQCvAMiBh4SnwMtSINN569u5QuUutw0sauThh9
gWz5aO/FkY32qe/UyxPHP3tDVqgU7meBTaf800Mw6lWRhhG5mqKokGYKnGVtHdrOXtblT4U8oDyk
cmnAZtIau+wMdDdpDLsZzLXv1URQjhsp2joZoJWAaxtDCN2vr8cslG+h42tkoey6N8wrWt8n7x3X
QJh38bMnrfbfdnBTnBOCsQqas5eWXw1j5gad2kzuYcE3rEb2hJowsPAB0iMWdrUWhtLLEom9kFtQ
USxWVxkZwIAnTpskHNblqgnJCRuVwH/SpGCLnft8oA/FUp9JOzXvUbX3AN1PkWNma6F2RQ4N5du+
ZlpLywgdkpyQFZ6Xt+q1m4WkCIfG7y2W1WjwUfiuhRbRTa9T9H3jwplOGzYoBU/j6uSI4SdV/M89
V/hWVdVCwplcBnGrRSVmaEssCpRxbrQoCDS5izrJKXdwDHXtrndbXKFbdBkB05ud1bg3uNxoSBFo
lVAJQDFYsu19aCg9U7uiqvyzNDmqYDJ10KgDDXtCWk1TRy/6v6eeqHPYcAl1aZLR8t9+vfd2S0NB
wRqWNrG67IUfOW0AZ4THhmklStjvYAyMr0uSk6Nvzv225vUi9jDIBGgb5BaeqlvBIpl3Qbx1SIS3
W81doOrkcVzGPo/Vk8dLhGIyMEoMcn6zgQIUmwg3NJyMhghBrCUthzVPEtSHVlYh6NocWK1U+SQi
M++WvDxFzCr5gOAPPvSlx5pf4s36/MwihJSypo0wgd9roeVgcxKWFDTII9C+owcv+1RFcQTPU4kS
NrcfssWg7u9WLcRsdPkwv9jQgpSmpIulSK9h0l8vd8cX/PoqlV+7T8qPVcyheKuSmB0Zh5O8Cbkp
+hTMfUst9a9FF1dNN7eXd3rLVHMt0Vo9RzwK2mgwXndZwhsJcP3LL7AfBZDVxe5+LMOffrof3aJX
RpAakXbJNYCTV8zvLeuwjkAMRBSgPJBJq5FuxmvXQCGrvvlieGkNr1D4kUh29KgDzNhJRbaw1vof
aQv1KpHhmKTW2caWQiN07QJNnuNO8h39YrhOb9E4dlgSvZSc8qVs6VuNJEZpzJlaPatDNgssz8aM
bBwHG3K4b3jQh5g9b8+zPqllrZNK5q9Y3+HrDi8d28vbbpUVnxzHd1zEbp7E/26mUZRHIKivx9Of
YOlhwAw9zkFJ+m5ff5/8OvNMg+8ggocysYvfRpQzCXCWGlq1ggJIX7x/Vx+YyBdJfCMWNZvXZVMA
AU6hBjtha0OjSAq+6vSaM95PYtT/IOb+3ZUi5XI/TI4tdjpsogheCIU7OSD59v0C4XoxERn7DJp1
c6BloTa168Uf+bRh2uKb029ceH99ldUJTKqjKJd+MCzEZydd04l+zlZbC2v7ugona4PX42uQEaUJ
8XGpoxWq9xdD6kR96npTXlO0c2IysyojV4RG4czm1kJkinQDF+jnDklIgsNgowKLRyPOn6nDBCsb
Eb0QdPEj87aZfOSzgaGAYBf6QAqE81EuyeaXMBY9MEU6vjA1GJJ0q/dS7fBUDklzOcnzZNwy3Fot
T767D54wSzU7NcUSyQMdFKQV6IaMuzIJRaH9sGlBzGuNoqMGNyO6YlBVhj2f9YAViNO0nZQJc6qQ
HEZHNKbMNc0SNvCEyXrIo/mJe1ws3Vll6gj3RaFcGxId7eGtNOo7s1jBob0gEwF/LpnI1oltnkm7
j+4j5svlM82s4HRtdrdlcX7G//mMIX02rKmytunQOUlrbsI9N5bU06dIuojOx+m6eepDTdEEN9Vi
DpHKfqL+UAqo+aEdZ0GUX+u+9ZD4kxxe8OGt8oHZenxZX04xAqgA2qvxF5/c/1OiUajUKjB5jWNn
eP0ukT0LGrZCE408C8C2xgJ00W/myyNJGiP1vV0jwVTXB1VQmf8/VVjqcH8On3Wfg9EqFKF//59e
m7lqIb1Cqgkg0nZj/wbgz0SWPbSfy+JewI6GkP01BJRdc/YvZNWaSQKtzY9/xQvqdzXtrhuG0LFG
z0iAzeGaERmpRRBKqYwCPdaMbakbBMdeLr0pkeEeT+EApF670At7CAb/GXK9enCJmZLPhVe2ytN2
1//dSknBhBbKhzaiXAYCatJkcUO3kqyyvbDwL+kka9z3lfWvFSt/7tU+lOeCFwWPL+Gu7FX7IzLI
VAjWwCwabM1ABrfI0FxJlsU65SsIAAvg3XP+HeoZLRJH05bama6ymOemI0fRjzW/b991J2a4PYfq
0iB9EmxYQMepeghWSp4s/kfOWd4lNh9ncObFv++t8/3iAz9pMHDxbRFgqdtp0C2GwV7eZRaixy9L
7JIRcidtlPL/PyhubXeQ6qf+sU9Pe01ntjUtPluA6Bl+EVvA6pNHk81JHsDbVn5E0fZvfjife/Dl
7gGCBTVocIsuw0poBCOu158YsBHZFedcixXNFrv2oSEf0yLzK0MMJ1Vat5qge2l8iIWdypHCIyRE
EF2AHtWdMgZI7i+mlLFaKRmyadJrwvl51tIklZacAb78wCxEvYbXq1F3vEe765WMhsM0JCVOy3by
cRNaMNMthcEyyYImX2JGiQEiBAdJvPn8gtIO8NQa45Xftwr2Y/2lQLY7tUQZNRhmjlhBdEgRc2Eg
vc4Md7OeomchkNcDJZuJwtIsgDleR5rR2+YudHCUWrzqhZkB8PdBLcfSmAlNnn9aIwYjrZJ86m8j
5isAgFN/G/KftzWuhzE63O6R7pMIbUG0fAKBBnEu1iVKpb4UUZLqjJJA88hz1+pXlcW6t6lgnooP
ytozO50KZBJ5py3d1132oo2GfZw+j1z/94cV08HwCbZi1ukIdyUfv+z7kXraII/JQyhTs75rE+8S
AKUcSf1CpV0u+Q1yIdjJmfZFy9RQ+KTPzH936cux8Oz19MSec2owgFnhcbI8Snhsy9HFGMlOq6Ca
pk5NvKctffgywXenJ5Ua7IssVelRQIQ8uWKjZPfT6i9458h/zskmt4w+3XNqYSB5bqKVhzlUi+E2
Fs6BnAbvejRKMB8Lrxl40553HHxIru/uAhcyPfMPUE8RZ75XmxQnNY9wEqAQsem8fJbS6BcIRLtd
nBq0KFbmlcTddL/46R8IpDRUfp5tqF+ZJ8tLacJpSh9I8YsaKTfIKYj6aq+BX611mfGO1oI0sSi+
qtjz1SCSB3fthB35ndRoietNEkkTjKJy5fItiaAY7jfw7SFR+G+CDqU0uDIIAG3reb6qSVC+6rjX
XX1zLbaCKfVk70NilHwfA3xci1N1kU7WEUp9lDXJ/YWrVxfrWq9Hm/t6LiYIMh09+yZ8J7XwQ9iT
gdUtyJ1JSnX4mNxzX8Kk5hO6KTwOJh1lT6e4gUMVhVevcZJRRPluYvZdHaxaykJzVTNQQN8Qicxc
dyww5pmc9Ucb4Iqxv/XQeufAgVqtLA30jQfzglaZqiry3bqfjc8lOUAvtIX7IwHLniSwgpkt0+9+
7+9wQnumzLIGjr02YOyeDWiWbgOG2F1X4PEHqdN+B9bvduUmy5IdWbfp1xb0o2KfAKun7Pr12bGk
pgPri+eOjd+sb0y8U+QQZshk58YjvwjcNJ6bkfDqrnagnIiFXhLjVf0EOwG014ldfo9G9dt8sctN
B9McqL2tl0XfTRevQ8ZUyAIw3NBF3kCkGJcFnmrfo0/mN1aSXcXR3TLCyxNDwwanm+QKQYTcaF8w
Ex5jtNGhxW9g5hNwMYN6U1nj2BG8rMj1ec8BeXAUVUTg1QtQCUOaOfW0aYc6KYOqGV71Wmcxn9dJ
ryzkcn7KcuRuf6Y4HLjW1J30704gKBUHOUnDs1JGkABaNS9kmCf3UL8IeMzWTalUTdfSpzSHN4qu
N5qdpIp1EB1SGtLPWyF9DQA/IYqXJnJx2ObeczJdBBSXUz1jR0RBoL3JUJiGnCHxDlL3quxgLxup
9th75r/OE67qRvuziNNVcWofeWf3m6PCFtGnd90Euh+MK1eHM7yGai1m3mq25RaUnwp6/s/Y9WB9
veVTr/3+RMS7HadepLDvyKxE0BlICv3hpuXFBD/wEU6vQ0Blf9uzQkBMuCxzommowr8YD38ySzvI
d0rWeX3PSDFL7EWuNy4oXzX0dPhfgwN/W3m1n+OkY9Ewknd6HVkxiW31qlay3FPzjywb9wXWqmnm
4CnICrD++YNjjGe4nn/mXk9l2gY8XrR5XPIFgj3ixd1Pgsx1ZA8423kKBBcj4ft3GnSwW6Fe3vDN
mx2p0iY6j/3SeRZrtEplU3q019z2IQ1Q2D9B+qFGph4UQTdy2K2KDHn6vVSlLRcnH9BMkTLv/Bzr
k5TbwCU77D+WtEsqPBmgsq7HmcyT8Uu9kRbl+oXg1OT6fwfNO6AAIMXBCY2P5dLffaf4BWCSyumP
uyTDCwaNPEYbNBq2BxsF5eQpoBG6lXQfkVXv8VqiHF87X7/M91heOkJE4mIlBqQJ2zhtnkYzMBri
1CIO5Go7OnRiI9OGpeAWRv17w7niEikBwYmD31JHyMb8vR8V4qLWG499hkIDn5EkbNrfwkdxAyxK
Wd6AEBH+xtKq4Qq0jm8nwBTKZWwBahfRDSwZ7JoA5nH1m20vUIAGacwjYqqtc3wegziHIpLOAIzN
pBqoxpVGiJfaudq/3CyRZ294Disw99akrk/5HEz/x45R/Sa9SlGVBzaY2Ntn3DnStXBqjVDYKxth
qjMpVvM+aWmdthBcl9z0vIKRRwscaRKhEvkBC43L0/yvxd+6jQqXGLDAS4AmUTdPFI5iDAh2qpgp
RyEb1qkq7ZEmfKY5kOOGFeCt8vOv9F6eQ1w24Owdrox4vNyuQr2x6+0amcyG/D1kXGtyJ4QkTgbO
POIkRZ2pk8b/1RUN3gqutmShxXEDrmRgbZHYdGfokSm06hiRE9QQY5NNadWTPhVoYeQV8Gq02wYz
mx09tJIm7c/A7r9Z1W9Ogm7b6lrL+T5i6NDJxzGcsWSatOSqjZ46ySuLuJ8V6vAx9wvvqIIedzgm
b76TgidCoemYkq81liZCrETK4kKLWDeD7uID+826eQDj768G44Iw4+EM/dH6sEm4CSTMTaKwJdXm
e/srlUkVAfInEQ2/Yg7KkIEF6tI5X7pp4JhnIEoUC2/n7gNtlRhbpNNANJ0RJxdfZrANWlUz2dTG
8oP3owoolESRCX7zmKrolcYKwczt6jOjRVmc6W/X3hhSmIrUqmtp1Hm/ckpIogD6DHbKIP83UarV
eqVRHyrwPl25DW64MSJB6p+/FB79HvbE75r0W+gAfpjzZuLfU49Khul8EZwA4hFrEOBr0C/B8lS+
zCtPmORkm79FQVIfwewpI8Hy2rk3O62URQgFkV0grXdZCOn2FSiOWf3xh/K5TQ6afuDWNpBYt5mv
zMfz2Rp8YX/72pH/a/azhBqoAALqEpQCjIADLPILKO1rHYj9Bm2y9nsmlYMECou3FvHViqn0U6K8
QpTlR1NfB+eAp0l7r6hlySMstpf/KdNz3FdM8pK9ftbjFfU1lquw4SwU7bbjbhUgj62q5GbJ9i8L
Yr+X5h8rn454/KDYu2/KEcVGOgI3uVOJrY6kmg/nlLF4mAkyWV4XeMUNR4mj2aBFtegrOqQNDJc5
jpFMFZjNFxuVujtemjiHitlkWZ2tKrjpTTYCY46NZcnORsUl1rvoHaASMc6cte6igh4VTbBsbePT
EoFX1xx0v88jTAUo49u5mUBOSyySdWxMkIeP59/Krv8cIt6YDNskUoG0UK9xtjA1Wegx4okJYT0i
IdHKKwcFobmP+tvtsTuXDTS7PtOR3CY1yGSbNOABHCdJF3baEtU+VthDXJlBpZWTa7XCsPgr+AOp
+V7rvAf1RYF83sLaD+KrFbYXSe7jfB1oTkETSeUj6PSC3x8vh0G9pVP7CpX2YaLwT1dbpHbsPlIP
1hdwJIZzwhhI9d0+c1O1C9/Ol1Gl3yPPO0jlDEqdCNKyMlXzPSx8+xri0d4cpY0C7nMN2XKVsEM+
4Bj1CZH3tfNg8klNrzFqyDwQh3aV9u/Ly+ZwPz8v4GkwCcgX3p/CTLVcEvK3qoy80KDb1HOUsFkO
e5i9mBIICpucxf8OdwYJSmO4ABr58ZZLYiYLF36jKvbdjOgPL4biOh0CkRjFrbjTR1w22XvcdWyI
jqqoMdh9bYFOq6vWD9hEOab5PeqOfh8QcgOgZ5zNDlGuHJY9ATE8skEwAZOTJ4JyqfszsVBdQLY7
zB8bUOa+2F0/HWtNOtUIpa3v4g7OctGMKTVmlLzoE81lFVkMRXyKjfgNu/wVI1bbYXrkzJokeI6a
K8f67iS+2O6BT6naryY5lSA+vorJO7miZ11jGhQDyNCKcUVho6ndJnLZcvVpZ7rgJtQR945OK2gE
S1H7ZJ0V2ZZfzPFDFGf+GKGK135cZ9fS+GJ/aZiqwG1yKVoep/0KFRtDJQvQAWYwT2dD9QTPxZi2
6qFPwU01C9p/YctVUi7vXz8+Mq4pthrnbuXt5gmHsCGIlxfHN5W3SWCxvTtLY62A6s/xWPS0mHnH
nbwDc5qkTzQVxBG39F3cOdYIZn9G1aHY72MU1XuOVg1tqDhDvNuJCAAnMTNWv+2Nb7qnsWXruDYQ
GP49ooz3ZR+LX/4pBEWgN7+o84RjYVrVgLGlVx3qkQAqIoxn1T6UwBUew9jCyqIDtwS+cAxZ+4YN
AenD7xAB43hq8I9gVu6iyInFRwoDpcG/aka37pVZH6sfiJBcRlWXy/4OL8Jq2Q1Ia4Ry7joV+PyJ
wZZfQmSfxtIzgIHu2uZM4XMxzAmR1MdBfkdE+a2Jx6Aqc4xXyEdgxIlPbEnTtIzaI828fFzpz4s7
ntuwh+8p+2aKQKn2kxtY5Lk1Ed28BTjLrAQ5a9nDjwBZu9TEK8+M1kUj3/R2DfD1vhPzaQ4aZl91
R/tMVkJ0wGCvuAi88x+KjQ/Aw+HC6SkR1m5ddiRhpvQWmDK0gmtNz7fBJY7MFmYCp8RBLsMPrGxr
42mAJeScCEDr2P/Rm31j7SZuuIf7paRsTWqs4oWZ39xBdyYLGahr8kehngux0jcUHBJZbE338z37
GFu/xD1jq3bH4TYTtaNw0I7JpAFyUOrVJ2Y+DPsqWUsVmpGZjFrp9Y9mda/ktfQMAJnNrlcnB9gN
B1ZfrO4QtjswoxJ36AZCSNl3MOyMEoTV/TDdUTu/n9zA9oiuc1hgTUiwdJqhT5+hDqVUYq46krz5
6StGjcqurIWQwgOpgyEq9fiIr44uqCurA7YWHWBkvpvuivI8jYvs0J7+oGK7sjvW5CynT/Sk08Tp
/qGM2OWfMh9FkTdmThEF4qTPHJwvqt9+jF3vReA+FEtFBcrPpuw28T2X8ejg16syuhtsnfvxC/Cl
3AYGggP/jNUPCvcu8m//mUBlwLwoiz44lD8FuDPhLj3yU03WL31g277bhoGkF5oThFl+wRvRYIJf
XYEOFGWlBxzK2YrTKZWGlEt8AEc2TWil45oJziSuMhsq9lTJHZQSTSjwT6yukMW1OfyoR73rhsOp
jsW7vstUQLIuRNm3qNuBAL8Zb2lwshcrgKyrcVLUU22G4TiMmqgHX7CaAl6YazJZ9dOq13DMHJ3I
Tlm6Uj1FOUSm+Ya2rrsdsGtJBImKpk+A5sZ4ferBKcxYztdKDbSh5Sumw6utlX9w0rhZHuDIin0j
w408ucsURkm341Vj1yE/QEu3VaRvon4nsi6YgvIFKdJf13LN3VZYlIP9h1sorJ1UxBgImBrHOEgG
Lh/y//imPOrVCRQiyxMYDuFSJfnHoC8k2+0pOsSxBP2rqFwx3ZfaodGUapzs+3flROzzgGDthW3u
L4Cvq/br132XX8GA+OrmhRax3FGcjR4kQfGZ594NR9iCnx+3MjUEWSji5880tVJWEG4J83uL1yL3
B1ie65zRyBPUbPq+k8/qar5DgW/y4PL1fhYba9c3euwr4s0Id7OxPzfGbMS2jDoCANDYPBn5ts1k
ayxaHwm3anPu7Oszmrqt56UTNDZhD1dcsl8Ax2MVWnuyhz//s5W4fT3etAMLuEojTaym3C0Xl3yh
Dyojlikdqb4PIWRCjCc1tKiMO7cDCinkMUsFI3zvA85Dy99yR5Of5/IARQOMHRF2zb9kuYQpNuRn
DgkAq98NFHyaCwHm1arc7sf6QCHVYZGL4HDOL/0qsL0zgI4hryg94PV3TW6zmBVlbtGgLeOyL2pu
DfBLqSPEJLqupXSzdNHNEC6wY9xOL+7wwg/Ps7c9mSFj9dqnmmwoP2Ljw60ooA//3LTePQHAPCn9
XIMzHsoVQGAGy+qUiqDC0K3iq3NGKT3SAy8TVjVaeV6CT++vbakPBW7hp38DJMTEpmN5fAycQFNa
P09BYflF4Jb4JIsEbZ1GT1+gHIzlIsOUlia6Im7Yc2Z5m414+Df/ehX1AaDKKK56SKYgYwuMwfeS
7aULaKrr9lHxGJr5tO87whhutcUKHe5F3i4ts2dsJZg77F3nvI7TH3vIU9YhAPzOG9g5TmtePXFB
0iwbBRgZQUahBvEPyja5NCLfAs2Qg77EPdcZWhmVYI+zbwIrHc8SHARubySfZpMryNOZGjhImubG
4OJyhRrzpMvtaYSU2KvevxaWVS1XcFpFpG+xyQ7op4RCtfxgtvRMRz3x3hil9SkZW6P9Bjsc2AXw
N+Rf5qkYevVK4m3WV5SYLiRIl8C6ty+sNlXf7sfUbPJLL8aBun2ae/E7ywcSTiMdBRxlPuRRpKGe
3NIekQ+gpdkN0xOG3tmXbijyycP+OVIMgBDbQdgRmNfBkt4TB7tHOqwCWwgHnMA0VjuYJ0bEAAzG
75vG3oBx74vSORU0tBQJqS/d4ZEY3CwTI2PhHEEmIv9Lxusq0tkzOO8YBqrs4LKOW+KNrmJAv7ZX
YmNDlMDhyKB5jarUDm+wTueUPuyb3Bk6aMFpLgx72JIb58tj01mWJLieQQMWpPvlHuoPmTwVR+Zm
aOPHCwenjrsCb9ZXBDDbss/kbowmmHxsk6aL4Q7jnzMKNk9UFu5Y1QWHsV2yoa7uMRADs3P8zAqP
Zje1xXu2G9G+JMWjnNAk6Vvv2u0pkkQ2bgDvwn4b8MsDVOCMdrtjgU1qTY/2oUq0/QJlHN7K+nMb
ew9B98yyJ1dCmgGrfBuBrpg7df8VLUMBMO5AOb/LG+GTWbb99GBiPmgUqmJDQyOFqdcjUKuQWea8
rEuwystFFF5Hon4FAaTnaL644OIUr+FUDvUmC8Kbg89TsExGdn1aJjc/Psn6GIuoqEnFvKJt5q1R
p8wiHv2acmbH//ISB1X1hwQ7/pHmPM8fxEHWAptK2nP/UMDJy2BqOeZUSq81EsQzy1kVFroNyaks
ut00sd0OYieeXlAy8EK3JZnxlqQut3dBcnlbhSlpFAD+XDn2RCrlL1pdP20xoA0kwqk/bSwNpXmm
+tJFADu6mjRhdTVrBhOaEIxKCoTRfsR5gEE0kArWgUndC+/T1ay3cz7PJSHPgWKjfDAwiTQgrumM
5QrAGuCitPAMGn/HAqJZjqf6OLwby40DPowNUWQhnNc9H71U3ZIIoEwqLW3dYL03b9dL5acmNf9c
KC+yw3r6rNQujWOxPbBvO8Ue1ki3nfFuNH1mce7Z5y9kdYqqbVp+0bcBy0G6Fc5KqF5y5ye0MjN8
sXGFDbehV/2+udRtTbEP2nF9uV3ItldiSZbgYug95XGnm246CHLnEc57zAE0P3GHakWEeFlIj2BW
vxWH0dM4yPeSnfO1xFVGbP4HNFqsCRVXMV9ZCyNe8ZTMeo7jBcRtF26/K3e27cu4GGKzkilWee+/
hRuYWCKv2avNqtXDtL4w0eDLyWTO/Gqff2JykPqf/rW9snSuXmEQ7rr/mCtf2HpRY61EAI3vKeQA
xhJhZ3sbct40XJxPAOq2K3qYxXLysInTowtGfpbofZOQRhR3Adj4uyKmvEFCWFMVrZj56mxmOJds
G3CapILWdWu783h4vj8IgUiz0E9n6Z41nZHQhlfVejCDM08B8iAPRHcy7FOsNWPaE7YiBG48AD5a
1lOgvIeS9JePYneZeNsue083waXC/Y9fn9qlxmrtacJXZfJ93ZmxCsIn8WKT4zEPCYv5JJtV+i+L
yblXGOJBStCr2RdbbEtZ9bhVNVjcMJb4yUBkqN/PMWFIXs2vsKg5fDotvNZaORS4jjyPFBVwjPsd
IaRSJ1Zq8tR5sI3T/CYyJU7fBbRT62Jr6LnIqu6eXg21UQO8AijplCtOxEjoiByOzH+I+I5mL+Jc
pKu8P9uYGIGly6R8qoxaRS92xCRCIh8VukNgTiszYyXPlyk9ayjRk5u32opr0d53Diz4ecmV05Z5
ZYgDOrQ3UiQAZUSK/t9KLXjIscB3oq09f7uypD2rpMugoX+Y41Jn9KsfN+KPHNrlTsCvZDhEEsqr
w0gdY3NrhaQUUzZV+omkBtnm34dTyhaA8jKjV1t1HbNTVV75JnIKDFD4kvdaQi0WZmsRuHjFmkNM
PYmM/JEf+2zszC6ofANyCQ/ZBIAWBrA8b6DqFfp35/5F+VUo2jWX8IBFNz8oOhpbTJTzams9mcWC
K+82Jr9UueeUuVnXkSjieUC0dE6jk5D3BfqrB+90HdP58ZSC8D/h6UWwnRfJgGS6vXMkXKJAGIrY
tAvFg1G1MCOZYyRAXjot9rpwqxV/JJvrDG4NQAbQkcZccuNKm7TyAgBc77QscYQ47u7Qt0d6Pdnc
k6HURUodvOFSqcBYAseMiEQ6xA565rJB1C5FOAkpBg3ngV5+f++/owkzOs8F6+29KMIOeTAVs7EW
rDjeJ3DnzdIgCAuK2T1IPh596F2271YFFmnkcR58Ar/IBsYT7gifYNhOeaN2apKxZlAtTa8bb9WU
//blmuGi72MPjxaUtZYWzeuzC/0qpnenIw4jR0vQEVgSWItZ+vHRNHs5b8HRIjOboumMJ9+2HdOP
37xvTBtlcuPEqmrVveY11hRqvYQ3AodwaRWEMugVVWb+VbWf4hZ7AD9xWWSzgCD0hWbYZNwxd3Go
tP3TwCN7WOh+U7Iszo/euSWZW2sjMu6UUq3/HKJUfet1yih4+ADMyKdY9pu5pWjhEszUcwpTIZ6W
GsmCmcxWL12+Oca5B0VIRF3ffE6pnR+3Miz7t7A23vF+hzwZclf9TjcEb7Y3eJiCyh7n22uJAkwf
5/fVKSmR9S1IZ6U3Tgq52yvZwmRiQtw1Al+yUiZXUhyJJNM6w+jU81RCFcxz+vjToFvHF2L0aq9F
6sqSlzq+TEJZukLZtqhsYvesqC7oH7vOSirYgu6Jz6r//iIjWoL2xXEFTthBLontUDlJYQXF9iqM
1YXs4hUnAI7JnX5R3gjeZNCez2NN0q5e5mB2RzywfPesg/Al1cUh8esZm5rr0b7BzX1+XvQQr/Wp
ATC8Q3RFURWO1rEVN47BkEhDre1tYRbGW4ymdiHE74MbsymVbV8gJP8rp44sARUu3eMf/5dYWYF2
n3vq65WqxtD9PVsxvmEv3mryBF81pjco4xialQJf56DVArLIA6K72WJ9nbfDS9/Pe5dVA9Wq6bYL
v7CYg8En7mgdhviglhS+EUWoCJs43h7K8WMfMoUXwAgFvpH1ui3te5rNUgzviguswe2EBOcSP0q+
zngzdRR6LpYz/FUyUI68eKvb1/7kc5iu3aR4BQjiWUHDqCM0N9tcdRGkgk/QjzX3LJ/X0qzMWk6P
LCnvt1RfmNsmrMojMqE/O77Q4zR5RpaTtmMDw/CvvUMY1iPtMoscJhTMgZY1V49GLP3/TmmMU9Q/
aS79twFHHs7kYFd77slRSgQUVI+hohx0Yfe6kVbzApHiittACeYTjq98w9ZyjVciRwlavXlDHKxm
l8Zo2oF3npOnwjyLz8e58/Hpyk8osTzlLOLe5DOiN+lNWxtBPXwmrMnFMupyB4NsC6WPrKu5KElG
iyrMXl0cFfFS9BnBrQdPkSu/tL47cxi7dNr59wqSyGPfkSyUvrLSC2E5kswWPDcVhsXleEtQ0+2V
JU0nsnaBhtT617jDMaRk6yWdWrEKGl1dJwH9U0NK0tnttOJ9TsL2VlajzrIajFryAwtoimRUW6U6
K9CvWvFklLpVJMg7kdCiKSbX9SFnO3XuxI6bsnW+vWvFmcEY13KRHBVjHoKraxLcHaVHJpgTnQ+L
Gni3OpeSBxhXX/GJaijUgnt3xSRpb3OmVAxpZZJvfiVvdYtr0ZaIRvaCpthQX4d7GBTwlNZc64oH
kUV7MfqpBV20wFfoDa+z7dwstPAgQPtQd1PzlU6iOYRdeiksb+DoCCmgbk3PfS817Yx7Mf6CyTZQ
B+sOHZx39VArXnaZiMby7lIlUA7cJlRwwqr6gpoC7aGB3u0M7d2W9fBDqDHKvn4eF20mmVQg7o68
ICBpuyIa/4s3e57JotgeP4bsHMusRvAMV4CsD9HKCY6pD2LB3rtIwfOf1oRTfTw/l4KQXNc6kmji
dI6MhqiuyPskYV9/pYB1w6orEprRapLWX7wC+dbCnmXSREtOtj/LA88rq3fQ3Iu+zMX69cT8/xfF
S3h1egp7/6FwrI3rlBrLmezNnOPm6gy+ZLbnIMDJnArZpwddftyV+RhX9gSqdO/2aB8MyF2WoarF
KzqaiOrzzNEWzoPBiR/khM52eAT5DZABeOrs3Fv4N2+qYxCKnhli9qJB0IIKi4xdzE/x0KvHhOpY
Q91SvBoUI6DVFomUc4kE/6ddKa+kN0L1quDZQDAn3i0ACHrKDIZ8zxRZixEqv9/yRPpiSaM7R8E7
jGPvMGJ6XzyZYHdOCLv3k1dTdjNCH1RXF2gjsEOD1BMXqqTgPbLUj+0k/GrDGmyZoW9MqPKQ7EQi
Sw9ojOyrYgvvgKaKaZxVEvEKZNqb9hVfVSOhLxZrg+8D5HYAAp9g7JfUN4Wb9K2l4FtbFRZC6sfK
X3oxLNo7hNsrFcllPmdqKbPBkkzvoiahNRGjEzwr1nvnA5hmnasSMDOFPGv6NsTdXZA/GS6unw06
/S5JTDgX1LCCkaKfZn+FMPeRJ1D0QLZk1xm+FQpYlAuwmfdzE6DAbxvyg40NTC5MfR+gXEiwZ92B
f556Ys99VhYMHnXZYlXekh6gPg0JXZtCIWlKQY+gJErNguy0TJghRbhoI4esecBbM4C3PB8nNe9X
sJrWhow+BYu514R7q9BqHG3bKEnQMchOE8mlhyXvRwbUcu7NT2WtnYkt1iE2pIdRw0dlCMslUl5c
QbC2XLBszaUaMItPOhXHD+iaejqMrwTsnMktz4WsxR14G6rP9jIZdLJDlrrQv7HGLJRkOh09sRPS
4SveNhXxNQHNg8AMvy1j4tuJ7ggDtr1d22F5QMopwJKec3FuIIyS+KBLiJHJAib+wVxFnZBbzAf7
d4SzHuGNEMHbpJF176gYIRYWnvGdfL8J608NIxr6M1qJ7ykl7efTpucX1TkEsO3fFvSbnbTW7Ayh
Ioov2qYf6xMcogcosoa2EHeDYdvCsHPrgKDOWUeiwJk85RSL7hD08/v0ejZZ2uOUL3HrYilHmvmf
JdloV4nXGzAPhwanlv3GABHh0d9u0VEOedGSkWDV0aHTU5zZ8tYYTjKiKTgKNG11RKnGUoc2vwKl
DnaOb3tFF4zL/3Nm9tCzhBkQbUnDT58dTp4m8iiwk0QKi8/q3VgqP8DXP0mSAFWTgvAAmtIYW6iy
B1LiD6f69/OMM5ZFCMF6g0aIzqWYONvVm2pRHPSEujj72NuvC0OHw5t2btCiF1Og5L5w3u9HqOEq
nWxDNvs2DFJyMk+LehdixxgVGOZSZr9jb9vlgISa2Oaw+JYzGKafbwZDnePIMG75Yegt2zzpUOPa
weJRKEDDENTnMG/VTsz8dLtlMtB43rXu9Gl7dIBpfSTdhErjV6yq8UGiWx5QxvJbzUYVHTol6OK+
Iu8yeA2lz+FRUYHRBbffOczjDFWgE8HBkz2wqFcRvS/XFNP90DIlMaZpVvoqUMBMFwPvWoG1nDMr
o7F8xUHyMjqgbuWoWQPSewp0DEXL8KRK7znoRZzJUZWGzrlDEfEGpj+bL+L0euUsgB4FSKIh+jd4
44HkMBWhDjzstCSgZfMVZsHMGZunGT/2E4doWcJ01QtzQcfFsTrQBr9hD/flJ0QgSQkgpQBIsit9
+ddeU/77Uhw7JUqlz+ZfqWc5lLH/uhUs3RUs3uPrOGOGerzvfxZ6gIFBDnri+alK55WqY2T0meog
RkgqfZWg89kUC1DyXfzCIFStWqz66F/W93PK2daKe6fIGjHL+BeiUnACUxVEiQ7SBwPI98OLPb2m
vYdKhLxbydLaE8VCSqf6NGAGPhpUr3U+fI7gsiR97Xa3vD5oFRwDYq/jNdNEYx3VTvDs0m8fo+fZ
qdu6Hm+AskIqu7t7vczVoup24pSA2uUUdS+FJnGD9u3ddsw06eyeFn+WJT9903ieqZUUBEpZcgk4
g0F/yiNjeJlIUt61bh8QPsExwOn0Z8C5k6tLMi9TG2KZiejuwGmxIaj5UW9hUVd7wAO3Uwg2c6Qo
qEVtOYBusnVWmg2TRS/GtEJhlVuJKeAWYGhj7N9N+wS4RevMRf78lxa1dmNsmjbdnOd6nMOrw4k2
BIyHaw73otsySBoDzU9AtOA/lIrLvFdzd9MQz1ENTBQ23o5I8GBWvpd1iZ9iu7Aon0Cpkx9HEYsB
4Ze4XoLTKNKrwuIyBuQVr69ntG5WlW26h+DjsdfC2hIc5kZqFH1aKy90dpTPkhNhrkz9Ed8PtVzi
lJxTNNglvFg1dGkY0draMLPNpAv0UhjmQ/0Ts8FHlxGiJWBZl+9Z30ZPeXeXZNbRcXUlCbt9flRJ
w3945c62+ZmkFBoaeAhOgAvkIpYZiGBiIlVi6hQ/Km0vB0/JiWxGbCtX3INh8+Eq6sLkOZK/YMKH
lhiv7I6+3KJnmQgvTjdoCQC+24qRhOyoLYwAeKdBPEOl5APJV6LHtA0XFIOuICHhUYYPuq/Ei0A9
cBCf2FqSAJDgEW31Jtca3aogX59hIEE/5rF+//VPYTIEAG+gFlmiIE4HO9rVFdX7R+5AmjDjtsIl
/EARKatzy/ZUbu76okKxT1wO+laoRKqrXWx/jhsbUdQ5FyVNLpMibH8RCDpXs5/IaTRbs/fsYvCg
rCRZpQAQOKemckXY5rzTSDJc+uPLQMF5FrLLpm0edwyRqRN+PEWcB3+ml/x2iSl7sLdILyOXAbF/
fD8iYveN70l4YZH1JSmiZ94L8/ujN9n9kcsIfCLNewQy4Z1a2/TCMjjhSNMJEo/rIXz10YFDYVp9
zR265k17HhrQgOMej0IKYJ800BCBpnySLPIllKC6w23kI4AAVgigvsZs/JCU2CTAQXfkaMEJJpMH
jjQjbRdzjlvZf5FCZv2RR5zdxm8ClP4x/CGXevp/UOCKoahWE8LNqhR8JBoQHlMVJGXnvy+BRkwY
/UFVHyKsTHtkeZLRUnyiFUW1XS+kcsOF/yYsQMoBKYECw0CY6CIqf40wpPyH//F1JVJNsgQ+ZNOL
FRofNDRgh72P7m3L3hTQlM23Q7SCA3e+W32QvJLxpjrC9i8fxfqyp36h5wuoKKLKNBc9INd0md99
HhH6kXriXbTQjzgoSgaYvmAJJBhpQoDb2RQCSTA12B2Tg4TB3szIn32As4V4nLwRMeQS2shKltkA
9WgHiPsMV8k6sRaQcLbmiIcpeeisGiL5f+Ym19RaJLUKFFzpW7UOFQncb/ZnbZ8FpbfUoyojEffR
bOy8eFTVbseWarIJoXyh8tzWTfq8McPacAyDRS40cMsE0aELUU7rKXDwFRep+kbVxVcWL42XzsGh
F7RWYfOKdGbTP0JqXkuW5SoeZJxmpG4l29xiV8GP/fPA4aw4lLSiAwmIYZGIo02IskYIf7Ti2A7+
+XLq6mlnlecGlAh9ndc4aVA29Ld5BSfjcXRsM4VzWJJ/PiI81up19DuIbVFIXBddMYw6DCOKX31i
4kVkwf7Q3Q74X7e+1FzY6bUFVUm3upN2Vmm4YmXS39whAaaG6jDUltFgypOc3DsSnkIk+vHWpl0H
yRjwujS9HE0zJs6N/FTxWDHQ7gsorwIEfEyozfdBVx1D4khIxt57UTUSNNcvCi0KfQdOjTEqt6Qc
NVxjP/PBe8Md6VQg+kYUxcB6aRAAAhFLQZFtFbTWhmyHetRPBGZPTRcqdXHsKy4B2eb5umoQse02
X/8JgKFfx9EHpOI5xRjzSF2xpeQ/kGXfRtTelQtg7GnsQwxKys37jvhsQZiBvueg+DBC1QHyXCju
a2TkO+Xqs1dkmmj9D5TLHPojiNHpn2GMCZCzVRKApw7N3p3luMSBgZNyyIdU1Zj/yLzN6foJ3IB2
As7ljhZcLRzfS3U+rYjf7kHiCHAkjl4zLg0XDk5VJNH10uvdsEtPWQ1K7lIss8NoJzxZpYQnNJ8r
K14gokX/Ha/WsMVAU01wC2cXerxYXTF64WLY3kRZUS/0Afz36sKdR4gu9N8Sip15+unKysGQt25O
lxaHqsJLzW9qjnbIrJNSagZ+8QRAIUew1HG8gLLzwtUNglfjs7HyqBKiMr+zFpKf+o5SKUHjjnMN
QuRnbeatD2yMCcFt0GAMi4oUH2uPayncWHT5z7XpDWrJOwadzQvpvoKd93sqMMftCgNMFUV6b2r2
jnxLR7AAp/9qvKCJn+H2zjMGJipAB/3MgCiIt2oPf5vGRo6+A3NtFBNJSPLM+sEd0uBY2IVnJAIy
zMiokz56i07SXarMwGK+ZyCv6Y/blLjR3yW9MYJudSl16DjWg3Xs6+4gkGmJdkNqB9+yYdCj7hu5
Id8D44uyiNgIN/bYGlop0A/qaXFWSvN09Cw5ct7ai8mZJxDdu0WBTb5noPQuCBnlpu88bK7EkIAH
2WUtcpjQ5/L597y1/cjDJQSNRNwziWh/JZepk2sXz3IJcaS7Yx2yqjFsYFNyOgAZneGVhMazhqiZ
tUKX7EBqp4wA/gzQL3iM8MCNHtPfCa7om1MPpomAn3k2fdvREnd2V0pfig1AF/cal1Mm23nDuijK
2erVJ/Z/LDZB6cS3cVU6P0tYfPWsz33qjBkHZhtRH8ptMzeu7uJVopJczPXlhzcZMSM9p8MQszkf
vHh71fIePAzSGpy3baHtI/xh4zmw3Usdb9Pf49i+QvUMr1jZxBnPK7bFLlMSbsu3jcgWcWx+WSep
dkK4lpHtHA9mUBAb5hpth60T7XT7O830fb4Bqkk9RCE7XmJCnLh4NoOG+ctKb2ERyoRzmopbWk4F
4JtFbQNyHQ3j65JVM9CE9ST7ra6d2RDxOs/tkeQhp1bZ3DTPyDdK3rXuAe7GZUnxL9SADe8Q8Z5/
ghXTmpi4AiAQf8jqyYDoZvlTk7qFaMeV5BBDMfvX9deh+0zVmGGH40lKlDzJ5pyt6CkQ8vWzW1+p
uCe5F1CDVkFqM8+0B/NamKkePmONbd9o9hSxXIKWEfwOdHKxxEBfT9X2ULU/RaoBBOuFSIHcAZg7
JRDt623htYG8xllXYNnPeE+T6aYzKvnppMfeSTkw2G9UMOszwFTu5daWJ1hT5ZYaKXWPWXyaT1/A
6E5jKaKMeVwTO77rwf79pn2tSiAVXljvijZYDMxLH4uvcFwCWIy41pSHrdDURLJF7h29PyCDPKE2
JOQl7q64eeZ7evYMmkugLP46tXjKvzW0t1dsgg2TWVnNr9FL3XGt9vztqU0fjtTdD0bKGgAp5tdC
IORpZQvrhhq9fs0tAQVoqfBUzZUGLPRhq1Yb+E/TTjpX4XVtQAZaDUd7LUR6MAjpu0YrWTs+Tr7k
UUjCKMUDRDHZKuvPopvsxPqVNp/Z1vCOnq/znFSkjmndqH2v7u11t8MU585o1FUOlbtSShdQOuBf
qv7i+3yRQE4DT3+iG3l2X2rYsXEBZqHiYPYiLrhf0jcHjc8PvH7O+tsh50+ca4/OsX9l72gUe4C+
zqdY5heHvWXCj6Wj2t0Yg3HNxjxmw2LWKt8Oh2wzNw/mOSXbCCqM+58b9lr9jcAOUIHRXyhnU/Cc
WtVih21/233438X1fBFhxLNUe6kNw0PE44qNR+mfQwfjoQiqorIJ4hzwlas/lneyApRn/CuSGUaq
xF7danH69X7cnTVKFkNSwdgiVnd7iSucnRd2fIOYIZD/JOQM9mfrzyFFFdsIOCsvX2Q+GM/zTR7k
lRN9Nf/etGp5p+9D+aTGxC/xj4xf+aOUKFwgG2jFqEMrpTgkWP5IxM2pbvm0ZDxUkeJymV8LmxD3
LTaUwiBHLAXMeTAMSQmA9GaqepKc5jgG+WDui8CSPIOUP8iwSRVkw46b5w0cgYTIIn3ReW0NqVH8
PnoP9cNyrT/yoIhDX2fLhbH2z0l44OHuiaHaqMOZskjV6ynprVXoOPRWyNytGUFqI0MjoRBBnKBr
4wq1ilMLL88zBLJp7MT5MKUuE/9Y7/62BF1LU9fhryuvPeFib9xBWvj3lmD1uA724UhqARwU0fpV
K6pJvfbanAGfiRw8uwhxL8Cv5Hj7FtxLlyzMWU9TT5R2zYp7l31ceFsfXnH9/fJ+oiW2++Ri+mnv
PbIaWCkNRNPPCLKnbrpsTW9sB6EtSpL45miz/kStZ99MxM6qQYyecI58WLXkb6YRkuFssirW/jm8
3eKImXAvgNWIiyuVPyJYqq+w/6lXSNb+axqWuF9mFXbf/3fgQJMKTOyxb3ZTkM1SReAr4+7HHaoM
xtpRupnkYh07zIr3hrZdCMJh81mJVvz7mLPB0DWFwYNbgsZ9co8YIge0L6sRUMM2FC6eqlQ0vHeY
UlM4FKuGN5wfBid23YSiQdiwHgAYdTmDCyDGTASfPuT0SkmGqnBfxYw5/R4M1YYLfAfT9UZvqMag
PszzzyIWdf+VO4So7/9nkpru8AWNXSrjjZP7da8gf6+T1FxBhPunFqPdPgilM7GM7nQP+VjT2ebT
SOizWXoZdeG5mG5SX36kUY/E9aNnjcYo18JVOgLTk/Epv5aOlAxs/im8kfCP0P3SKG4JT36GtAeQ
CJOjCwcvry/okijXVNq3N4nKD811hsDjhGHAGpXVeUoh06yxdQpFN9x5GDF+smoFAYFI+nSHrQlM
cE+7Z2SgPXU5j0ljVFFGdWbYIZheqDO7pomfpgzGD1nt0XPqa3D3/VQXxgeiThuh71lsnlY/16YG
RdBs96m2mG5TFvXaKDtkG09IJlA932JE2cW/8XcidK8xf3mUVF38kWDnqVrh/UPCyslni/F36ZJA
w5S74gK44ns2nzWQh7qhSMEmcHayi2QXqOyA1SMrv4O1fvArHGRTBq1fgO2NFAnC+dp28CDs4UiG
DcakX3qfa45m0zy6nMpXJ+MaXdrZ32SgUhwgytiPlsdAIxInb8Zc5DnJdH8m/eIhyCEoYJ8EGxQX
OmFi5MsS7o4mG5Fl4r2NwFIpRiojCeCafRlKfSOzp59BIA8C80ElYAc0fW7JyGbYKFFrL9W/5bq1
frgbDWy3ZSYIgmIOQhrM0DeF6/KV6XNcC/wNxr9LbwIcQTGKEPmDXAxiYBtw1EdB3DNama60FKmb
nKpLl9b+gXwH66vCRMBPlxHmIGVWOvKhBkMeDx+AQgYVAdR+TimJFOQcNte7mVu7re5058Nim0WV
wjjyQZNx1QJwbVL2vU7Fh2uEpFmUalzFV32aG466QKu2o7kELNdOJplCCF9GmpE4kST30B+6AjfG
b4QTs2nv8QaucMx4RB0UPKGB5p7fEgcqBq4bxJvolVBQMWrWjON/YTZFd2vIFU0NmnMhR0J76k4J
xx2RaZrWf/IpMzwKIl2d5F+lHnW+few5nIrKOhzNHfJxRTy6s9M8Uqs8ekjePas8cspzS8xKCM4A
yoO2NM8VMXVuSnQYKECID9VyD+HL50sXhDPeFRGE3XmAwubJJyMMTejFxvqa3x868ySIVCzD7RhX
q1DomFUEI6V9LyQvEozPNJKyzD3w+34H15bIeK0ZmA+j9HnlGRM6VcFr+0QJzStI+0PbzkuZbGZk
ijTjxILZ8TzvK6O+34HS0pjT5UjWg3tMB/ZAPR0JaH0/P6zX1ntj6WeQgV3M8mx4vrfHdumMwWqY
9EOdbVv6fDEXFSw7jfdFqv2cXtwxrB51PK+ijWurugAfDSjfJ9DNZ7EZUGIgSUpQnkNmDxOjXJKK
ikoFCD8jq0xwQ33A360XV53UYip1EIKJXtDKPMP6HvuvdWkrZ1iTmFq9r2oJMl0XQPVyxMI3Xnnl
hN8EXMThsAbVPeMvPmJ+K67BNEIuvP0eHUisY19xSVr5CcGZnx2QEfTVnmFQYIBdHQmMt10Abe1C
ndaLceO6pPdOxfQ6dNMLaM915KfZjwlcc21b/1Em0mLSSkaIo5D2/oGyM5J5coXyIcSY6j97rJbg
KWuhF9f3/VT6RovNnUqXN3Uphzh0ZSJgg70EtbUgIbf1cvrIknC+c2TcAtvnK+8kxtx2xJZyQZhs
jyx56XFTntsSBE7SvcbKYaBgzahoUs76dcnVsG5MjydNtrVAXnhCwPb84wULpv8abPMn/17t0iCw
XBNXgeUvFs65IY21rw4WHbGy0TBendGPVV/GrtDMBwrNVAmfRUJQ9bXPcvhytzi+lN4eSVvIvg4Z
rv7Qf/KB9SWF0fpbKVbI68N/tKC6PZBcOYAqV6NtG6Vg6KFEJvp8sN9e4yzqOuJ/NAhXBk/+aExb
tCOclO59MGoYwcvrfneKw1LNxU/QK9OtpLQ6Fj9dr5TAue66949cnZp1f7/ZGWS4CZ46DSa4nEvE
rlA272fJP8n96cYOW+gtF8G56z3YyHMrIuRjbFtI06b+CYY+kAxyLYCMXKtte5+75W0HrxpUcEQQ
26ryAXqTY8uiS8He3xRW2IG8xV5/ozYtIrN/KFD7Hy04qOC39IOPQ9NPFP61+NpRq2esyNWSxRxs
ZvXS12oHqEI+iMI/8mLiqUmU2OYo0uSYvaqH/AJ/dmunF0106VEeQM68nQ5F51hkLxRMSLgpAbkN
xvoFNBaj1CMnt2n8v+e41IVBu3x1LJZ5xxPC/uMjgIGHPnkpCsaOVB6UdgbTALx0lC2UE7a9ZZG+
DCFTjpSLFC4cBZJtTYoGVoCbUFnHiRJcw00N2YVSMhBqd1X8RY+GWvkKWXwueAMcwNBT4v+7Yw1A
DuxAgEL+QFQFE0v3gTqued4TwHkz7nSs/NY2KsS0j2QzRRdjuEMXkUrdLauwk3tqrcNuSv0I9bVt
kXKzmL3HPqvKbb4VuQcEvawD23Iy1+Na4+DBRrh0GsKCs1VxYCXsF0EiqQv6t7dHcjxeSInH5U0Z
DoUk/GU08OtKovPX4eIQzW5UpPT0IM9FkO0thzHKt0If3YWIjNDnaGgrrMVcEIqR+Z5iPrF8+E7J
qlFHaOITpcA8ekp1XrMzNw8QjffEUiV9oF0K+wRhJHV//vI4ToJ9Dxp8F3BiqUceaF+PMFCh+BmM
UmtbvvR2at9tcOVLg+T2mqNyOG5eUD2UIX7VOoMn9OGxV3WWmbEbbGJo53gmxfuiKV4jimV5yxaw
cuG//rVW7ViaG4IXGDccDsY/CHnrqsNB+W6u+BNyyfspEnSVQj42INI1FfvPEQ8tQWKfQAi4Pc7r
9r9657TJduc1zgoIMzO1JDhYQJ2/pCnLcHqjBblcdzCSutmtDzTAgORtSMZSYbYaaBnOp9mJ0uCy
iqH0e1SonGjb1jrHcV8trFWPYEFFPnIJCD4ADT4PeRiqZaxL8jm8q9YGiHGLdgdzFzQoIzWl70Va
h5MPkk9lC7YSQMRMVoeEcI7Z0OQGBPfc0KO7kV5rHXhC2RyJ8/n8VHsE9EO80d2ra3MfHvOYjuKR
G6hTYItV4vMmL/CwQaXFUNRTS/zihcj0/tma1A7jyytE+lpKRFm0HxUgSLf5TLmRXdCK86kFWl9J
5uvUrAUI5MjYtw3AjrD7jJnCEhtJEHVmSP0GypiWMoMIOmvXgdmNq054BZ5Slu72YufZIkpELq7p
n3sNW0HpGxS96Rr02AoK1qVhs85q18EwXt1zdg/2+C2KbmIW0ElBm62I+8Wg3uC5jjfsrGECDQsx
1iyS4OX0i32Xgk401lyYj/W70P2RFimp1WFhKI8YCXxtLF1Gy2ryNnwKrgtOzUYnOedM/EuhE4Py
TcIufnL1oODW5wQB8LKbZoI2/voa41/UBsAcXYRLBbpHpZrUJTRvPCX0x0yT9U9skBXA7EcCffyQ
otCeVPEWyqDzS+Oy3s6YORgHAWiyN86uIA6dUhY1ctHNZw07i39cIQPJWRm91pEokr5wHt6VoKOy
afOVoDlO3O1XD+t04jDIYEUTtNAdmq5U4r+wVWpo/VCB4uaDySqQjsRqtgAz7hCVI1+ZaBVOr6Dw
Jw6NVBhNihS3eFnHGSRBxq8fdN04bP0E1YkQoYUjRBhB7ssyUaXn7PymMNwbJmfP/YOp1UFpD5rR
FREXc1Rofc1RMgnjZMbynqCX/dWLbP0wFXGYVvjW4n4ySzHmuOKntnLysOkla2UDBrLcaPIUL0Oc
2xUH4oTvLbA8RF2z52u5RO/zU0F29KZasHSQNSCeIWx6Ul7Ak5QQY36kQLXikmeKDeO87KVxv6c2
DSZBZgZpW1IgMUU3lY07G4AqhZrKoZ0RuYDLWcUAOX2nxiKuyVq7ENnigG1SEGTrj+2Omx9WEASf
K3g4w03hevqk9r/hXBVvlaLGc2OiOxGOnqXBI0fBUwBN2KKJeleoHVXHJcBMPoxe6lr0Y7EXvOii
5xqhYO5osNv8hiwLL2yawHiIMb6uMa56G7ilkX16wjTCA+nP+6jBFFRYDJYU6gu702HxrEPP44Q0
Hj/xoUasjngwg4PJsvnsHKJVTxavca0HOc2qxTIj5b/Zy9fxpJWaoQoFLUENm/QJFGDKnRXS0pUH
Ha41IolnAJqHaWdyWIcpqaRdxgo0xxthBFj8k6Hpeo1Bk/cDOYHgHTfYRKcHsprNl652qh5SYzLi
qISSltUEdmwVWDwLUfpvICjhSj9IzjHinjyEcHj5JqzjQl1enfWMPrRjXWeaA+WB/6SL4f4f7U94
tts6FtJrVLyYCpt/tlGnUzzhwIiR4Z2EboEyip5/V3VhWmfn1Iz4+Oei/8YOgL24Vv3jvYUmHoBe
2yzA9Cs3hVTtAD3VXzrUzJSENam7jNfP71L49B28ac63w67MvAMsLIi9+RoGXhbnO6zuozcXYbM7
QvoYPSAvKGKMZ8k+r80RNd5KCQyzcUaQoUgFTRgnsLz54e+1lcdBW+d6f6Byz1iSMQLpQvj7jux+
HgwtMpp9VEORjrLm00sdSHoRjQkMh8PIwCFUoC/Ykwlow9ekybxctXGfXu3Aky2AV5Yzb4ldMuI2
5N6jc0BSg8xSv21ekeBIHXlIRapdiN9NYzrP0ZCT1FZNevpQGxQglKLpc3w0Fq5IAIiAU9/LkFvC
gb7Paa4ZabRpAozFv3LlDSi0+5fRa3kyb5u65aoJYEgJgZlx+UEnTDcrWGcJ9FqzB5pfDDG77ZMw
p5AfJm7rb4COTVJUptge57NZM6qR6Y/Xj//kCXYjkkOp3yOLMxEAx5J7AI9nMgXLckLMdWf+S002
TVoLUUhR7wj3o21x4u6nAmsnPdLC93O29t0m4qqyUOODY8lYjCz+pwaKVqFPjpUYx7dZJ50hp2Tu
cfthpW9Le167pZ20atbHCFkYh7W+J0VB6Wo+4BxHj6wAlfJHs/6cvCgtbnDfO23W/f4cQyK8iM0s
vFaTW6srjFdBNbTNmQIoaw5AMRpYnD4L7ftuATNV86oPIBFtvWpt6t5fToumuXuoywVmKgtqgivL
Fy7cEHF77/aDcKPD8Xqt7jfTfv3Y13HHww3NIMyhgPeOeNbyeHqvJxiBh2KOmkUu4J4G2Ul+aibm
/eIVQEooQZ57P22XyH35GyqH1Gm9JM1UzbIix7WPNLPRYA5OXXAY5kRp18WXjWLmJBt2AikaSAaJ
sO+BioH5nC2yV95y+hEjy0q8qFk5iWFQ4vzKn/t/rMcJzL4aS0ayApje7+hVml/XsYMFCFgGsLs8
qftooMkCs4QUzi9rDPn0OfoHi2w4rnLPSLFZpC/ea73VVn+dF9xSi6m1QeC16apeVs5T0VOQI48F
Wwkp9JWc2c4YGXzjf/Mdp8dv/mxh34d5Fuw8vaPiISgfK1Vn9lRjuxgIOAA7OIjXrlqWeAq7omyE
fMLGLaENCoi3DUnnQSQ2brw/TjNluyhh9qgoLyCaVYppt1GsrvG+om42H9rJI3ePqVM2edDd4zQX
aGgdUxHn5BPqPXTEBOp3ItOYQoXKAqFNQLLgUXCx4J2MSnCLjEPmiX+p8nBLtEF+RH/gsprII8bv
95AZ2aAwrxuy3dh8RcRMEKhnNBI5TkHUNGyiApOIAOqMPupcLmIL3OWb29tqd6laY3+OZgvJE7cF
aboeA3gyvfo8V0rRtTCpn1AaXsyjOX0Indu5T0xAO2yiYHTaeEXjwx9V1XV73mvDILy37KMM8Jd1
VRkdJc2bWG61G9qXXsR3wQiTphzNXejHi/K12elZBp9xp5bGobmcF2LUXAw45pTaRY5J6tp3CnaM
NyODsNGXEUUxTSY13Y9PTw1RgGQUyS8/op5FmnPgfQB5KmduNGukRY7T0G2Lde6ZE8FHLpUmzJSc
k5lUrIfmdfMsdy9TepnOMg/nxymgKqEBRwA53YHrVmj0QmQrbHnhKclE/fk0RrMNSzBTNNR3iYfj
iOHbQ8cXJQkZBWa3q6iA196Uj0fRNoO0bs+KCpWeDHVV+5jRLILmNX8CWUVRDa43dZLblwmvFn1g
nA7srrWerT2wn4ma2NJ+fHMv+kKQefwh8SSWu3XFMMaowUdKLQAfQn8BphWoYo+h5XaUBvAZY97S
4yOQ8HzY3bki102gfnz1vkmYHsDotwPiFlPYhkON+QjaojffOE4bpaHCpjAKJWGQ2cGe1FhA7wg0
yyjqqhlJKU41c7nHpFnyvLTBvFH+X/sgnymNml+/OYtstpSLESzHtxTgU7VY7jQCwsVwToZTNWaR
6Tuwx939PxR21hfMu+DjvkhWrMtyowYyqOfLaTUsUbtGd/RF3tR058ZybkPm2Awqrdhy+f/rREkk
z1whQM6cvExnRU3Blo+RMT963rLUkYSBK+n+pbfyaKqy8ivUhxifL/7EyIQauOzqH98mtd2logEN
2c+V4w611VZ2rRIF6oU851Ro4/Ycc+UW2Z8yE73daH1uz42RBq59nfjuqO9NumdPIPj9ry59sda2
XXeDXbdIyQyfd7W+xD4H7J+6fhCeYtceoxud8x8VtwqafEK4nkXKptG0I3MzRMJ1Kf+Ew5vxTWBQ
8QGW0GWMwmfYYv5gdNkAvLCQTD4TbAlZI6ox6DqhCu3gOFStbkyo1vgqiXPOIDa/xdzm+raGYz9o
ESDyqFqEHFqtST4wsVzAUW6OfDamkxYr9SalgE3r9Yf2Em8iH8vHxnQ7nKqLxaYDTs9LYYMAsLgS
GfIR4WvITH5B6Ho61PYiXPBWS3FNyI1qeZf6Azr2/ybUq4i01d+mawxFZxqOcNPxUSSHXF7cacfF
10JeX5/0InnbWiF7S6LdpxBr1+P1Dok7KYe6+Lu0568GyJGhgRiDUg5lS15W0RPv/6Q9/2G2sWxF
S6Zy3/HiLGa3Vhvb4G3AQp/W+B9h9MAKxtV0BQxQh0XFKtzJ9guuUghZhZ+ZejFF2mNwvgslrcAM
sEMSqQ61XP9FZp9hB+mP06p8QhqSeKt4TdRf/WBRic3JTzG51t0nyDMmEHPhJQ2vfbDBBs1ceGL9
3upcDeIH4nzBtl69i3QCaGK/gnILBE2MlWEyq1Ph9ewMIXXAO7K1Cdkj3cNaI978JRhuUgLObtD8
B4rkpLpwABQUEqAp2t1QR5T4syEg+DhLP6AS9784MnUtmsSRoNAAK01B6qi/cqWAjlygj4h6kXdP
bNaZbeZTwIC5xGZf1mG4O6kOS5s8n3z9f94e56ztPJwKorOG8Lyvr8XvYEuohDIh6xXd8scsKqde
XFSnvBawKLm5ONM5utmEGty3ogsj90brdOGneqMBtEa0z/CVUzpUcdCkDEibBqy+a9LKEDktRNpD
H6mbFqcQKRm/wELlPqoUxvkoyRSHwVij72gyfjYrSkt79xJO4jClx26Vun0YxLytmUFUwPRkSg2f
SswxLIBiCBwDSlQOlhLmLm1hculznmrUhyNpvTQnbrpA2r6gQ50D6SqfB3IRVPMkhyS45dTsjw0y
IlaaM4xtFPvbc22cpSTMAZNK0XQCWUi/SxTg+KyKUlkoT6IODfu6Pvt/jkvlZRVTWK6cvkATanbD
Fm6fp3FS48PqO7kmXkf/1UTAA9zJQHbZ9oPWGnrxlgc5jl0Kcs2dTMeinYG9s95xLFrP1eQeJVS1
ko/p+QHnEjT2xrQcPNP2fNuk988jZoNxHVSL14bamFFjUrKaleOTVqBCGEfYUuQdu9U+oLXf8VhI
bErxR3wAphsrXSc+PlsFUMTYxavsycyITmpUx/SUgirgjnRY+hlSRiHV2BY+ybMFSYotfY1hkuFN
Yg/iVvU6KxexJAFypl6PRCqMFSQxRVAecW7uTW+8kj7dLUHwvhrF+ak7zAgBxWru2gnH516l6g/h
PrSY5xLjoFaePOBvMTCX2VwlbUQPMrAFIHpALIBUv275CeCH810PYehmSeKsY1ROq2EWEYxhW8rH
cuWcMczJAKXMPuyKwZXe1Y+rJ84Y/bnr5/s3uzdoS6MasfHK2OGPDFbHbuVXprC1kglENZt8XiSP
0M/k0m0VR+kyyutj1W2gNLon3lPrBgbVQi7u1fi79BRjt7WaqqTSWCEcf6dgP3jhPL1xzPf2CLj8
sxIlkdKJ6ZtIIyABN4qP7FkRn8ImxZ3xGOAE/NQUbegs7+v05Qa4sANSKp1BmlF7WP6VDZjR4LdS
Ro+jHVoj9xAJb2xLy1I/QfQ8yuGdpEh+tZibfxNRl/i6nuEJn1gxaL2w9b7JdaWAqvdt1x1Eeac2
NHOKsBQTOEmRQYj94sezuTht8QNh+S+yHsG7n4WSWBj8Awus/If2rzBhZlEv++bbMotdbV3KOxgt
qZxV1G/txKkYrfdIee5EnPqNQ4LdvFnaukgvg3GCbuSSD8GmwDZRcclf4r81Ry96CXTKFUpu3/9H
r/1O1brs+V2VXuoOoMREs9yJ085wdfSdHkDpMu6KWZoH86Izv7uJhWIr03wLylKiKOB/7ZsColjB
F3UfN7GOXwjliJAfS2gv4p0ypLpPwKLxdn/FG6nnqmZTNN9TS1Z/bVqxoHpF8RB7aPqFSvFiqR/Z
uAbqka0Dm7pPGKil5v3vYgQfc3+AY5U1dv0E40Z5FbflnLwtlJjl4f50giMGOHublm7hSc6SsqtN
FpeV34QFH9Sc/dwRqoi9kjOKwccSFd8PHjWn2vOMQUhNYfhY9L+3Awj+V2D7SdHGK2b3Q15KlhI7
aa8mus7ZBZfj5xTfrLPbM7O3s+POp3qsV5PRIqvLOE/DMlBIqrfU8HXBIfuQmpkDoH+6+auBgRj3
veLTBykwp/eNW0lUSrhJn4FeE4jm63AN5Kth53mcYM8d7FSScmLkw3DUngkw06dcJPjG7sfh6AWk
HxlcvOpmqNsjAOguKpp/aAnt6+MkNHVL37ibGh0GjNhtLXxRnJ2hHc9ASVismZ+hb6L9vZd4gre1
WGzjnnxdhtfRxI/MFyu8LjasiUhnNkE0f2jluu8dXXBHh7VSGN+g5wEhClWunUI4t6NkjpsBBpL5
2dX1+yKpfRcZeDJ8uxeQULt7wAF6wiwFPedt/8OYg+J0L8skX96X8EEVSxp1dk17vuoUpGsSnvmT
bNBhK7xXiIA0dCjOyIQDuxtaHCbeWXjEUWBs/piMXMqaTtHfefZ5g/CaJPXjX8uz7c30ZT6hy/YR
CUKaQFp4xaQo0SeTO+thaSYRP0tVXBpG6xtesr261iS9FyzqTZEAMTX5n8hgCI84KgE0lvKX4VwM
s/8c+F8WqCyqGhKjtTw5bpbzUK3rFS6hsKu0ZSuGIE5HMHvQCKSPb2Uqn0ewvn/tmRb8G0FGcmy1
aDxHz13gFJAOtMuGQOe1dGbQKWF547R1fvxySB+XAJ5QfDn/zCx76nqYknmWY2x9nL6Qb2l3mTkl
UBI/ygqLGmeIqlg8w4vLTbR38YHKBXUcJu007NIMWevaQOxcfVuI9sw0cFX52ggj/J2PCh7roBBG
ZiUvl46n20KJNBdnYwsl1nfsixMM5C5f+fIgz0WAFHD1l6AFvj7EcOoLVg6PGMOMF9Cnwz/BEqLM
4osUNHSQSum4KXiAm4o4u4IuG1RNJ+kU0SIQmGVTMV4TqO82vpNFYAcJz2xdzExG2/s/AsvhTLIP
Kfzzy/AhNUkOSCKOCKkn0Jen+CAug/Y7qc+dSbv8MYW6iPoM26hWTqTZkvqq4tO90Z53TX8Ax6op
K6LY76ZFMu/W3ADdQTRM5gwKPzZCVBpg0Ifw+Mp9rqHeahRcDkNo4wzVeTWicot7ZrhuAoFoftQF
RKAqKcDEEcOzvqRxhmP5h8rTZ5SOtkr9oI0i/SjMt2YsUqjIRuKBpgEd3Rj1jQhjtBXGd76pCdG3
P1cFz/Ig3PPvSIiEOFs0GWXEO130lX25Hlqy9f1KrliCUOzbncIMTb68yBnLolvu8cNKQqS4J8+0
CXeJRjfA3XVi9g0Rc9qQ3+bGTVAxbACNCGzmV8gfVKua293xZ1HtEOg2Feu4NFcjg6MgZgiViXN/
w6Srp54vUIVzLXERHARvXDd6U6UJg8eAxlgAO1/OwItj7yatqsOjzJ7ZtvzLEhShAl4nN+BPVPsF
noL9lfAC8f+1TR7MhMqRQ+PunolAa0g0KHDScAyg9YIfxTB5uPxoOssGW4X0HGZevWpPBa/tQlL1
09vGMWH82+V2Oql+I/W1CCwBi2eO8XnDDqWJBxRyxki8VRxHOOW8sl9a7jbSevlAcfQfoqPFefBy
UyWIgiVPzXuHruQVD1R6xq3Ob+kjeDjI34WtTCH7EFuvMik+9TNU38o/l63tdrRVjBzKNlgFWyJd
VnG000kCQeVBPzZn4uqnJla55Gu3Z7t3vK1lXPqHeIc8mV+oQdn7I+G31m+Q5GIsViEDd9mWMBp+
Muli4t5+hTp1Yl1o7b4/viSNhZs/E/r5pRV2wc7M0AmIPRUPIxHYfr4RFld/hVQE1+MRyAW1o2qH
EPPaGvBP3AyM3RRuHY1JP/nrstuZhh9QetKIFjiBeV+mkmh+QPNvwrGcYskclSZWL1EhUy0nuDv8
MvqOosfJ3Zyu2eY8mgUP/gCuHDGoKfSBY61KEwT/z1k3RfTHWfQldbe9sUndBjr0/ebH/pTRVZ17
m6FP4EQoq8q+ynfMUT3BXi8y22s8WQtXuY5iObHzC/1HVnpSIEujHnD5BSBHJdCk3aTx3ks/myFX
ovs6hlkWp3ZvP67Vv0soId3A8lEhxk3u2SSTBrmEnrgAhGvkEXJJ/TOG5cl2pGct3G0sv5ZaCMf7
PHz4kj1JQZfHFAxRLzZxIlellk6LXmjYZHGPxYJjrAeRzQpmZn2wb9CqAxcVULk7bneJsu06s5Sw
GFA1u++Zb5GOJKhI912tJ5zcW3xma+DPDM+Jkjywb0rXMeqViZCKS3n2146m0M9Y7hEdp5V29ZGp
xNry91mZjJhtXMaW8AF3kw5GrfQ226t7CzJAixifdyQo5lH86XW0XGSjKLBqlYSUHW9Nu0Qt7LDs
RRrtlOyi0L8H54F/zQJ0aUvg6X5da0Q02itLQ0LjojPqNNvmqy6lif+K33uk6ol0IOr5D/SQE1Mp
2s1ZNWVOJDV/4LGQwiqsSfrvjWh0MxH8TKHaERiLnVF8K9XkscxdUzaSpJKTXKviZJkkpg4kg1m7
609CFH+crpp+XU5InZo8itA8UWu//O4N3RX+7USDjbiCYXGMAgUsXaUvpoTqZp3Ect/jY5TCF/he
7nOPRVFsUTgpPgYf264Z1UNbvH5cFbMNhcaImhXnsOb0APvUi6RBel0v/KlI2LJwKB+rsCpaMTLQ
t6Vh9EXBkkIZyXsMykqr5T8nDeKMc3riQXe+b2HyuPBcaPpshvDX3UcAjvrOSxaOral3mVggKj23
FnPyxnSuPGoDWhQPpLwekk+s90wKF8N0Rjd2PoqG3F13nPXm1FhsvhbGsHP0bNKI9gWHuZc0+SpL
thHO6dydmi4FU6XgQjub7VVo70n34n3EhT0OW8374XTK1YELRT6A2IybWyJNdDrB/bDhmhhO2Bo2
iYfCtHLqXmW4F11UEf+lJsr2NW7EaQFO5bM9tSUzG+mGAO5qq4+j39XxjSjGIqGeP+u+RBiov2lW
9C4mPVyqtIWrLKG/iCJr3X/SR2d31ZZP35OfduH6DLewp69DL0ElqnPu88tWDXusxTsDfzIP7FmT
ZUw+FOA30HFtE21U+5FW7ge+lbO7/9I1Ho0+gt5KAQK6BIhz8OSf8dKXir6jAWqAy4iIpchbrrhY
Xy3XuzddTMkjhInkT6YUZDxInFjFwZta6uolGc/H+v0ixwG4k2KUxGIJk2debgig4KiuyDG/MXrs
O+X1YJyyUhSloV8MN0v148rHZlCIbXnanqiTmcuBaNiiNslaARLe5yaNbwbO1hN00ypYBBgkEOOh
3RpD3lGoQQAtVovlP3x/GAmWO5pyYy2/dR75EZPkQLBoZscw5+0OqDHHt+SRXD19l8LlEjmoipNM
Vs3E1Is362G28LOhrf0dEqtIWZUSGC4QtR6uQq6Tj11g+JG+HD1+9CO/jCBAuQZX3s7qlucKWYgp
LM92bNkk7rBr8myLR6zDovZD/7JAc2hx5tizSnQI7FE80+8rjQ/4cNBQw4K5a1EDEKB+XjRggyuf
L/Ir9nkIUBQtWZhVbESa+9ybElevVyFBxVGIKP3+GBInBxYBMpE+n4/Nf+5YKyhmzejA3I9lO3p2
dUeNezfnli8N+fKTC5YXc5aNLymwyd2KqpYBxU78oojeWSp4SI0HhcdaXUKbN3RxpSo5x/aeIMt0
8ghksTfT9me0ZH7y9Eun0hkEJahfFzoLFAA0rw4lDFBbuuyg6dCqdDJkudMoIIXVLu2dikZ2hEkl
q59L2BYqdWmNxV9LLlamioD9r9mD2K65k34JExrUUt9CyenN24YRvkwxerCWoBfntg31gf7autW+
1+2hIRNNWKpof6LG37uWp+r/kPerXlxAbc/0Ue33aVvF6E8bDV0It/kk6OlZiGo9vWlkrmu+8aEd
oQXfSi5gNZbq7aiCr69yoDSvvnD73z05uVBiU0lpSELFMUOt4Fjj9aZAcLlQkX/hlJ8b3iHh985p
mV06QaCT7DS4wDacKtoZn0MdpJawwu+Sy/UmgYCRtEY2Zu8ZOG967GHtL/PfO0oXaMfB+SFsp+YZ
uqFEvu9RtjoBXINZyDIok7vtmhGI9G7YgNZMhKbyre5ZIHtlEyK8NyjPCjgPlBx5awdBxHChRnuC
4UAfzoeJpIgMRBGykJCr2uFQu5a9ORL9EEI1R0IboC2hQwEGQqi2E6FDW4AnDO/m3AkcY1pLUZOh
4SW3iR+EVQbSVPRhbC2NXcDEgRWm7WFA+3HqFcWKF+w8q2qXuAa62y2tYJ0jKJ9NKNi0C3hNMy9B
h+r1HedMdiw2JodMn84tfRwVW4PY1EHp9ZssygIpWJwQR1N0MkGo7B57rANRZlgiyh9RBwtb/nQG
IiMPoFoPIPa4Ne2VAo2JKtPOemh2e7a1oYUlwKh0JVfbxrbaVvAzoeyNlr1IrZVBUc9B5CEK4HXO
y5WuUAPcGOHmsIe8SorxIr0A3xsmUzgXgCDGgOWPr3dTfBKF7/5R0PMvJBPYsVmKkuUU52pPKRx5
da7SKRagXg+HG8s+ZrLjWBiwHY9tKfEWIcDPHLlcva/jqC8bTse9dPgcj6JuakNzCgtN7okW7vys
0O28YKbCXQMJ/sqpg+w+8xWsi/7srQDgH8PsqrGXBmBc/x9EuSOxNW+EBTCnFMQ4dHDdlJ8gO2lA
riTq8CBd9LDdwwQrY0M6+KrbPa7A5WObdcbTtB3kf9J+RO0P0BTK82MJvXP68PFkzDqMj/tfKs6Y
XRqXU1etrZfv/SI9ctIXHy5WmirKzr1XgLqWBwwGb/s0+e0NQO3mQHTNUIEwux39Dv2EVbzAamKF
wqlkrpOIjxQMdduAH/Rm+mrGSj+Fgf34aIKOtWrS5TL2ntEZmpklOZZ1Ekqe5vMpQYvp1YDBMiGa
v/+I+D0hyfoS1MI4iLq+W4zO3Ild4vBd+VOLZMoFzIFIEp65KdrskYbU1W+uO+Y0LmTPDCOvkX51
iNnCZum+TXrQpD2j7ZlCvvBSY5C3VoRxhOoC5zDLqk8094iU9cen6p1psQQFdolBFtjOCYI3aPsa
Hf17z23GPVrgyoTgGpAOzqMZK5X67/2QS19aMVIi18/FUA/IQKpS/T7qnZgCtfeak/1UWmk6GiUs
4v10FOJbhzPvacTAr+b9dFeVlmE34Qo7MrzH/dk49HghQGZ5nDxAfzWxOiUxGDspkVLS9ta8KzVY
vOp12/NYoy6m/z+RAZd64zYS0kAFUS+UDjkxBh7zDk0TJ1GxK6pYTIP//KHdmMdm/PV3jZOuKdEK
NDg2H3FehtXutAQ862VGOlqfIvhtqBL42ATlKo/WcdqT0L0XDhSquxB/W4Xym3X8xCQk9fV/snee
FtD93MJuozdRk4YKtXOfTlmTiJnQ8M3PCJgbl+viK/NQfDZKpPtgzFfHHs6MdVWdGBN/Uzk2DZFJ
HWh1+2ZtMI4XVrQ4VrfePmekQbdlkH/tC/3wQlAriAP94y1+CcXDOxcBo5NWEn3bSvEHaQhKt1yc
ceuQZBXEuoMpLEP9ENEwTziyMIym+ty34tcvTMLo2H7ZSmEr0n0bxoxk7w1s/7KgJ4yh8TYdKD9Q
5jSF0+8vQHNTOzSr5VjWzHxFFCX4B8TNh2BnsQROQB8CbvFPmJ/woKjtHLnVP8PoYQbvxkdvUcqp
+GNhdnA7e//m4DPNrTubbp1oNeTZcnkArmtSqb4WFydfgGNJAJl0Ockq+VUDo5pDDfk9OSEGNXLs
e/saAgF4k/D6pj3rrwBAIqWGA78jxj56tLm/PNVlgp2pzZvlpSur6c1ccHq4t+OPK+QHFAhr3XeZ
N0ADE+Zv9O6hIj7Lk3p2s/uD6ukawNt1bZND502eeE0uhtjEJ8k3ypDDBjV1MTD2dUNTPh6IPNjO
Xv8rPE1nMMoUJofBOVG5k2API/aJ5dROZp31DV9h7Kz3UoXnbmIpIli6NEP645UAy5jo6exiojvY
lhqShNNaoOmGiVea70F+IHkYtvkB3lll2VSWEKKfyDI2MGUC6ylGhlgpYdieKVf0D+UPMhb4tVh6
GIqOiBTDvOEoufOBL8HPBSU7TF2uG0NDiF9jBXir3+zdP6Mv0J6PnVELblEQZnz6/hRmSZYSHLhy
QGh+tGMWI8UuN6662q4MHE259NNiWZFhkAWHLgQ2qxR0+8JJnzZU9H2o8/LoXPJjpCKVRJNsq8hw
rU/2jvVQZCNchAIFfcnp48LVtmkQ/3J/Dr2WucZaJJ98e/jsgAurhbX+UkLmHy+1r1FlWx8yK0vy
zKn96vlOca/b7xgWjEBnTvXR7QL7wgpuyB4wRD2AbkF2SeqlEneTf+Cw3xP0gp6KVkhSMFa3kzMM
XdfLwWjToOg52YIrlb0KMbR88xlA23/9VzDOGns1lOdN7RYcbUmdzl3gneNS+dFRrJ7QKNcYQhug
pdCnpv/+Nf1pdG3ECIbeDusuvZARubQWC7Uf6M5UdTK1WuwyTsO49etebPEVj4fbSbSgBxZhvbzl
vux4YJuPW1th0l2w4+RdHp6VNk2+7vfoz3VHeNM5JPYxEMLdwWKzLg7oEon/2xVbqmhao9x55Kp8
vCG7Ca0f4+Fcx9LCYjozXlmPVCXVY+VmtMtF5G34f2ADju0kh6jPEtN9Vygp9OtVfo7BcZTId/Td
wC20E4FIHyM3HCreh3NWtQNXK5sVqzxdsmC4KU4icFRi0l8AZPjvuCPeQXZKOFPWYzCSRRCnq5nr
2FINSjYY29LRJTC6t506O48b3OU5qDD6KHDUVn3hCmlILlBHf8qAbzFVL0JjeRdkkYOELq4VqDSN
42gIyH4Jsi86rJx69tpEN4Y98eiRnA1iT/eb9HhJ8que/6sq88RQYgQaEjbqsiL0PctfuM6UjDoJ
Iyh6uh5f3S9OT7VhhzNp6BJgOaoW11/oQkJhI4KP+Ih5GEloDN1Rxzu0Dw7dFLAPTQ2WZ8IAmHa0
flapdFZFaIxFr51q1x6BaTWkenYiOSpk9yqutv20e+c5meOebigl6lHeyOPDqIHU53BYh+RLtO7e
dtrrqZLJ2uHG8yNbeaBQfpxT6oIGJ6/8kF3uUNcrKjGk6ZbbO/QQMieDKyf3FygRWTqU+yytsI4B
gR0AHB9faKLjYDNLgPbAJyJ06FE4OzoXN70Jkvs+YHdxCSJN6ySUDpCE3q6ESpXVKwL5RUASnOgb
o6IjqceCFNJU6ANgRs+nEIykJkIKu36eTVHCIVvFZ8rchnUiI6y3wjeHu+o02Sm/BTwiG8x1kvXS
WAp0FyONM/mQdIeGh9m7oaMG1nqR4z42WqwuF2GR3a8THcR4I3slrK1CTZ8UB5q+ihP9oq8skG2f
igAY+i6dOtr8LYpESrHsqvYzdQtT9OTQcPzkmp4uWsy4C93T+W+M6xJRbTHSIzG9MQJF/BDySDHs
N1kLQPo85RMYUm4N8aajW8e40mDQv6hNifxDHVyZ7er3vKV/E9o0RbwCE04bD6fxZFB/J1gkiWh3
PMrOyY66y/31kfPtg0MdpR9c2GypgPd0mveJVmSZtRrmc1u0r3PGGCkxt2pR39VgjkBcRamBSuC4
J0ei/14yVqzYoIEwz5jKlkB50F7Ykh/bOZ11DntrbfJ34OBzpVapO3+w5WXthPbv8E/tuGrgGCWW
3mGBC5Q8WDlSWkM5oIJk32BBHmiqHv3G3umkZryHirLPQoSCxWDr8FWQA1fyfDI6/usJOOAJwrQ+
vPJgIw4YicrVkJAD0aztZx0bRA3DwLGYeA0se31hmdjUn4iPg7sVEYfOsV5lxdJCYk90HTx4INl3
zATJwnP7s0uC3jIkxmRzUF3NYO3KRg3AJMV5yuobH8TzdoBHYWrwf8Q6My0GVOKIcrPYOvFI2w0i
MZfedxzKsFMRBK3/yYToclRBxazSw6gQLl3eqcK/pY5ejUnk5jCAyPWSuJ7Km4WUVMnTmg76QovL
k4uUR1ysD1cmTKoBFyj0VipsmD9hvlwM9CaDX/X6a8Wccforasgv07jA/G+rp/xVI+aRQiIQBidq
Y3gq43reQRlv5UIkavqZV14kWmsp9eOTKC4Eq40TROmIze/4gNAsm1aXrkjS0zU2AmyeuSiJ13+J
5E8/0vanBAQtGfvI7Jc0v4Az9JjqNtUH944+LREh051uTPdSeRjw+qWrz9d3XHkNlYMNrHFhJ1GT
jizBUHMxR4sullrtSq7Tb88OgcHwsyLD3we0ismHelx3VXsneze9s5HVZP+tPJWK/0qD5qbqkei7
K32oR6ARlSj3Y9Eu2YajHHpX7PhvKIh96IwugGDwV8F3y2Wc0RB3oKxsEod9zK8BoeylH68L2BqI
ap+w9y8tRhxS7pqovN/M7BqjlvlBLiEHfBxzsS8tTchEOmgv7oOU7rggoOSYMQJFCoNBrfWG01e9
x8o/Yl0TilJ8HAhjqJM3hfHXmHVWccbO0/iYl4Ii/P57y6ZrH+29DFjIZ42T8DlxuiLk8chTQy4o
6xWBCfcvF5OaUrU9xiFtwLk7PzryEIADk3yts1DDr7wnTJ+A2GZcolC/dqgpE5sx2p1+dMo8DrO+
L/Tur7x6UXcM33B8sgTeL85Q0tygjvofjQHVztAYFsg+Ide0T+xT+lezaQZQ6V6pOuGk6aux/kav
K/qV9Fg/JzrSrCyeOrRmenuSACcH59uKw5pGtyNaWwritJK8wp14sf/pCXD7ROhurDrcBAo/uLRQ
lHToYRagNS2jk4a7dg0kCFLh865sbHUCHUflCDEnflV/90xrfqY3uesX0IYyVoWsZDegJ5vtDgjn
qrzizzulYXE2OiOSHGtm9L2ugQA4S49j3nfCASMKvIvy7+TvW9lQEIsr/V3JWg4yPCnZfCfeqkvS
sTIwbx4sdtUNb0wjztNIV/fSl4raygzdegaJyYfG8KeTmI980TBqEWaSh/5YrzHCPAISBLA7G46q
HAkALoZi6z51eM7785fGFuQuMpUCaDETF8/WOw4lA30ek0Jfbr92IcH5X4RHZT1e7HHC6yeSuTLU
sd7NXXVG0rtwlT0aE1X5jWRtclfhrz2P8I8rOJUGEr6P6jOGjEZMXW0s2HhZu5MsJoGM9yJu9ZUX
jAWuAfXCsmJz/ZgspbQbeb5VFB2+g8OKp/qg5bTI9WPL3BWRph9Xl7jQvlDn7bK3eVq1RxfgmOgJ
pAUStIdpMyIxwLJhrUMQcFn1QwyQImy8Fw95POBNFLmQsL84DilvQ17ldsN6FHMx03WuV6Cm8ihx
pahfq1P9zSA4OkQFYnS6V0Hw5HJTIUNYdbLoi9Az41C0dLSX2HlFB5hr0NtvLWairfWTVPM0lxZJ
0EnbF6uVuhti8GHxdpZdvwvVG8QwVg2an4O6vyXc6fmpMhRVXK8YwlkmloBQx17P29FduTqR/oEb
e/kGn8rTccwTpnTtT2SdNmvusMsrwQ6VKLGMTFRybofKXZCQ8aKxVYbj+NWx09QpfWtBNvvsdwa3
ayc+BLWaXrzn2DqIyYwN18WafNv04hGbbi9auGSn/pFzMdudCl+cu0GzqYOJuhZZCCvK0uWkFNdQ
OuTEB9/RgmlMG2Nafc1Dnp7MDb/enbBbLGLdSg3VkvqzyfcvMGYQ56M6gDzIYPZEm6reJNj/MRYj
2q+NZod437YdRzvc+3YCVyHWng9rlXAoqQKuGh+iIe+foExpjO2I6Pd03lK6HJ+R2lr6g/iWUlqC
RiCYZalCeOb0VdM6MA9HUCU64GSZRQCZptp+xi7rJkYzrPNWbeCjQ7gnlSp1/ndLNpkVL2yYYtBN
i818/DLX+AuKC+XmbxYxTr4cFlk8SAFJkLs146S6X3mecQD7HNxbV9OOA+RM3iAaZRmMp8xSpWYM
i1Mhh0oQGqVJDbLgSIye7QSvDopbxauXBWleNii3ZiLJMYJ2sP/fvYNsuG5cV/eLjFWtnwoVSISt
M0EBaxWMbkp5p0ZkCOnwMDn4uD0XGqfaDtsr71/f5Ggh9wsqheYoN8xYM9GKZap6zuuSdtgNk460
4AonHu1S846oijgmgjd0kIHQiV3P5vb5TvhHi9oYxcZx88n4NkFuH+jAsNShBfAa4pPCD/u6RqaW
tnUL5HIwJQoJ7DhBfVjZvX1OkwRf7U9vWo31vKEeOzUShKTXOfxyaHhIKv65XsR0xXd57I7JaTYI
rLii6MoSOokBmGF0UyCxEQMp8vK6BODzujpFJsRhJNfS1lz4HGofxq6ZqTKLsrdV2xIrKqBUsBBO
ZDcMw/025D75tdaOpmykNUhETUT/NCpPruNj1Fy1JgOLha3vekwDq6u5/JjzwAfC5uZjJZQr4V9V
BAxs3N8W7YrMZMpYtm6TJaV8ZJOG9yOIg1tUJbrl57VTa6yTKs7lxMbc9Ygo9qES78lmjALvpaxc
YFKrGovkc1tVzQisDbNp7s840HUW7a9SddJ+DbT7Zt6F5zEBFvFz79uKSVu9Go32C9LK3IqDSEwP
Gnr7EnuUwcVIAe/c+cPoraWuc7AGP8Da1PzmlQ/ugu48cyiRoZgx1+5xY1nnLD6k6224leinMXD6
5f0IxW+9BHF5E97wz2h1oSU59GV09R9oZC2jQFQsUBKL1HbdYWEwYIy+GxI260NSGbA6Pk1eNhKh
g+tRWE/1hv7tYgTyEDkzaMMZG+R7d79eGoBXc47nC+vF/TeCtq10YukFLVSAC23HCG88QvRS62h6
plOFQr4d3cp5r5ooLg5ndKcs1EVUbNZKReADiZ7f6/wCCpgDyzOrc16hoHfXjwfXJTJ7MWreA9DS
E8M03Ouu6liX9s3no+H8JrrrlSs/9gLQU+qc5bPrrLZxOr0GHl8/2e/8feNqEbBmRtWMn5XvjJ53
HU+pvIadqmW39Q+nnR/Hbq8tuB3W91JMgKrPMSyypMv7U3WuAdTo4pHtwcupyF/PpibNDO+XMhlU
Q+TiOsEVexMylhj8YKtQ8FTAlw4V5KHW/z+8kMOUvpSbGaAgyr6ry13MsZQtd5U9Xcu/iqnanNfM
951OnS2+FYMlsOP+9pQQBqXaDmFaUahcBcmStziRSfM1zAKKiyxU4cDwobvCM+M9pl2eBdtZX+hk
IHk781PqztJ3wObZx3V7t7GL4Nj2qnCYCXiSYxDLLZvLNIvb68+17Qb9ax6p3qk0UW+viF2Cyoqx
HDgaylpeFLf21ZxEeJ8OmfhRg8UXLfzQ3arE8lcrP+XKifvQ1yTe8UzXrZw2MfiuxNStd8KzdtAx
wQyqR1dbXvSo5SzMwcmTKp0o6n9onBkZHNT5XLNURqjiPyM5bTXrw6fenIhfIIvqI3nUugbUTSI1
TfygAAIEG7TDauVbv1y46y3waJCE9YpFdutmghFJ6hPAY6euFFI7dsB6tSX89IR4a8FWpHe48ZY9
ruImVmWCEyvm/0LzjuJJEmrz3/8gt1SJWbmhI9ADJJ3ih/IchiiquqVUCwKLM8YTYAhL6XR77Rpw
vjZ7wc3OYh+RZQfObMP8rygpTOzJS3TiV5rYmTA53ebU7rvywwIryUK1QBg0zPYWWYRLPe3jLPWH
iiA2ocARsTqTLOUuLaH5qoRJlHpMF7vrYHLjDQ+1A5PDFtiMTf4keYy5OyJu/a02GsAe5vLpEW/I
TQ14FAye5IRsSB1k520GNAru54bYhYn8yzO3H/+iRuyzOIJBAe9TsctQ7VGI+Mfu1hSYms4w8rD7
tlgc+PQzt9SUvrpkRuZIRSoMaxZnUaO3BfMFG+mtPB9hNyhnQ06p6yWdT0MPCGrMjDW3It5CJZbq
rLgSMfex8kcaPqnU0c6VPRVY12huxZ/AeZJNfGiztR7HKErdexPjMUrrJChtzoHen0Bjfg5etTfo
jHSmLKxINdpoNjSSeFaAvC/4oItPcOzWOUuDYAwxbd25bUMBnjtRt/L5/DmXiEihuThVZy/Vyry/
4EP1uvox+h0SjoNWQJzr96D+06VvzkfzM4EA2j6LOHEC7rqLdi/RLoTKUh4+LqSPj9ud0Y3RPKZP
YHbt5AIi7G/IesmN3XMOql5nf4vRFizbrXDHknwf2sKXu49igETi7rqD2U5/JCXIl0sDiyZKq00u
4R0Bdnq+B25QKIGNk4vkrx+OLGc/MINr+QOEHEPaTVKfox+Xa2fMqDCbaxmN3xJ9N42c18fX5tSY
zEn3sKrv973YFFCAD9WZ7u7uBa8X/Bou1Un2RzND09uw2e2jzQ8fGhrj5CRrZZH+XNxE/Z0RYTYw
ntSvZEpGvZsv3zUZ9nqHil9LZg9Z47giEPbNl7eXDjNpO7PnYYeGGrWUokZmfUdvQagqOdbv870L
yrkorhvr+i4mt6GP98pDX8Uwnl1i+DgrQQY53vwg2EvAYcrprR0xF3HoxBzU7mXvW2QBdtZepRRq
Mnd8A4Y0EuYl6B90xkghPy1Oq7gPS0XZEVXHen1eb+WmrgKrG2INtnUDUurqJIvA6e/iIuD50HCW
YEB5IxQ2rCw4cq6CYbZI9en0kZWv6s5DFLFU2sCC5pc0E9nsNXX2lKhuvCSGbWP/4Vx08D9k8rbd
PLFyPuuVETkLa7h8B2ZLJx8FxcZgM7QPInJpkof5hd46A0E4SlenLw9IYG95uVn95mida4q5Up7f
TZGFmGswA5XYEGwTNr6dDh2dBVRPeCOxVG0mZSg7rqlLrdSt7U1GqHSglXqzdS/SJ/x9zm3B9yUr
OdhOjcjXYJEuwM/nHPYJ4HHpYq5cIrVKmTqQewnsUmJ7Jp5YA3yMa/4XKqQCCRPDjlu9XbPwKPQ4
Uzp6tEBrzarF7L7mw050CxBkKIMY0EH3sgHJf/sqqc7Y3cqz4KkoM6pEDvH3KwBTDXREEb7SJGqh
lnUiWpv7LPlz8z23rSs8eY+3wMu8MelDjELlApI+R9B3e1vV4nYTTJjvtlbnsFfbmQgbHg71F+89
2vck3GmZrBpnlDofOsG6Kew1TrAvE5KuLPehxv9/FaaMUBqu3HE9m/malIq0QZs++XCI2KJ8nQXl
zDA85TH8M42imErzCek7+Ujk24qZa8hwkNZPbhRjIacN+JvZ1BLqc8TcIqqd9xe5Er6QaPD3Rt0Z
y7Zjme/5SsI+zPyUbLjRQbc03YGK4MoGIAuckWuFd0UYd/lKa+s0+EYY5X6ru9qhgMtBsjdbIWAg
9D9OcNIkxtfEDqXqmNYVZuclT+w616WDT7Gaw1ewwcqg+tZWThWKoFVl34gO3rIiiRcANOZNnjvy
4X7l6KCFN1BL6bXqu1wAbOP0tdS40A3/XJ6p4fDckSFx0FVoMQEeo0MCktrJXK9GilwdhzLRkDsU
1LxgghfNbIXGKBwg4Flw9H4EoJ6Y5tRBwC0NVmYLXKu0HOnxwQVgjmyspOjzIgr5D0ZCymEe5m9i
rtnWtCNAW4UdeTj2M4q+TUhiVb+8fU7RgOzsylFqf5mJv7wwCITNvMh7min37CB5OnGVPnGvsqgF
o737Ec2SXVlQ+mrvtb/hJII7Pub+yGtTTzKc0mFBw1sY+OPubnsIpVMah1MQN6Z7adGuRZVDvWkK
Mr+Bjf83FB7q4OtOpdGZKlhmrDQe+3fRFmFGQZP8yg7+csx9tm/g8X73CX5lXn1DmGG6/H+JR6Fx
uk8EcwLXl3S5wTWepBrZLX8JxLtISwR17E7eoGrE8xER+2fxsr+D9oO+wU4IerDcVhAsczoa5H9j
VwJAUsuE+kkj39oz6YqxCtT4+MGXFgv2WabqUKDoP86Evy34OL51fRfJ0sqKmd/xegeheCZmbiD+
b14rXyZ1SFqFhnKKCOqTGXIhwZ5wNiqZH8pAHxkVHcIt49J2DuacjfICty6hT01XUGsa6NW0+/ur
kK+/GorpYpZp45zceI0t1H0aqd3WYJqcvGVod4JUsnBsvmCHFbCsiLfWaNAewDU5LNpgux+vMxlt
mS4nA4Dh8Im9hD6vcxv9yPqw/kyNRHoHCJH/7NkG4imHGkv0HGPAs/rOsPQwwjAcwGA8WX5Ul0iy
TwgSoC5kb+vXnDeJcKQiz0a/jx/BX77jHQWoLQUlR8GoI8e6o7E77wsVCsgAJfc9v8M6krX3NA/2
NaFhTHPr6sshBBJlqlEtaeWXabl31nL0IVbPKnA9XlsYxBwi9xuXQz0mBwHeusHD3St8m1BTds4u
hJIXqPmiR0/GMpb7L9rM4mRWAvqutLey3+017yKpHtwz+qP9D4NrsuOdP3kIYG44YJfJNZE/hLDh
8efLE63hiWt1KaJ4l70Rnyx0K1KGx7wag8P8iZZ1IIW8YyIJzjL+v87W9ppWHec5hz4LY/teuG12
y9YNoiwtd6feQH1XQ89a2gkI4Uo42zW9tDZX4G0K9cICQoApV4TrMuBAG7AvImY80wld6P0RIjLo
yKSYFrABdjM9C8vrkTpX8iuqjpAufuOsvB4hvHpjhTpbWibvqmwH1/Tu2o7e1RzbtIZ/JXECz0+P
BZPXG07YrCuVUH9rfrNjhbLAzMdMstlsDtTykOaH8YMDmi3l2XaPmdnCNGbBwNAJGF6AdbZtcc7M
DnM4bg//bIQc0Avy+WNFrN3624WZz0UVfdLGTUjdYTILBjSteULYKZ3PFugcUHA1EI7IxyePGO3m
NObhz5Vkq4yyTy9digNDDkhESb5NRTBI7qaStkBxKszlkNzc9BoGo70PyA0kyXE5EBnocJD0erqe
ay5S6Sl7YesjL+SrxoMLjx/3PI68Ny3dogUmoEiOwBdrN6lfdQ+aI5iqXBIblgbRAdzpTCpN3s8s
7KlaDizdqy+O/nmAPNoaTuydLUmusHMxKopYDCptvr8IkFTDB4JuVGDrt1k8HQ6/6n0ogg5kpl7U
2+xYZRsI28P85jZZN4ehsk7cBZFZC2lId5KLacJi8142T/AElKV+dTVU/+Ch2plK3oyOEZwi11AZ
8ezl0/5NV3FOsuoEhHlR/5ZSM/gw5G1ljV84o+FjWyrcahMwup/Rjf6Lt0TQkUXulAmeLY4osjdc
08qoWG+6nICYKL5b+bjn8RiL1ALVh+Pr6fBQoMY1hyzMsLEdgBPx9GaaJC8gcqqdzKqzDjPFHLwe
JAFreik4gztR1ymIAWyN5IocE8gImjREtXBhNSFwIF3/4hWcfEIwqoAv58F7n1m7aqb95i3+wyMp
pYu/QJXv+AXQXPRSRm08wrZN6KjHI+JWG0b1vTFYmSp4Xw3l6LNvrGJ8jzYBDf8tayEutuhavaVG
rJ7vFkgzHmprG+SzokY3WiATBftXeODB6nqWwo3+7LX1vENccF0zN/JrBphx3hji7lhYUvBTjS9W
V/wamMtFt2W1JhUhaOTocZn7/4fmJN2StcjTS5b1YdCXMfnhE5KJSm4oednl6VHovsFXn5xFJsF+
um1L37PIum3P7fIrYx4zXIy4ncHt2MWsjioI8lbbvd/dloVzelBrK4lUSAM0E6gd08BKbxIn0EDi
R/jdqjS9+WVw4xTbyBUCIBTAttivIbgqCrJdC1pd0NmfNKI0Qc1vUh51tX5k/UC5b6ngkle48Hi9
elWzRDnMMoGHBDUakEdR+vtoAyGEEDs+5Bb0lhKgo6UIkB8Wd3dr5msb4Bro4YCBHc3xP5Wi638D
NoAJJf4mKeEwzdBQ1dkCL7wbo9vPiRMiXEgka2iZMfaPPhKxmklvq/ozCQUqP9cmg0K8WVoQXbta
DgEJBCJevS0FqicFIRfLobJrk/wjopqG0vPev2KnOM2V7SRp1jZbDLRjEylBoWVQEzibV/SyEW95
lmMnY9h33wEOGg5TOoUJ35oSq6FNb5P5BfOdm1u0NsyeFeQ0nm48ZVl0m51PYsua6d1giZ93AUEZ
V6B56zsFaDhgvRMae8XmjCCCvXESH7OJ57J9MLzs8ex11fGhav/EqVbnJWPc2zvNhSJNPawOQdVX
gHVq7zZu/EDHtT8mZf0Rxp/lZm2955GiEtZRRLHk59KYgr1c+s60gNVvcuMJ5r08CpCh8SNit1d7
SearDcaAqq/9df9CJ8ritAHeLJ9TfziGUEtZ3GYyRlrpx4hACL+IT9RNvWzQBy2uxdW8/kjIhFdq
5YJdxcQJ/TZhQn3OQFz8cqwlIyk3/j/08xeOc9H1wdjV6gOuYsPyXBDeBSmkHEWWFcuHZo3HMKli
prPN/FdAOyEm0pxwdxbH4zNLQiykIH3y8OxC8llPfpODC3K2BUmTs/sKhcRnx1JZCKgI+tg0PHG8
dQDkTt0P3jgUllwy1QSnyVwjput7vYZf2F0UUwYBk7GQgAqo679hMr7FB8YuDruuTOsmNoear+tf
kTLL2F+mXpV3wfw4CmkaPfwodg3ISdu8j3T2iKhymLUFWb0Q/b8U0SxgSFm338pnk6zm7iPsTV/H
TzF4vfrpTS1VRS9UGwWvu51ko50vLPtxjKU4IPXnqsAQ74j37OJe0IrdvdOM6e9F61k/4Mq+O0ri
cUOQevKTJKjXWts0wSJX7hINinvvFB6soycqwer/3sRMpjxiLoXS4LQfUi9kwv5MBCeZ0PyAUXPA
QbTMT74e29ZwSGmIzqh4RP2EId59kBth1iC2MX0uAOK+PraUFBKJgZTMKnhNtVu/RJ4EJoAxH9TS
nhUce1+YFHviQiUJLCiVwqOxifckFohp7fRML2T76Dp3wvBeVC1H8KKSxa6h2TpvvxkAu4wk1jLj
S3D+Z/kcyAGN/E1YkY4RfHuL6hVy1NwdtMFjhJilmWjt5+/z/ifBXFyKxoiv4pUy5llsORG+sDz6
Z7mORK2QsLeqx9NgSLfRG9AdZF+RUPgSW1sBINeTRxrxjsQx7QvL1smobuJeNMqvMgVDLR8FDz1V
rPxvv/dGyxzO7y5Nk1hGxK6aX7p9OGfly+aMFAETiZd+y5j6yC5Iqrrk3v8qxZjl0Aob3dOQgRKJ
7x956pUvmyoRJoGQjqVtNo5Rlw/1NlVc+lE+0JDk9NOaxZKVilrxj8vYExyxm7WR6S9onRnRAl7W
9CYG5iAol+/NRgpx4CQE09oiZK/kg98yXt4f0ERajBSaC6dj6ZwwaM/n0sWhMN6ydMdiZjtf4/+K
DoIoW2dvvsrMAGLAnrfbQq+r0GcL9SBYySgM0lVMyCMTP+lPOgODlOk99kGMJqPYfHBY6evLwFY9
7L+Z/VQcIeobj5eUnonU9WSmyHASayWAGDAtNgcp2b+NaEdBwt3aoTbz7JQ+atNlEtpCUY3VbSgz
Ir+zs8pPleLK827MXecCR7ivGK+Q/OyZ69yTo/h3KPZ8jt3yWx6JB2trSnC7LAPerakCrAIvP/nL
/6K+zTG+3WFGSysYuxYOOTEQTNaLIxAK0IRwo+Kh7XX/d8TR0VH6s1ed2eZEsug+b2uzfCyIoxqI
VFuiOI6KY4O798ghuJfadWboNp4gEoFrqW9CxpSfNQwGADeSz8cdiskKp88wKFEQFBrrmZueNmD5
Ep/D7ndJZX63ZbHk2SK0YMdqh6/YD9Pd+oLNxuv6VTHPRCqaDBURvGjLAQSzoopCFsNhBZaGn+ps
MaX0rufLJuLjw+cGGM2pBuRBIRzu6O4dCXkzXFSY3SsfyqA62gosd9TqwtX3TwYuaIJkB1xRtq3V
E5PKT0p3AQY8s08pwAbp3W6OJ4GVTkEqXM7zmula4A9j4qFR2h7Fye6q4i2Mq3DAnwOwBXYYXKXY
DZ6gl+tUEOpc8f8OWZjzM4vKOxZZlijeejW4fKynXe3e8wIvH5ss7fHwuDIXyQ813ao3tp6KWN1Y
0A6HTl+XCgwvBeVC3fO6q6AFsESWDqhma7AJZPlD8NaFSPe/s7tpOZNefHSMGuACd0fOzkWKnqRR
212sfodbwGwDldTzxxB8pfALQdArn87DWanzV09AbdOhXV5jVWuBc1IXxm2ZBxUU6jn5Gsu4QdYb
3ly+uyrqqWrhTmDpBlZtnkWwTKuVv4IGckmU81MOOsaJPoc2wvqbl0E/HVqdJcE6dxc4diszlMgG
mZ6Z1kQPjNsYNeetC86cMB6LeX1iW8HyiPhEjtBSfWjouOiVXUcgIbc1mpcl77fnszGVxkJAzO8u
UW8ohWCh6zkCBO6AfObqt/iHYbYecUKmdpMGoIdMbiAG7fXKMUXqFjQ4cULSAIEgKfr+TUQTGhgb
5L0hToVsjz1qfiv334l+42fRMP5bxj+hbBvdJeUE4EnYbcDbDgqfyaKjrv2ttg3U1i4tIFbxAPBY
w1vMZAcvgB259Lzn1P4a5CFLdhDMMBBzQQEJmizZS0elu+cNyqCGIykXNRwntqHvgMyYL09X+lzg
19MgkKMmsLLDn/CDGevMkegdDqZwZ5OPmeSCRYtGALjTNxFbQ7w2Eoy8KzOi1jflOeFUzYhcUrik
ZP6R3dnhRsOD+ga/lQxbgAgw9aKUxaXTBLgtamjbnoZ1enczpp5DBKSQXY5rzK5sBYCi4h4GKpe9
Cg2Nle0ovoRN5pKBLYoylDtJ+ZT7PzeBdS1UMyhg8F+LQDXh2kx+dbeq+QClZIJRnQrG7ys0/2Pq
EDKfWWdOk9hxjDxJEdsbwgjwp/ry3iFEX2Y3IJQw5r81atLZY2omCpADeZBaTT4jnFKdgKMMuEvf
gOXLEusKC3AP9IbJE3ZnscqgNsAgjVU75KzHpK5VsAyn4oNIl276RXJ/2NMQi3ArsfHLpu10Wh/8
hjFxfMgLz6hGeRv/h/Z1JsA7r3pyvYJidK/KkEx4DtV85gGNCZFEEWkJ9OrxCr2HeeuLE/aQ0NYk
zZ02t9whL5zH0l+d8rnwgpI2wBo3DzDtuLCwLvq3EWDDeADLucu16lUvDKycwb+BcO4z0Qtzfxny
PyWueQU2EU+YJZg6bfxiKiF6KRKv8iwZpaaCDaY4FJURjy2rMRM8NUCHYzAHQD74k88XBgbJ4g/p
voB9omPodwu+y2ABGQwCzaTXgBWh6gMpvFCTYa2N998TpesSU43CN6U/H1Wz3baUK+0Idc2Q3e8D
VHtGWfG0nK1J7koZR+1vnxC4UBQlHImD3ILz3OkKm5pVF4D/qteYqEH+bj4294wRGPZE5652vr3T
6hc/j6Ksn1LtZ4PnjIYPf4z1oWNLm9SUaLTbSVhFA2+0R7i0SpMAfX/Pe3C+IAI7j+NLRzEKiMnx
VDAX5FeExAVrVK833bMZAlnqvqsLTtmRuJtPuuDTJ/9mjPNrmHDmzEKcskrvy/Fg6EWdVnzGB5al
4KnWze/GCWe98w8rDf29Q+dLf6WL/x9yl1MXE7b2mX8EFW6HOjkTpfGJ1OeEj04Q80Cyabu0mTjQ
eqtARuafYXZoWR9/HQh6urrEJZYJNsJEWQcB/CL4LAiY8njJ47Mlf1P1ngxdPSENIG/1unHA1dk7
aL9+p2ZLSQAAkbaRcoKQ4uUiA+UZ5RliR3UKh3pYOdyfpKFzOq/XSO3KY5ppTgU+ezLukGmRpQAw
Fveisi/MlZHhzBmIqR8KJUfQ1Szz2UPVv5dBTvtQABbJqf+0UsYSLkqgBs1UuyZWlujHdsncXEzY
vZpKh44a91YBVFVmtJ8AGhWqAmM75I04Z7y6RYT7+OVp2BLVEGA/x5ElK9pdtJTpULjZVTbNctkk
i1GnZ33B7rnIbcMp5d8UlvvVBsdQQe4vurGVkwcWIFX+7Cy3Tp9Ci33SepnMn8bqloogCHo0ytln
rRYUecgrr/qmFG7H2kPxe6dioj8WbWyYtGfQIdDDAoj31GEgNwE9A67jX5C7Hk1fEtFYUOYU7I5N
2iQQJJxZ6T1qot0NdKJsOfAOz62kA2W0MsxZ9aXm40rQXGOmiVbOuB+DXXM+oivH37ryvEwbv4z9
RdRnN+w1uHQH3Wkli4ezKfzhgAnvIsgBCETsqLHBuGKw6QxLSRha4E5A5ar6Vq/0FWugxPVpxdPU
98KoZwA5Wnyzsua/KjkDoXxyHDH+ikcX3zLpPtqeGSTV0YDVdPLrQIC74gHdNGO+mzMGDDTdfknW
rbuZehRIPAOYmop/eHfL8jNZ5pQsULtc9qLbBF/+vsbM0sBIJdzwn9e2z5khMtBOsidsNoLgO8I+
+CBfQ0QLm5cP1EZv00pHTGI0NQiHoUdVW2tGczW6j+dH5UW2YyZdxVWMlOdh7axYDZNRPH6SIk7P
900IBG0zfhFAnULkmfYijrZzwFovqrKxdQ5sFmT+DTg0hcs7cGVI8Wwg0g0yfNmsVXNmz3n2BqUZ
3NP4oA7gLxJ2dK6ttB6CLMDC3Moad2xgCTgw/7kMHGXIPE99ml1As7TKrRUg6jb4nVi9rWxTPRYH
uSXRlQjaIOBfmx7lcOAVlmEu1ghGfrI3omQnRs8BdJxTRAhZs6f1WyShO+oYnXmGo9DMsQ3t64Rr
U/SYhjv+wFLMWi4n3E+NRn9Q5Q0KuMvO+9K0EjXZSiHsz16Y0BuLFJ5OQoez6qOG3KT23iK0oyC5
1To6N1sV5stFPw0lMSi9sjvsi50KTcgL06XfTY9Ci9jrjurL4cV0Ibb/gfZ2XQ7AyKs+4yBwT2Rm
ExxUetrFA+fGHICP/RSmEckaM2DWiOiDFYehHulvi5dwVhPlqcUavRMGDMCKTWftROtrVBr7CYjV
vOhuGVGdAEto9yaD3bPzUtcJRHiHfiFxksyHlIJIB78aS8YA4gzBIK45uBX4hZbD97X+tP1TMcyz
wf76mbRppmmUH0FyvKCuqfr9Q+jJv5+HYXrtfAgx4//1jyFE9gYLC8gQE6pDGRaR4rBxnnD9xbZR
TjkSKGlduqbPbb5dT7vgtXNGkEekk6u0skKmRh7sgjnw7Io0rEK982F3jEdBhgpWVgplD3koeqdx
ia+DFZIExQVXiBD09Cp3VlLi31n9Othb67c1GAIiq+jc4H0hcUMPup+LsTtZ5zYocE//dCLeMGZc
Y6EMcu/udBqG1DS1n1qzcRkWORcasV0dWd3PzVjE4L4p4Zzo3kQIf4MAnY4CvseydM2sLEBQrKJs
wAW8s+DchxEApSciqcBGPGZp23U6wyNShCk+zWN8fbptNpT8EjEBfi5+ciGYdSB11KeIiv5mQXVu
+qaGmj+SRsU49PHdE2+6/RsxjEeXQdWtDxbmUtLnYfDcHK5C+Q8EqTKFy5HlvXD46jUqEfUcCvfu
68oV0uhwMRtvN+0wawRQe0V0xKK2KaIo7NVird+TiRFL+NPWxaGTEU1oQE4YWHwP6ViYIl0A6fGd
24pJxgZ63N3O065c0pAxe1Ki2fYDlM4b4v+A15kPZv0OA/jAomK43u/QQXFhLym3mr1zx/WrmxEH
yu3uLVFCRFcg4Iu9GdOTupDCwjaXyny55JsB3HrYALcBg4MnuDow/PrkuHDz0kludlZgJnE0WXMJ
xkWYoZiUW30VAdUdxuJrboIXt6shKD98i7OTl/54BCAgjmA+Cz6yZrEASD+eF0USoXDWOpmBGKEh
KX/TmDdHkqF2DXSSL6vfPDWQeMPh4UH3hthnN8AgyKBDynukwL994GJ5BQMpaeULua7Dnwz7F/gU
MiAyOZ4DQnm+JBnY/xtiDZFprPAvDCQkY4CHcEuYVPG7h7qNA2GskfWl4wzywplrditvfLYs/RVq
VwnpYsQgBLkCPd2+IT62q2qtC+zmvedxa5YXqaxTCb1dxbLVAvcy64fbuapQ8r5lfFgMBfmCFp6O
0h6F2/gfD+oH5sLWTLUWxhI8TT1NpCUPhKAoccqi7dsGD4g8FQnCpn0aTIH89oFPF/KLKQgGY4wY
pY7VwYW8GLhrv5gKHS/STGtD9nkQh2oajy7BHoJjFVCayzyBw68LzlMLoskQp8aG9Ity/6sucuwP
KD+n/km9BHLfV/jKLlEbICn7ejUDeCUbnAybahw1aH2uXi/R78bpQcPoLW9AD6g1iJfrZc/6pa0r
oHTTnhmlEe5OI2f4tXTGZaMaNS7ScEeShZX+FjVDu8DcseqjW8P2NrgzqoRWSdGjIV8JpIxvirjW
g4FWENKFOFJNX8Qb2zSTrgJlWI79jl2X+LJ6kbLdCnC+H7c94aqaw/+hIi0wr3LosR2iTmlQW5MM
9oDy+7NQRzODEV595VPz5P78PsJ7IULFKCu4R9JkGiycuEJ8axHDWhnilPaTbvkS6AxoqHkhpQbv
ZtSDyHHROUBO303xy/gKTNQ8tDUkl0kOGY1cLWXY2tqHHB7bOtG1kbZNaBlsKZGmPv7u+4ysNC14
P/S5QjsnFNhGqoAUnONs+qC8Ta6UUObzTzMcBlWRWygcKYQsiUspXSroUriy66qxE8NfvgOGEGwp
UOBriFu/sT6kRmlVgcS9smvw/n81t5sd67vYx9+XuD1KE8SNoJazFKueSYD9EBfHufxuCSGbnvzh
lQvIaP3VvTBoi7byoIIU2Ti5mRkdHOCB5318QB8+/D58deIfNY9xndS41VG8obB1Dr46hetyuYlk
zfBxk2c8FmmoCXbkKwfEFe728yKymgtbe679FBk3qQabLtJoqkl4aPl5hZQyqKN4D5x5O6GeApYg
ZPLbVTy55ZksTF8VtVNJfBx2H0PfwKaeKadERIKYKyK80Bm6OE4hW9FfFHkmY1eg0nRan7CYENSV
P8z5pIuwm6UnmCZnW4jaOfpU9J4VldPs1BY+QarSCrQ55wwwN8AZh/0TItgcNRSJRW2MZjcgXObF
dY7ZxKwG2F23N8OimucEOsQ3hNqGH9FC2TbupAhEu2P+jYR5EVq4Da0P8/cTUgL6y0dOfmOiV02A
CFFuHHllk1onPCrXbUKHF9EmwJEq+yXaw4GOypFs29XKW9N/V7Y7V16UHipU2ap7E3cCmPzDqLIq
Z1bIuwbJXMxiBlMxDbRX+eCj3M+nmELZ92RCc9Pe2wu/L91xmSc7A6hvRz1Y+OK5NPTCqwsrJjGB
jFNNu62UommQhHWMpEH9lHgBwcUGrhLSCuhN3Ymde4qdK5GLt2sUrJdE6PAdgcusl+cZG9p3Nytz
aXKh/h/W6BUFx807xp1S86v6yrpL7aefwoYFm4MOxcqVqqMIx0CTkpF3ZvFAtBhZeLWtOZ/BHUPq
8SYxuNN35kezNvsnAp146iffzVgR7Jurn+/smRN2YqvdKUN3j8xXipEKdVifpbyV4cyNvWBesl/v
nkGDcJRp3Y26gh1SAO5PvC0qmdci9y+0pnWvtZh+OQNPlWEng4fjCQR3cc89BRWdEUMdmwAXSXmb
K6wDXtglqIRCeIGiBLqUUcYGYcsEGeAWpoxYfe0qOozUSSy/EtKhiWR9g/6vn1TIo05bN3wg91H1
f4SwzrrEAc5R8BjAHpFoGH9sXW88ESNNM8rvKG7FzEy/Jvs5JIaUSBFgm3Cy3nmnar8IrGTsZjQW
a6Ur5jOGjscPMEDy23oKJnDvCRn+Bq8KFB0+5b22HwdaoKSqaH6i1pxSC/5aoxcVDmsh2RU8yhz3
itmVxyGnoQQ1r1llz3+espZox/Q1AFzBdc0Bih+AQltTcuJ3RFwY1PcBLdF9kjRbhtvpQOF828yD
gTvaffmFi68QtKbP52rOx0Qt24mpuRgr0cmIzCXJSEzyjo+kOMpe8/JvqHFZmd5O0ZjyuNC3GxNE
9VzUT3fX+Sety0DZPwr6icexoN3gfuzKIRtmNloo/E3hqb0v5Xn2RAbmKHoIiv/59wc3jEwulCKa
c75iUpHt3dA1SE+YhtKiXszTsF7b0Hjtn/sypnWF8OMrfORIWRcG8xIUiX4ci9SA/uqmnGdUDAjS
mRQNE6DzrCV6QOEmjMWd1r64ZsBFbqSCHCfKzkCwiNdHwRM3IB/dZNzxJYuig736kFf/ZIqCRef5
xk1fy1pOwGedCHTRdnrM/4NQqpOOUtA+MITgxYpcfNsEMcmZMTaj16Cgwf3l0rDZUWHd6EwlCj+x
MzfKx41vBf2p20lz+tSBWiWy3v0gU22QzhOn8DwfVFKr/7/lGq828MrOBemJo69MNQN1y05YTQT9
hxqamGegY0ieRzdVqONs9l0mRAFrzRaR6vOnfLNOhWFoz4ygb/cWGXfRj0SPhd86ovP7/yrOexdC
5we6MQOZzptG4CKB23ip7XiJih5kB48vztEcrQW4aQMNWp3Ei2qoumroZhj24Ec1CU3Fh8YM+LOJ
Pteedm3nNmSG3H0OjvWxbMzSb6kHFHnCUHFBfGIrPGnbB1xUAOYpFk+SByM3P74IwWJ14L+6F6Ne
BAhFxxhG6bJj2NQKxaNuie38gd/2/tiS2IfACW5yOPisuFfJcPNwIcGNRnPxUa0A2d3zSFeQH8og
SrpE5q33ik0Cdi2i8ieAbAjiK4JLfR17eJ8daT/cpo7moO0jEXMOOOB2yhmvFQTLmSnxUc4NvTYd
aMAEzZ62Eu2fVTwaQ5HHYn6yqAmvP9jSiPvs5An2d4ANVy1g+poYgj6f/KIMDK9mKSYTi/2R0gIU
kETdTqfk6jGt789WTCDT6ZmbqovTHhUCRqMbdGfFnaX4/70ed05WK5WEReI19/19ZiofSGeC/a52
ocqzlBU4b/G+a7f0G7aql1xDCyPu6Fx2mAYpZ7SRbKob+Atc1M9nPGLuKd1Fvi6nbk3jMKTBrEjx
yVlVCFqUK8zaXN1lB7IItOmSPETv3AeZ1Ubrv/ICO+SGXSak7DmTGtcDKAtoApt0AsKyGpqhM04E
Aw/ofyF9+uRJTpQQl5SNZTljB5xkPImebUMkc2sRZgyN3WWfFrLo0JZAoYVDb1iRvU7VD7SUlnQp
Yzaz+pesltNC1l3KJlqPromsVxJ748u3J2Ab9yjJFnSVY81Fk4WXxVMfxpEgs6FVfDTR06oqZ6Cv
Y9RUdmZ1JPZ/64vWPNoHvGfjVSnWctxg/C7OqH4JrI0t2q4ua80TlLONgGlDyTx7xaitYsaALmO7
vyPBZgRnsl65ULop0SJRjgNaanZx0+SLmSmWk4j+aQ9UFPO594v9kZ78tMBaxndUyhy7x7DsIYA4
X/ZK+3s8xCCnqamYFXtS+gRt6/wRJuviXjjKN7+g/CesDDhXV+FezOYbs7WbqqqtVqdxZXo1rb7S
7Dj7/ig0/eeK9BCsAqk+Lma5OREiD7cvRJFiFcu+hzap05t9fau7bcTKgC34ZF4XEFHoxY7TYWmU
ykY4tnPzae0mvQHW+ThFO0RnVSmF10Ggeyy63KFdprFtOBeG00bVXR9n/IRMANCThd4yztFYmmfs
QQ1hu7FwcEXSn31nSXhls2An8ZBSSo7sSPCobSAFwrBa5ewtOsyjr4TMQpGImRTFIrFuKKHr8Wgq
RcVipUhaOFXfEjV6WJjugtU/Sc+rDwqaWMGhgnkFdqBbTZxguS+ZHWCMMewAHg2cUcU2SEv1dQpn
msCXVnlUCgZrgK52yFROgFiXcD3n8E8fk3j91XTRICKDV8qcjcY93BgpgtNENrUHW2eTOYkxSgj5
DZLriq5uSbo/E6ElZ4LefA7vRX0Frg7RUKzVFUyqlysF6nTuKlAtLCoqWTn/eG0sKQy3YUIo2E34
JFQqerprymwuqWGdvwp2Z8CW62p3Ajoj2vKAun70XSMC7sI18bmthY+oHK6QuKfFUfufUqFpmeqc
dd4F9Ub6k01ORrRG22wfSEQdFCPvgB81e91YhYK+NyaxCfOPW7eFjI5CB35qdLwpR/0OOJej9dev
KSG5vD6ANRriSPRKupfO1am3kon9PxOhVaWgbcclPF77Ip0HOm6hB0DAUVF9ugfzHc/IyXCif8rX
NkTlrkwq95M5TAPrNgIoE5U/4OdbdBQpOEzAKVz2AHbElLHlsHHcs0yVEfs6W7OgfWW3twFR+KEE
6YlrnN1iZunquwm09lVRKVaHsqygNGPo8B0wiYOoMuqnMrAhg8wR/CrMObfSiMnC5fo6HpUfZbHA
/lqLv6n3JDXtKmUQonYmGabUIbWot90iv8AiFUUzaT7X/lbNWasEXx7YfRj3bICHDCPYSLMrPGeN
fm9nNNpSpqZim8lNGwqTHB4DV8dmzKPosn+j193rbfIwcDCseZCtULQZSj+l7t+NkHmn/C+Kcvch
AswV18Qm3CWDuD2bKb+Oh7v1Z8/RT0a3VhyhkBOuOlUl13wXoXuAXcedAeJMm6n93bO5KcHu+XXy
HLox2cbzqTfbCoXlVxVxcbHXiMBtbtWjzUxNk3eQW3BVb5VQsjHXPQ8LB8wndlECwngmZC5Amj7K
rG19PQ5nqH0BQusR8j6D5lEP9F5tPBC4JNErERj4r0nTkSZoXbLurFemfdpnl1K7jdkUtq896WRV
s5IwbgJCnmvj4LYTRnnm+PF1uN935dPqYJkq0ZUxny+9WfwCQUXKbEJsIxyYqWLeNAF7G/37TlxJ
NT4eo5B2Lnpa3sU2PFulF0/RKmqNWcbwasDnU04zw4zx7ME1dXuy1VlNSPcO3Hv7rbnm3VqcYUC+
y/BghyNe7YrnTkuiA1+4I8z1IOnniC+LGpr7qGBCXw/JL8t14oKykp9qxo9QUzm6wjaH9ziISaJE
gdIAHMXyX9TsJEuIjhv4OnCrLwlIy1j7FuoJn/QeoIbsqVJxwz7wEptMXnTBSv+xRtRAPKlZjD0Y
CA7neDys5+CDdbJP7NOaoU+5JIzYJO2+/1o0om36uTTWJcrW/1YuPHnT3pTUXx/xsy8BtWgYj8/j
4ak1iYsB4URSbjke/PhawNAdRTQWkvKpjrtl/TDXwwqtxof2M0R/te8zEDxH9nagJ6TldTOiNXUR
MDtR5vRr+LOV7ep5mSlioPlpPDqzoj7Cw00GgbuTGfOeNFKbwGa66S5uXJ7KkvFYi6o7Y9Dk7sh3
nNF5RW+9q/Nl9TQRDEa0pWFHn0ZN4robmAE6Gku2CAuV3XhldrgoZc4cHLr/EHHVl6RIvJoGgSf6
Ec5WmykQ6DYBnVHwuPGuLjxrg620636YR6V/B5lho/S5vnhf10sf8pTnFNVP7nFiZygM2rYebDHR
niHQO4muoxLbPH2oIzp/3MG+zaT0j3JeTd9fcoSrbvDHqWLKGtiJy6Zq/X8lJoirM8KF/waytK9X
K3GV2FiHUeY7/n8vk/8qlomDjiAa+9b6vMhbWpcnqQVmdoK2i/9ULQ/YlrqNT09JdHu7DobTXeMA
QZmKT/XMAUsE13BVuET7WthbE0dFEq4H9OMkPAg6T4JjXPt78p+1rg8i8sfL+gPtCQa16xtY+pZL
O78nIeoFrji7ikfK5mNH82G1gpZEl5UMVJJz4RtGgFFr4N9SZ9kDRoWhOOW7pSfs4tVqmGXBqpPE
d5yArZir89nlUDeUmVJvh8QHRVaHx9blvTnxgbEjoifktL7IuGeCL02iPGBciIdC2ZS7guiyEawI
gXeNHLup8pufuXqFCwUC7Y1dkyenscZfMKXY9PeVg4TwAJHJn8ARSRncF0dCyj92kfCZKgeoRaXx
FM3xiprmESsRh38jEoQTMNbUEzAyONBgySY+kf3QqwQae3i7B7PVSBrs4P42ysqGBKmV8Pqhc1xS
KaSMOklxeBlltA+Pr6vo1w6MxJ/87jSqV+TV7Z6puWW4ME0heG5RBq0vvuxxHCoMKovc+14hYr4u
IShFENA+LlewP0KKaepMoMIjR3sBVthjl9eGZ8PVGnSFWTDfegrkUz8RMtWhaAAF3cxWWUmiICn9
71K+rycAZ9hplmQpf2jFP6gpJMnO6UVljf01nI6LHvnman71VMdLjLc9rkbSJQPygoHdKF7M86tS
va5AzM8bkJKkAyTLEQk/f3vbzUOKQls1bbtoPNg8eAOTb/yAQaNZMuwQeqsKSbCm8fWeXr2CoKUd
FwuUaBhRcePYsci6e7+/h3Ps22qEBsrW8HmkXwm0kYDiewsTDR0Nuskd1K44TYK7awPvyXIZnO/M
nFAyi26PwZ36Nqfr6hxKHv2sKZ9k/4a002aQMxFp4RG3FW6uAjs0Z+yFXSH3HIAmKVAN5SJGd2lG
w98AMuMODdrDO7/IauD86yqx5+8GRCP7YqNKPM/kza3eJhFNFyBrI4aOJ/psmSH/zA9SRYVTvIpi
YyF0Z7yAF5VR8MymIZ1dvnQPE2jf32V8em4fQzPnKp2t9YwO6FQspXBFNp4NrdS4WPHeA12zBhrs
gex8dSSJrTcQIWq4xqUPEcov5u+EsUjQ2qSs6Pl/9n9hhEf+l5yAk8z/BhHgHhDSwUjzHstXZqvU
nFB8Q0Vf4UpuBTu2eieQCeBjAITlIHxHjOT3bwnODYlmThpyqZnbpPYIy0wXfC6MX5OSRDRe2a/l
wmUWTpWtyItPY1tkWzLjMdK6jGaINYLfOo8NmnLRYj/7kqy7JtqOOLuXSz1JaLWWxc+s7Bi28pBH
7AiJX+QwyaUjiZhQy3wWvxREwMzdwX2dHimELwY0Abeeg+TL4ItnlquiLmDfhbHoGIHySMU9MzLD
lIZGNs75zU0dZjuBbKuZ5Kw6ol9OiHZUNB5o73vZ+wULqYcvWh54Yf5ktFgWLoMj0MOD1G9trcDZ
JjPN+4XcOdXWC/rqiKXFY3aDzpY2FYejauzguFV1SjrBKF33nG1GCblv14hshr2iFOL8zIzFUTrP
rNG/mN4PbYYtt0E0nQyu40f4LpysA51VrQPKuLR8zkN/aUEkjriLkcfM3hThLdlZDkOYmIk0DubR
w+lox3srwgq4W+s0cCaRoztj66b4PMjsraGbrzNNDvwF9lVkqtpfHwhXteG7grh7BuA9gaMlAuab
xrhF2PiCw4QqTkU3BBWj5ewm/4DdundhnvPa5OZmX8RLDn6NuqoudK1baTK64mQzkW4dXW9us1ru
/2drX4l2ZyEuqd3fYMab6pLDgIXIMDio2Dm1wMRX5jClzLd27Q1vKyr9V5V2kyZotUk3AhoRs9BY
6BN718eLeFBwQ19zEfERoN+aK+en5NhsACDcmI04bmuepyFp06Byw3DF6NGBwPjqujBv7fyBpNKy
gzqzj1pLcRhakP0z2COEuD6fJjg1Msh2fao2eymcSlTH+/2KpYWGfszxIDHfYCc8yrOICRPP8QdN
DlK5Cgy1rP8zEsFX/Tq7c+GoCm/QXp+smESmOJNMnRHMXUpNS0uK6zkawIEUugxfMqfu4SvqnOaU
0SKUAsPVcCYCSZaxGEWpfKSJPFtVevq4uCey+f8oazKs4hz2HpzqNfMh5roPW17r/Sg8/1Rsf2Kz
eKLWaeOgmy2vIZMpYQeilSlpzuTFbWh6VolkmU5F9oA2F10W1rxlc5AGeDF+OuLGVKU32xVG6XHq
lfMPUNSW/PVSm8jsDKgCzSM1MXFtgT6kUrw/i5uJhM3Dx/I1AQRxRo3CJpy2zA5mJKvAHwVTd5uB
+rnoURFZd8VHqQ0qvJGkNHWdqz8LOLxmeKdmhYBfIGkl6ghW/PJ3IVQxS8Pct4Hyf866H7PN9PSw
CSgrwYsgcElTEd54TF3Ru3Yi2jtuPsEu1kl6c8ftVh6cfF5QE67fDzFXFPlB6Ztz7IMPoi+FfyCK
0EpRlsfB4z5/q17Uyv6u/37x42MP8HTSgQVS22xerz8EJhq9NnmO8tY2nYdGf5goO5w+kke23WPt
VtHsx67mJB3GfOh1PTEKmbkT8UBSPdxWxYrK69ogltkKGbZ4xoN5j4Rzd2y97VSV5lpxq1xwOxIV
h3lyoCZV+QQiHEovEiuSKW45Eop0nrLaEvWYYW0pmDKSnXUz6kSIpm5VWyjLemRq/doHIFTbQ807
316LpG9JFQQ/90yFKN2/qgQcD3/jsNGDcdsNGFz+lGH+RAVIBnRwRcbIPAG9ZjOD5XJZ0Nx9BL5m
1uDLIYZtze66JaxAmXNgahOU+AV0XrwHg1HkZTO+XGZKZkK7XtlefulZzx7ZIS3ZucQ4wfdcm2HK
eFfWQt7MwbmVCnUI4gU6+S8OB8aO9Ru+7SE9III473MBOqF0Eqj8erC7asbcurZWZtG45mEShzAl
yZ5fFOa/6hIC41qhyO5jsuF/NBamJiNgQpcHJsNTV2/ggHZIXlY/GhkeDJOJ/RS+Y3OjtEX0Wzbc
k9LYIhv1Q9SdUrOWYGjCD6okqNT246DoWjqPuRrD8oYiKZX8QLdWSYV//0fXNK4OgHA53RkFxtrq
HU+OCustOjKeDehrlp+k0t/LvWt1QYWnXCZlIGZVwQpIZfqYGx89I1ypnxrR/vWXU/bj0/LXo2fW
H5/vj9fEYriBQtzfZacGmVT6pbBl6EQvur8eKbVSXFRaNM3tYcRFnueE5OdfbkZcnFR1ipl6iFII
NvD4RScHibUO6tMV3IDLs3LklSjGHwM1csjG5n72Hm9jMmEAqYHxwfjK/Bv+DTR62bV33jHBSCQ7
UFm0sc0F8ICxgGmVKp6RRVl3hvErJKsJNBiU3KSnCOhCVzx1Kfjxbw6+x0/z7JrcdTRyuzGkIiUG
osJsO2g3cLyVm5YGQGL36oxfs954VYX7ObasSQDXguh/GNJ/dmJa4l7d/50vSADq1jNQEHd9afJa
ZEqVqzOSjIlzCDfVU4nTS1IUwCAXKZWvLjgQcb7fiKdCq3KbyyXkFFU67D3D3Z/6TxJg4iCt1JTf
pIfPBaOqTitWAnKQJbLO6jnSPyMDufn1RDfQkX0xSj5lznVIol/ezNtGVjwczVeZ6/JlPnBw//93
N55kRoMaBKka/AvSOXw818SCgyDHgtAoNthlKPE3M7wiyCf5XDUMtwEiXZbDoN2ck5E4gGos2ppv
iOiM89ctZQF8kraK69gf/gkgbXliyF4/rnJeFonmV0M5RnroKTeUNUAnVzeHzMSupwaRdik0X8dv
252xCp6RAleldlk81vW5F0bOvATa8ZQLYa7Wrl/5wjJHyIA/9y9Fvnj+M9NZa/YqwBjNq8WNVdWw
xykZSXj2fQes9mJii7ZdFsTWVAXJED6jPwfiLF7ceSfsYQiQxYZ6vcd90xY/6F1O2nmSP17GdaHm
r+P1fnDZhoWPnSSth6WuUuQC0HUG3K77W7jLXtHJxFyqx0XdmB2gFGpZB3czeBHPx7VaxY1hdltf
sZQu0MV6VUmw52oiRx16liwGMu/JlkF62CuM8YAE20ygBOA9Bz6D7KKyPmneV7EUKBBKFBo5Muc7
/u8XLr9Fmoqo83y27eTSxtu2K5cJkXd3VPLbXobMBkhmTqt+pV0hxG5bgV9JSGH4gyKoURwMj4PK
EK3tLCKbTlvKZR5ghKAHLgdsUnhh/8Gmi3R8B+iLxUyzqXIPYfWXkMpWeovBD/ZHLHov/onkEvAE
GkyBZy0M9lEAyKI2rQJkFeL5UVyrR3sUfq14uDIyU4dnGvv5vO8N9/Cfd/w/YjwTHKZAVgTztcd/
p19QszqoPFpb8gD7f83rx/b5RY3QpZIULuTpmz13kZGPFI+hMfZdXim73OVAr2Ysant9TNUfRjA9
WFyNglYs/JI2a5PWP0HcH0LIYlXva47EoikRQjClPU7Fi9Ke2OBgam7o/uYUWueIr22qUcWHoryL
YHnslNo4T6W+DwOET28FSy4vcxpnzFzAwJNBITahjHPx7QNFp6C0kXyouztI5mBDxPYOyKsDf/PH
t+BSHe2tuGnPKgBALEvmVmVxhnmwVNJibHY30Cy1AkSJS1va55kykEizOJjbj1CZgPs3xgLR7pBF
jLKEOTCuTtg+trfEPBlueYMrUMrApGQ91WnA030BfdTdy/u4DTKylPjdBf5u8mpMGYqUmuoTPaDK
dD5RF7xe98M5g3hchwJH/8d3/s2g+2UN7z9F8fD8vP89vxaIWt1aCwmKNs91X7imjvLBrVWRD8rQ
sHXUj7RdQU+51ZeWacz7awrzWjbeOyT8AHLKN+mHeYKPcexT2WvF8afB4Rg1Qq1jnFcCR1G6LdnV
W+fJRSMN8H1XGAj633Gaq0sNxPZf4Pp33xHNcUY/nak7sxjsXJBv6R84QKA3wsEPFx6uonBjHXFy
5wLQDb3vFUCsOnNW1RZ8M30qwq7KVb1o2zoTRA2qry6IQRoXkXehLzdt2iznjJBboAR8lQgoDgon
QD9p0juE2fdkJ8R08Dgypgm6BUY50SvJO8h3dJWsE5VFj8O8BpCdMV2hjuHD+B1jDz3mMt/ZBOPL
0Sn0efvn7ax7aXO7/Q1R0q51vrf5Fu+KxNmSgWcQOC0dgHyHu08/AC/TakwLyVxgLO1G7NUDqSr8
vj5nY0sxhzzg21/IFJKiRAxBuWyDzCan4uue3b9TA6IXbgKX0fgNRMcYF3gpgU1kbzuX7GRqVPTX
OCAa3nO1WuQQ7KxuJFGU9Cq5bl2khHwo1aHIiPYuW/gmGZYP/zoEwF+P3uoFPgv5bEsr5aeJkOyo
8qYzrtPIb72QR375800YEwnpl1V8XUIU8qjvZrtKvl1IFcxfxZMBGD9pzTtuTmkNvzW4esliC4MS
A5kArQ/eUp5VhBfnN+rkDfcBkiJwGp8VVmTaup2Y/mnhOkDjdifZvkAW3m4Koc1STUy1ed9t+yPX
fow94d++HBFheaR45RijZEYCymP8nP3CKLBoppQn0DGmY4MV6a/KikATMbzcn9dZ/sZu+QEyMGnq
Ve5q8xTl13aVxh8L/SWu3BtUB/JesdAzxANhyJeoV4T72dyXrDq5FoDdSRXLJkGISu5WiqJno7d8
sz8bgLGT3b53mPo549bvFhj9K/r4zSUtnvWh5jKWtsYabqJ2Ip066aKLyDYv6f16Cge1Ku6//LYM
+L3MLFYOCo5b64QvAhk3JHun9oYtgXY7gR9ivlP9yQfHEZ5vZRzMGEtPEyxw6bOExOQ+Z3pC0OYm
lzsTS5Bst8CYh3siNhCsY4qrSXi+C1MQVPM+kRjgY3Q3z0Loerr0wGoxslV8uughvSasFP3uGaZN
oYxqA+l8ZAOS1MQIOkWGfKOSQohL340PgWsQV6wWOaRYNmq6YlQLz2cDykcQyMKUVs2BoJdnQmNv
mLhJmNmer2Wwp2OL5t3kakiFizN0extK6cfF8NghDW/gSPmQ7mGPj7eME4TOPCTQcHM3dAgYib2u
NsuTFdf6v+lbun/q2iYqqBfK0+yjKZwBgn4leWsf7wVoAnJmVpUr2TLwqVKMgtweWChpSC+G51Mm
ISX4CUlntEfTeNgGVOhi35Kw4Mf/xDv0CRCF9Xpj3axNz71HShQngvRwQQ4iSlXSTXF4P8Yzl6EE
yX+w42TtGZzMAmgEKoeiyYkPRYj9A1IH/+CYvGMrDVjAHqdOTsSBBOCR5U+MS/FasnI3anpoXyIV
Mp/aYyp3okoS8ZJKIO5vxqQJeFJFm8CNSHxkOKwb85lDXbSVmBE/7S3L0ZkJ7p0cRbUoRKZVipiH
34IOnb5iteCFGU4V7MKFR4wcPLpfb0W4nkLzEjcfGDVV2fRCCYO9ZO5jHDjKsy914h0ZRYplsgoh
aftTs7CpTjxNp1/u40jKp9nitk9tLNajrgVmtVrBGF7rwlTFCXbIXHH/HQ4crFPXe5fwdQEnc3hD
wr4B9IA32+H3UTl7pRoxZFo7IPMZLz8WbknadIBEWLvReC76o+7gHADgudrIFYJgPqw4h6hl1Yzv
E1XaBCklXv5VooRck1Uq4546ecyWSdYyvwShH9biVgFsn2kuzfXpEzLT/jl6FR/zt/+jGV4BxbtD
c4fb2HobA7ATIEYPPkYzb9I12LEL1JL2LTu10j3HTNvj6Khc0Ge9lCwi9dciWKlDHGGltS+xjFzr
etkwNBLhiY7oTw7TFOq7TRDD9c79rQ0eSxggR7rgJ/d6r2XDDA4miKkFQ0x7xKKIAVPXJ2gC2yCe
EjImPjHRW0f0jZC+IiDo+in2jBiDCz6ewTCMa17/xDujmTfKIrnx5oftI2XzGPQCA1r5ACfMvqSi
uDCLXXAkyBKkagg8jxjTwZJ7CakJjGu50Mo+CmCUhg3m+aNy/qN6KU3GajdfbBKok6MzAFZrupAX
tlWuSlnHbe3ORsCtuKZlEetJkel8QLV4mEIU6+b4vYX/TgXkm0Wy9ihCJyg8HRqYR3TMHkp8gyeE
NOr6+rErhVhqq/aREDeiDOQ3iOwIzzUMSVSGxMYdmhELYHUEaymPjd5W5LPwivJaZPhdlcAL8KIW
5NApZ+ZCFwkoqcWnlWzb8rpFH5sIr7JEc8LJSJiMcxJI5/aFEcB7HplW9DpCgRrH8gx3j6KJyRLM
4548178xFz75ZbiuL5zmBXri4oq22NjGi/srXMthvrymkQBLHHNvujWcje1neKiewJ0blv932U/l
sCUlmfVzvYqjzX+BJNN/dqcvwlMscYuVgSpoFIdQ3aTOawVKhuAQCGqkLiidZPmI1ryyvEcd8aj2
UHGUWt3A9uORZdttnrhd4aMWiQHeBXdgV0Ehz66CmG2eSqeMN5AfC3kXqf3grVa88cIGc+jRnyUf
8CXJywYl4C7IVQj3IL8eCxpPDo1kUNTnWFl3Rm6iqAMFLdWB3ViGQhgcWCCPyGIo0NqpNevAU8FO
GUhN/PoS2Q8olKWfD6h2hZax8nEeCD0AzlhvI+AOo+UhxAFOXrxYa+SaP9fcbLZJf2Q+smqnO4fT
h6HiANBgWWM6Iwu4vRrfp4nLjYVl/S/K/mAidAzqeTMKJYhbaeK/bl4qjLdYJ25jr2QCjjtZXoF6
lcrDWuM4SppVXdJ10z1zwSCZF9qaQ5UWeIFVG5nbpYGA0Wcz0pgv9KHR8zXDeuE/pmpbZKCxVPcZ
vl/b0xbeN1ma+wJf3UZ5G3yeVzHf8e3nztZJtnpk030gmor1NA+Jgg9ok3uetbOy8O5/tzPXubko
fRcV3V3EnX+8IcmB07UpQu9j/Rrom+gjIjysUgJdjGTFJsJmU73/p7dMp2v1xHjiqqpm0VsUWy2p
xt8Mjr8SeJ+NdGh+Lk5dleIEMVQ3yX1oZ8i5ORBNmw0x9ZWxe5S5KJo8RhF1dLMfmGABr3LVfD5G
GNDFOGgv/MPq9oNiNLmUZLlLrSsRq1OfEZvws8BKWmcWbLtjCePSLkUXo0uX6217yC67FodkYsNM
i/c0HFkgIeA8WL7vRvDqsPp2RkVw5VmZmULrmwOGCgXIgn/5LJ6zUdUjyOh/sYYvmsvXeOcaQ2WO
5uxIrOuZTpdJAiDwA1xDhiitphjyXZrxd06Rk3dMxujO4dh5ZJr+bVTyQJ/rzaMQ+KvU/DOA+pHL
OYE9BOuYCmyQOPfC94RafBImTqiVbxe6Sul6vWVuXikNd1q0yq+YZhGRXUjQOW9CTQK+u6p/Qa81
gcjKAh3ZyV5N1AETsKuVf9HeU3YlIUFg5NVhVL1O5Rr/2roOOLG/La3A4geQEqcAVEK4AoG7TmPz
/nvTj4rQfz5ncftSi1Iy8ilkzUe8D4f7JkPiDQVW7qqkFMbsv5IsHa105lg2Y7YoBpEmE2rOlIjJ
wHcZqscN7ITAiBwvqQffbEr/uTpt43pxeReU0mmElwxzgOltmgiHIkz5w9HBUAkUKx0JMNa/URfs
2d9OAnGTocPmNnBiAUlLO8hmhrApwgYXXtF5q1hKwT7ZUyiP9wa+VTyscpt00AeZ+dvCuo8QIaeC
HUoD4yYzdcG9D3g5emer6+qLsX3PTNeZz/4l/u3V7cOaHRDDM/AVmR44Q7UiLRIqS4BdlDaaMnjc
6BWqny3PkGTNeN+fUuVVPe98hfHTSfnJyUcp2cKXOmqkl4b3UjH7KLJcUu3EIHg4Lsn9w1rRtQm2
N2EYdOQGCMdOsK2V7MwNbhC6KuXdnjj/XKAqZkG0rcsNS7czxrHXQfEqPAvSsOPP8zc5kYUuxYxf
+Iggp11OWybdn9w+VURgj0IXH6EQtQJpBAMnkEW6GHgtMn6LR8q5v6el5xsFCFWLUtUToSQxQGnm
rSaYzk+zwm0QwuoLM1k4DiVvGOPxshE/ROH/VpeiAKD/FLhRQKhTMo8HNRoO/G28P7sT8qGs2/Mf
Olhp8CcTNsSZPXrBJB47/Fy/6UezhMs1rQVriCY6uxAKKzws/95gWdJt93ijdKPqcd42IDaKTgGa
i2Dn2uJ/uZOYrWA61kFpCgfYes0OqiB9Ejr7x2+IPsem2R0tOoTqwH3JGEvIgyZRKaye0wWapRg5
krwOvPV/W3DbngYUUpQFlxt0foMYTYoSQa4ubjv1mPcPnDxr0AqELnGLN7ZapRLyvPjwiouXQ+ia
oIbAL360ThhO4+bjrTaRuiSFKYwI5y2APodYPDposL/XGOWV3A1EZnZ7uj/K7XFxaRv6yyHTcRw2
Y0Elh1w6iPhuLtHwwx/nZOfqpHzNrCkV47Yp7mgJMdgp4O4a2wkNTPFT7VymLFFy2lxrIxR4fZf+
dJ76upf1bgyO1x6X/3eo6DYHjRmH4OvJSv9KoEU8fMzZYOxLkF48RtyM3JzaTHlsyIPTSlp8d1m1
jKZme3GUikDxTlw2bUw7di2b1nUYRVw6SgjNfUcrv+6IYC3yCoFXDAPXwSafnMFRhdKle2hawvug
QKDnhHd6rpjHPzDXND1LbNggLGnpscnfTHgFUmmFPMSWRQuRW7gwAH55wBPr8yXzVTWTmxZGZxwd
fTYuBOJb9zIwSy5LfIy35NCATHSlJXEFm6VtMrGUXdAjaMpQJ8YGo0A1xtcVDnP8T8ybuvYPJnDE
kdNHKz7+iWm/V2NRU04oi40AbZV9+Aqve0aYHmZWXAOBPtUzwT84F2yhse+yrpf2FGEcHVKUxMqc
IlhSTVshB8gXq0PQrEfYD231V+WWl1+aP3x/chTrPTHFjO+LR0N8kVH9FVGAt8jYb4I7aSvuH0ZE
VutnxIhkx7KGzTpAUsPqWinZj5MYW0ildTILpoLSOxnH89+BoIh/Bk809LVK9+rEomWnJvUTL44D
lcOKVsqFb7TIxQNkJZ8tT2/Idu4PQiyMLSQO1HWH6X3P6sXnJoVli1G6CvLRBszms6HObwEpucmp
QzBH2fPGL5thWphaWXp3VZR05kVxIewpofnVc+at2tWxJFzKFb3lBzPjPUQGGc2by5w56dCL1QPR
kOR3NsZhRGNx9G7hHSMrKdNqlFs/qDKdAdWMC7x59Tj2j+PubqtECJQwJyi6UmxjLUfmvFATMPKN
GdjCbNpUdlomVvW23KCDa4YGMn+aDRMYkXZ51H3d8Vb7vKX/0n+5mLQ847R+J63IW6Eo1Ukg8maN
Q2OoWYK5lR7e8QjV23CaJo49yg+4ryFdr22cCm0/kWfkvjIB+Q+jzd7dmiotZTFwH2TRgZ/KD1Dd
3fRfPJUgy1JqfgVGrshhXtvM5EGsdnPCvi/2mulpf8O/YvWqZxCgh08RTsbZlAUZLPzM6ulwx5gH
v/MFZw7f1obQWXTcpbXTf6SctQ8Z1FTeKf2FQ9IjY9xN8THMBOI5Z98RIEReqAMuus2D0pGz550K
1Qc843kV7KclP4P7qdB6p3fKmvf7C0JKauhx2bhCe0lNhvMbdL77I20TQ09YRIGE8jBJ7CGcsFX9
YTAcmxSK2uNwuZxK2fQxDnHiVbj8/qRD+5LbWiMJPjEMX4UEbfjR2gB/Z/y68HzJjezI70A6EDQD
L4Cyvh7/44kSk2JE82uOeXvLjulHwzONnFrzDTT/jUeO3DrVTAScnGWGumeQV2is6mnLNV6BEr3R
9+oa2jYFY0TW89sb22nzx1IQLJXAXvoZBlNZuamwbBJf36Oiw/FUGzyVUeebouMQEuoS7sALE/ji
wQ9+1fC5QzOGE4VDkPn6vilkJthvppEhMgtR+3dDkD9qdiZhwKVNNUsSCEycQry5y+fKXiBxdj1T
q+d3e+SSdBpHmHUkbF/Ezttg8Po+w6dV3aMWsaIiMmr7OYdBUKcc+Q2Kn9rGQB/gBIYUAgmwJa3I
KtDgdZcSLLg7jcawMuTZPKHnXqlnuB3+r9rotK7DelNX9JaB/IxjC4Ov4yRk/dBOyYdulP/+5YEd
ld1n+KdQmmINSz1qbrzDxkEB9dqwyEHumbXqAW4Etu+wgJ0ZHZ5bA+//kjNk+W6ryJtlTFnnsjx+
1cRdATaEh75efEQwZqXxOmhuVPhkw4iZ4OW5ynt4UUg55UPXb0taw7dUxV5d+W9MF7gFCnnreaQ5
zWOY0HOvC5KU5d/UIHOqgA1XSEM31pB5OUFw4lcNtnnVks+33AI9SR+Sc8z8HitA/E/FFwmaJ7TN
0EA+4PNmKOzWT6VXuAkgbQ3tMXccUbAFN35Gw7bbTLvGq0oVP1QVTpr4dkBjl1YnDHrK9hN/RruS
mF6Sftei74a9LvKk5J/74+GioEGdB0UReGfnbj/2JvcFIuO5FXB7egmk+I9goN/9cUJ8QVcEA62D
GW4yPF4kuZtfmR2hgMit/k1uXowFQlM7T6qNMmsmy4wv/PG621g/hRLzKuXwh28ef6J+t+xxoq8Q
jwY/6gqh2AgTwb9Lq9v8R8tKHRKF40KTd5tHxct0yizPsgZFuUbLJjgPzaKjC8HGZENcSDW6ahVk
TQQgrrdeOYytElLeyXiSvxYRKuFeGFqwuBo6JVd7j53TKrB066cswk516D2JR119HrESEoUwfA4w
VRLP1Q+4ZpTvC+H0khSl/tkH44VavtO1VePrY1sHdP9HCUqxF1irqVR0MZWj4wk1bHvyIDt0IFNF
d8RfliuD9RPAzJdtgP59x3R8qox/t+auZTN3VFcHkMsTp4x/78370XS+fC1gtS+2OGgDRsera1y4
l0Qf7FMSXfgenCodaEDzyqLPFKOt+FZOQrj2K62ud9apqVhCy0pXCylNPlcETWgaFtrCXbK9Y+Ez
t1dBzWfIHN9poszVvM+RIjJACAAz54/zlnaE9THswcyGGG4DPySlnGjG2zxOlYbMZMt0SlJkSzF1
fFdBWXnDV1umOSFqJAwGJGrmr2rapbqMlmlKVVHSq8kWFx8q9eLxdV7t9x2uSDbf/+Oyj+4nfqY1
fvPh2o7iBXWOTL6i85UB59kEK9gINL0jAsVVps8ZJRbsiuF1gMKAtg/M/ueTGoYzEMttc2PxZpMM
iNv+bVnRqOzFp0eyDuXtj3nw1oc5rlU0PEK24iH3+AStI16WTv/OQ1XeEtCjVT2Fr9wTWTt/SWbU
chqZ7gNAqsVK1mlQMtrfwCKztdttym5bBKkvYRzrxbZOFl0z+ZRDSzeXGMFSmZGkkGZ6aOzf0q9z
0VjBovt2xWLJzUVksmykausx2uyLjRRbUtGvZ/OApVdGqWdfa6WlJZdtHW69/B8exbr3kXVqjwrq
44nVLaWey2tzrOKwMdZ18r7/flb84qt/0JANHQOxHtUFTXynGgZZJUoKEHJuu38rzuB6NkeAjDIT
3rhegQj8oFZ+2qFhY/jUvq+TMWf1HIapYeK8CzH+f7XguDwbeC+58/aWJ/hhIJjHsahnmndFF9h5
Iq04D/90W3k3nkju2k3PLYOZNKiBlCzXZ7ViRZYjI+fEDwRtJWYfJkzNwBt91vRsqW71Wgj6RuQQ
8OpRXtDmxXuDcWycUZTNFfjpmmbuv2OpC1Syu37qtFabIG/CJGIYQZz4cqMF2ydXcFltuC0GAJ/f
De6hhFHnWfdE2kTLCx7FoDFl6tb7WSIvkyTNYL6hncbDjpy8Kq9uJCl9jWCVrNlyFYW8yclB2IRd
gJUwvzqW6a7vDNHBETlpHnUdu50y98l9bHlvIc3M0CjlrCztNiGkKIJI9kf7xchRX1F6FxnZHOmi
dLfJTwB7f6dXMRqDkfk2D8I58UIW/mHiRoafJ7LYFrn/LrCMloRsAu5fJOWfnYWwo/WMM5DKAlI4
xKDM+cNzrq60q5PI0ddDTuVXQlGQdRUiT/sxTkYwBoNPkcEo2jYbYSiiApAvkd1f5QjY7P+eCyTF
0F/tUr4sLcTJVd9PSXNnI2rGpbtO8XHSPceFTXZ0OvUNwF89e829HLOVCXVb7qN40jm7v/z4/RNY
O6zGFmKvslDu8FMXFBtXNNWjxCmhBrFG8D3Ul7YrGOBtrBF789S4D7qZIGRUSrz4bBDrWa7JTdyu
UJfQiQmJP9Y9yBpgIBOe2jAxBnJIlvvcRheNbZkc/OFS7NBZCvXVvAE8I8+W9Qaf+iTMjgMUQtnJ
SWaJ9r7bAyAAsT3WsVcP49/GigJYWL4GY2b86CMgoYEFqmT5k636JpRQVfe1I3aJglUrSadg+30c
cDnmEC6IKiBf+RFH8ppRDNaZniVJH9jnOAafbBgd7df5vbVMJqwY1Q0V8sLvGtScLg++qi0lvCk7
0gLHLDbaDBPTGtLR7c9b4ks1EFpCDdqnzOTMM4Sxvb31Zm2tEmnvhB0qy/uElXfu/+PEI6iRI3R5
lJS9YDEXL1mkaHU92OQMG2/8ij4liEXDjENTz8mRIW0aG+WsfLht8428St0GdTyg7IqdAxF9ICBb
RS171nUnI3uFzdybYHCXMKVcyMohJWmT5c+Nlk11RtN7fdTj7nimx6DncIYMq1nGoXJ9CEKrKbeR
6IfiSReA7B0NIGfbJorUQWiA7q0lGnKPc8l3vWHxA5lxABWEaYPIEsAwa5q/KvP/p0X7y1icH//A
WayTy9o0H32+yWXWiTeHIzb7b/QjwQSqFpxhYbPiPyRZmD3DWdLYD7dPAso2ZP5oofuT26zeLQrC
LR5+GFSVwwDGmwml81jl3T/Rk81Oqpf5+UNFfjlTjytgBrfHPoy5xhI+WCfzQ/eHAcaMy/KeEEbB
rJsm6HVfwOkL3ZmLNvDQIWjbM3UPLwrfW6yE6h4nXXSclOxqfmRxSw/qSnAn4v9us92hCKPEzZqt
JyU2xcF6pnhpOrXYszO9ceHHqHEqSRS+M9SHDXOQClYBiiL3POSgmnmj2apyNGI6xfUwxQoiFo6J
wOAhQLi65CJltKv3cK8pPhNhHumX84hZMu88TuSupWaPunMjQKD3S5KA4KWvk/zt0ST6S9fQYtLw
aR5Sjl+KdfpF1SxleSVemdJKkMN/MfnBm5Sp34HLOBKqP1PfZvmOPqRyL9nauRZMaTxPaKWXMhLG
3I/hRZLJLaYgYgSmHluGVIxP78Yrp9zk0+tQmot9GUBq7tN6kLLDTb2sdwfBxfqJJMGnVSCQ6eh4
7vzCSK+g4AgP1XNh8lCLr3niS8enmN/RwEcGioPzHPsgroOjPio9+IEqBQOf3Fd/hSbIDpQvnZ23
tkysRGSStERdDtz+Y2t6Odz0UkomdKqNQBh6J9d8y5/Stcpoj6rtbwf2uyMOujhOzsiWQHCOujOh
IY1S79z2LDfkyGOGKWHZE0fwKRnUPhtI241zk4uL+ailX4F95Eq5XEdWU9qm8jLISYjEUtB2cizy
r4EQbAg7KuQYJYtJIou2wCffzIuCOzgTDqEGXnF4rhDO138H/uytsYzCNA8UUOVp0BGMofKchS/3
haAVGKqsd8UjDzQpyJjj5pFELjKPFbHUY5sFP/htDuHBEnUoqFJm80VALHh745e/xElLUe1HkjoU
vQ+z037W8YLwbbQgeE+j+QDPJPy16SblB6fmVJfccL85HCpcQQ8o1/M0NlTyzkjcYSZyu9N9pNqa
yzll4ORH4kb4WeIMUxLwv4dEzfqbYmGxtD+9UhoY2SdU3Sa+sxTdg4Ah48E4IdaEThXNViHAzSuE
CfUBCtMBHks7gk4Jp3SzXyElESTTt+mqdC8oVMMqBUGnOsiRedKr+rJJKKel5AU4ugmoopD3069w
PYBlD/Ro47KugJcuDkR6BuAxSNMxv7bQqTcGvXP75jEY9qBjlVFUqfR0EIZ/CjVztpd1DxGFiZ+y
HExKTsyaLkdq1Bd1cx94qj/2L9cykAuHSW2SikT67Huj6tX0lSSuz4FnuJIZ8e+tfM7zMWTKfkcj
YUngiMIQu/H3RhH0ryuI1c9mr9vXEQfw02eqbFXrPDo7tcIn7jWoEJaGFu8jqqCocsg/Va1NZ15z
jfH8RSnLLqr0Dkb0nc6/b/XvC/emabpXUpIxpymMA57ohHEV1lTSOXIaA/fKJoLzitIOx+BPzRK4
0EvZRKKtxWvlZzdp8o+NzjmzeMhnHcGfzZ5+Bi+mY5FXTdhnqkEZfRyXFCz1Kmi+YpHxVn7F6xWb
WLhIY5NVGUX668h2UsS93vrdwQmQDLzBvVx0I/CZfvB51Dw1XO0WppmO9USNyBSwcpLSV8rZgS0X
jrV3RPbotb9be2lWn3Ngvx00vJU1+axLc39TO0Nd9/VFWYOs9GfqLK4tMfqbsNQ/SMa0i12hQCrO
WS6RInh+zbXr+PnWhQQK1B+dH7pmg8dPh7eLDm2qsmiHMJm/F9fFQrpCQbIG/iQqokhjOF4F3d9h
yWjT9YpxgFTi9BWt4hNvvxNd9R27rjnaUsMb17x3bKCGuuEd7qLTfD2kDo748rJbldmNoNwcel+3
AXxYdUtkBHrvszq4MWMK0PvKyz6rgfigDxbrQ1/XRzloIhsUZafvgCX53smDVENhmCumzMomK8Ts
CwK2sK1QmPX0Uztc1+d0EKi/i6NT3RcOEw2klb2mYpGHtZdP+0bAxy2n2Yt1mlRJ6xyKB7ITEtGK
ZjAaSWK7XinCnVsvQIhnGN4OrjlmVK35gZzXTWRky0uSDWQW+bpDSXYEvRI2L/sgg6OigvMVQhXl
GkeKAgv2awMCIuQJa/4OXP5ysZnUW20QkIZojZs2lW8XX9uMoXSehjfpYJulQ9tR7Ghbr8tP8vH3
3mnlTXkcaGuN35IGyAchV1uNhCWpYUzK5/VFQtFdDNff1d7ORuVxnZIp+vq6cFy0GOLbo52xmHmf
b0rAqwLCFngB8ncXu4GYMV1hDzgIH5SI+M1DqRTL98Dedv2DGBWdTotdp/jaCrsVTx24a4tmXlnk
Z/UtfjxjIFFoXk5EYjEL9nB9DzssWUXk7WsUr98SX9azuUEMLaWgl982+xmsZTq+/bT0lC42tgVj
tp9DlYVtTo6EPH/eMQd7+b5Kd2bK37xPwEWW0nt/z0Vv5rOdBDIuk3dljTJyeLxmnhid5cHqKix2
mrpZDlju7EvXYdLtl6uai6yjmn16PdR4oARw/CZSpgQIRGSXUZ3SF2bJpD8lsKctvcDtaFKphPHK
YRhZT/E/g2dGax0hFBxO3bEfry/0gcQ7D9m7wH433qL5qf1zXeacKLXK3mJzXMPxbd/lEyyu6tcT
XJEKEUZjCVpyjmKtEeHzfwPXw2/xcXIY/PbI+jpfWrsa1D1c1UQeoJe1VTZXN7y9C/qcArrRmfzm
dQ+TKbzBjSCTL21vuNa6m/YNNc6aZh368SCrti1U0EVPvKyrYpg5xEM2Pu7JXwRG+zZyrHqwMlGV
lz1Dacxqbh6AKd+8dzo0L8Lc4wFyRyrsNP270tAARK5Mih5rSzbeTQB1yeCPu2bMBfDtI/34FEwz
9RixE9zp4l0R/W4meWdJORE5psV4Nv2n2rwVO5juDLFLhej7A//9dN0zY7Wu8dDTCTVHEN2ayMw3
k4d6zwB7kasR8O3qpXDmMgJ5H/xUe880C5swpmM1E4pobgb+7m/C8mcoROCNJgtFJMBf5jHx2Stg
hwcVMpZ6vEo4VAerpZijjbNkRfJ5YplQYRwM/m5/GBfXCuqqhc8j3udjTF0hGU0AKJivrAyEcefw
q3zYdrofb8xuJPiaztTgPUSyK8hXk5AsjCC1MwvsOWF/67jQ2UOwesy7Yii5jwOnh4dfpVTiqgKG
gXL0d5mvvDNlHw3XHXOza9NONMvth18mPqhfIPPsRRGOi1Ly6jRE9bYGo3ruykL4fEGyzNzzWB6K
ybySN+WGY93IC9bGhTrzDNsXK1Ev1kvuNtpw0UxCmkn+oQH5/hs8F0qtdyG90O05X6CBVH2t3gnK
xm3IL3AF8nUHMuFunHWU8aC26pSBqpk/O8Qe7d2Du9x/0RHRD33fWboo/dyuAsky0y6q5zd1o/fR
TAomlute/cM2Vp4AiYofFPjg+LI9bXEOIF1OfCtw9CSyEbabWasJpcLU1r87stSZsHwCUOV8gULo
1eYLEvSJwDPrUzGfkB3BtvxcU4Eg9wZWZ9FRiPkSYK02eWz9v8m8a+vXPWO53eIZBC6KXfRlZwZ0
JXqAWD+A8POR9I7vs3UqhObi21iTfib/MKJDfJzms5OXhPmdm8QCntMgdyFzqf+GVpSfBvIUTAYY
t0t7Bwk+4efKTEY3PS+q2JPdOW+ekrl4+7s2hL/e02P5LVDaXV5sMZBBQ+1BXiN4FmPsG7ogKbzs
IzDsR9ZrO7B31o29+RbOcHEjWJPL9RmSdzSc7dZnJu06lJyZ2IqLDGzDqFE7WpyRH/fiR1aCQRm/
AGPzljy7FKJXvfnlJBedAxe0nDwoWga062iKqYJBezuIoAtY7+h4g8sdJNS2Qu/KlZ0rM+3nYqXH
fzUOlsWj6RU1BoWH5q7AJ6NBNrvg1pyhCSpFhQ34S8k7CDgwTFYSG0phmtkbUKgLUtMSMigqn3Qu
z+5ZiGJZctrsNzWKD3vw1z3BdeT9CsSeziC/qQeA7ub5LmH2zvOGuoVLVAv9EDbHADswo2kIeNSX
NVIcBCp3/wgYsQP5h1EpxiRKiscUfFAOT3S+tnZjlS9hxiEqqNRmpXPVRj8GOqIozTwQG3ZKxSNU
PucwPhzvJNEID4WqYZyDum4RS7YSJR8TkKDkQ6a3kTomMwDNjBpDW0hSlRHhLd52Dns72/jAqALl
/jDwfeJwsGuAxic8OWXP0m+SN0InaFtrY/6DMvfV4Ov9wdbAJR38NCOJxmNumZ2B97XannH6KfU8
U8PGcKqNdQTdER+p13RJ0tDX76jUhfU/TZdllwkmRCKTBJ0Skn6mpy3OEHygVXVFHMRy1+IhSdCs
Rzdi3bF0mL2IHHt/N08LGRfbSSu6d3k18nE/5MeFsPL+ne45GRUCCEXVTRU3WU0yWuOgHUVTjnW/
OJujE8KQQ1OKXRO+cP+1KfvGXy+GVLOcr56a5J9UK0JWtRbehwfkktmtXKdpWRtkS9jTPsgbXfd/
LsoHG4dQqLC7HIGkoavSb8x5RehgCwNbuVCDfCwz/HUol7TEAdaSrtZhcq3r9ESJwYpp9odckePA
e+4HxzRf+QzKW0BwOwxCqbbql+DlO1VWJzSExREBR082MK7sJJO2mH9Fs1i21FNdgwWh3jKGLrIU
VHX22SvArkCdT2tLjJIb+xpXxl3rKpL9LjVMH2mcVWkPh9J+5MHE95Ep3pAMYgD+NX4wExU4M8u/
qYjdo493Lcix+lKENTszIH3r1HV4oEwi7ij834n3vlzssPlUm0/D7vUJqsD4+N8UP/eLRWhhguA1
IVby/1p1IuiOoeGp0J5lieuElrMqAFhNVaw4l4VjGEVwWhjuCDr1saj3O5pWgQ0EmiYN2SM78AHG
GvcqxqKX8HFK0tOQaXVVIBYtWCswuQIyqgU9pb7Tn6iJll/TUTe48la26hWWtMhD0K4uugb2eWYV
esZvrptj+lOiul/nhFDipPCLty0aaqQJZuuh3CSw7cn03CxIDu3b/0QZ8Dqe/6tjkUAES02gd9ew
UISbNERuaQOlv9DzNBXZMOEo/RbyvNE43YRudf1BhJUt4J8ft02rui9l/2l9303lffCwZEOS4NYk
tCQKYZrxKq7JZu90DA/mw4pI5eVrv4lbvup8VkFNWC8cFeAv98wW3THsBTkiiql+MC9DyTprOly/
ZgEBAfO1hUFQ7Mn0oW3CMupnI0KZ1WsDI7HlIAW5wqELNjHgc1rr+YrhyjtRVCk4zaQg4VguYZO3
KJAzcGGXOxn6Spp4W7+7OnJlovbHYTVPy1KRmIxZ47kcVO9I9hqv0iXuzsxx+dabjGSu3lrvRWls
Ajoafkx9n6U+NvGImfSdgFOlbIYqNERlRMIbAmykjLA9uvVVM7A84nil491J5JxgEQIAsk8WDUQV
ALlGakPx6IZUAUZHlzmiuDIxJx6RTvQ8mNMpO8TI92DtzQZAIHSZXt7yXeB79k90HNVZTHAGMDbt
cONY2HeUhOoqkxioTUZdFleZc5o3kUpzkAr1Y38KeV5ID/OZFtGXCxEgzdkCPHhxHLG+BNk3TEGj
yfwuqdsqpDca8XUNxRKralUm2y6BYqRbsOAUX585YPGvJ8rKr2KBrsB1FWHMxz0izgVEJDmDqw3d
01SPhPqzm7BnF2utNDbK5BZzzELg8zK9kJBVEq1oBX+er4nYs5stca5OrWfcr8lmY2fIEIJkRIji
8kPmlMtt3zkDP2dT8OcCGuglyErGwU4mgpuWuNGLq6+P1LvdIButTRPbgaXGAfDbdQzcyPiihf9b
QShabMOeHrmdSC/aXkGwmvdVXQSPx2gh5SI8LWNQl2fiiQETUdeHCZk+Zqb3IMPmgNHZXaPjjJJX
yaBoXNoncGqlTxBbpXgTACarYdY31r/n5cmldYkbFTwP9TLOeblmRVznmr2feJqLWwcVa+5nRlQs
H+tzwGswGVDgKpNHy0GGNS7HSEe9uioZ/1nBpC6ZItV4354tc0rShT1SborxoiKn4KliGwQ9+jvD
oq1UspIp4z4uhJtHgDJGoox5qT1jRwCIW23y+XJpgSeIhTnw0E7U47cxytWMR7ctxDhoCMXUsYIq
OpmErwJ33VF7JN0tA8HfrdrsKyFfCWEd/dCSJqIueDQVKadWkUjfR9QNpZvFy5x0kkjc+JO895lG
wWslqUXO7lT0F9hZ+baGIkF+cK0XU2ohYyt/cvktnGKijoxRcFQEV8eG1WCm5fNTQsyCJsw+0jW6
wt61AQVseO2CpuXi/oQhHHwmhJSSuapTmgrFzzdlmTveKbHVyvPzEr3QHThqptGK/QmaZikotkDj
9dhFjYnRa2xhdQuUeGGJg8flSMAye9a/x+S9BYCFOxT878o/nJmcRu7DMuh8ec2QCXu2/LwTmVuf
UB4onrCRuqwiUBKqy9po46S7sX+rOSyE96kivz4N+pBRAFEhZbMbvIZ2+fM2H6gntPtVX4VRwril
sjiwIrOVmovzSA6P1zGLuLHw6lgR4Wumbv08NaUq1UW8/kxfiCh138NqY5MOSVYpnVa9IstWU3vi
efz7iohqhWe/QmqscfIkheCSapvR7VPpe8NnPYhsQnMge0x+TLDp/lrNQnx8AJ615/3faqtrKuwz
G5NA6NAocj76mPVMPmkePlZmz3siTT4kQrwOthdFhoPSGVjCdfuwzpFNR/JiS+19gEQ4rb+PdMpY
WSiEJXY7UHnhOn/ZUYsEyXC8MxSsjz+c46/0SjzdVPQs1PCMpniwyW7OeV9MyqbUZ40N/HfWG+A8
aO4JFZqWGMkn+bY4rsh5HkeV9Bvk/RXmMIlJAV3O/cGHVtHgHcKTtBezioKCFvYjpwjsV36yXLsm
kaDNUQMwIJ74f+zko8OqWQfS+Nm0rzEHQffUF0DvT01u5w4/F4VlY+gToRIqYMy6wF6HXaUWy3By
/EN6qF95DulWvu2MSsBezVtUH/mIfg4MR48fUoHr4Bs1Gx1+Aqn42OvllNAhc/PZR1BGFuHn+vJa
cEZcJMs1/QNTeuugpPZPvBerIrK/obIqQpMn/NImEk0hRdOkH3NfUSleCGI0cPElVBGFi9ieQFEQ
iCURbCBbYl36jPn1dPvQDPyv8y2S5kGtQCUxyeIIQORx8jPUtmCQrgHyWrJvNq9Xa5mcTwgNYAf+
J4Jhb0tBRXMZ6WVZeqT7maezkGKUISUFkdZQviwej8Ue5n0fZ8uELospr/IgfX/hdy1uaFSiYoAY
1CYW054+HY/h0b6gM9h9juybwyDUzuOE6nRjyxznEJOQ3hXVBKx5T1QT3EJFiTYekNP0QeFydouP
oR/ozAqCNHBTnaiBUOZFtKKVAVycjF6/XbPY68AUC9s43hzCjyGekGEV0HH26iVSLhUuaBGZySR8
A3gLEbwynGolE5Cm0CcaqCYFy0OsCRV5zGPzZTk3HG8MLw/RE1y/TwmtC/QfimLW966QbluQYbrz
xBurMdvoZ+14Yk33JBDHjFHZ0nKQWY4+ET8QkqjwkuorhjzTA/MeUgBEY+vxNzl1fme9WRJEpIZq
HQcZSZk/J5KDGfOjyZTZA0eJ5JMtnwmaCw49tUlOx/OtiNgjNXjf8XuIPBqfl0IXXwBiVhXv6PRa
Bxc5O5XKrphKptLRPG9hC3omW57v6tzaCREZGENsomQ0RlFtqONf8nPeKXs3h6AtwLIui1fNyiD4
1sCMMUJLTPvi+73a5hAVYNEV5Ybitk6zyJbs0g7MNnESgvYKDpTIY0Wn/7bv0QaRrCgLzPNw/7Zl
ks+7znUEyBg4xDmeAn0xRgEY3sUdFXBPx4PKhQvyyAy1FgfaC+qFQmd6i3/tDlPf3+RBu/ZbA4Zu
IUq6R9klqu773Y/3sWl3pddJYP419NeAtC5aScCH/mfKTA7n6GVhdQVTvYV8LNA6Ymrnkq3/L0q/
xfHM7CbL8xXhCTILuVvMjcLgll9uJicZAcf6/RAJ9VxyS1eJicfXct7nJFRlSRveBEoPF6g93cNo
7ejfkB+gGDs3zt85mDTbO8uSekYp0UdUMJBAb+AKJkgRBKtOEcvB+Cozdh5PptlmQOqPZQcihyC5
JF65e6KqPfPbKLGuj1Jxc4a7Mob9JFm6K7GUbv2h6ZNHPS6sPEvg+FC8sGJoGoyBEY6R+LZLF5sF
+LqVkjXJc2cCYtOVQxRgIGFHsmtj5Fsi3o5zttUwuChzMpykMprhMgowkG/tx90by0aoZqExyk9o
k1g7L6wVAnz49Lnjg/oiaew1+pFijJvlv5dvU9tdPvKBeAopOUoRfeGN6zNhz4TXkGpOn/hI10jb
dG18Frv8S1y9SQK/oGJt/Qn2k/PKyGltuqqhPDQM6MqFN43bVXzb7jtmzMKRtc5oyOPSRZE8FsDP
zcp1YBrFZhkW9uacmhAu+A0NDW7zuc+Arnz9XFO+YZdPm4pgNQsPSVkWqlSN4yOPk9KNKfX6E7lQ
0uXPmkeYPX/jkICNB8OGbRvN+g7cJNUultyzOhbBDqCIMkyQsMOgguhkGNnQT8OVc7snm6mHA3nG
CdR85humWPjIl2/TOkkzZJqfPuhuW2sHAoUcnRsu6dfr51Jaz5PeKGs/WfeiZhJpCXUndJWG3XCg
5IDt1wtLFOsZZ8RroIbEo8egwm3tIiFDysI15WTfNjyAEVEkZ0S4544eV4ktY5m/YPgREW4CkfVb
ckW6u4iBY0CF5XMAp0kf1nFlLRH6SBbtshwsC/7FIk07spEy+FQCftUFGFPIfT+nzd0TIGsMB2zT
Uco77vtRt5nFIb7S4eU5spk2xBcBZmzHUsJWk61xAIGK96BxO2s28WCVa/2i2qYf20NYUiwRMBU+
riDf5mC/skUd227k5YCd+AdSIJGNJCTxNoZ61Fex3Zhks7snp1OfgiEa6oQLpk38IQpxgcDb01Ba
uxoFhqY92+0cGQ5xDZB8gS06xaFvu0clgnr0I4p9mXrPZC48ZloJD7asg7CwZzzVcvCrgZjv6ifq
nwYp6Myuri3UHAQUhUVtY0ugozuG+tvQObV129bVsJpIEf0J39RgC+QyB+gQWQ1t8+B6UDNqH19y
zMn3GmOgh7KF0RaYjQWfYSCPRidNW+hiHXdX42I/EgAhj6tZl0eXy0GA+KJrRuFeT3Uev5elOFoI
uvVeZ8hgT3hXcWTxIQ3APzzHfR5Q1F5m5fmoNvXy/DrmtJyf8Aa+rPA3AcQV5GcZdO8BkpNA8uXK
IX+Mb+W7PIHmyS3F5V0ZtRtm2ZqPHVUePavrRCs8jjwF+P4JUfqqxHhYbOnd0Ugi0dTQkGXxaUPB
dr+vVhTif53BL8tQkEhXzkTBfkt+Ro+IMt3i8ZsSlkXMpL0hy6TwAE9o4iEVWpbP1KXEMTsFv5l0
ep0cE0/2up3z3fJ69J6mYPPPJNsFawLWaO9FqguTHFSil5V0TVTnvSHKthQgbeJfTBPTVtqrPj/u
Dy/eSbyCPGRtpY7AIgI0druJLmwS+syxdcA4/99t6LbK7bISmFJKpac5UiAUKjz2KPnVoZZY2m+9
1JKzyO1mqsN3PvX7E2uwwtS2oAf0LYg4yGoszHyK68Mq5N7uC5DsRKD4UzHhneqDoEY+G+LJ3Ieu
eTELIUbhXSaVp3wWePS3TOe1UghzyC1Z32evZpbmXsBIu9fsn9XD8TA49yAajb+yYLbiqqUTb2XR
dO/eZAN6DVx19406GuqhLGOkZkxcoTlVtyPGOYjgaFfMYFbEHIdaqlZf3GMXGMheo5QzTABYaXf4
NhNUL272FEH0rtezyPM115HmrnegDdzSa2ZyNtfOMqVZQyGZrJcjzxPpcNqdaOo12tcdL89W/PAl
Eg3v+GTbtRL6CgFSK8ilRov4oze5A5w520bgPnI1TjkekA+YejpuEvlVS/LdxZbd7B2QE2kl4IWp
V1ihHb/RVkeeuMKNsbJw1VlWhGhLa/kuu7emrkbjmYwvZqYVp9HumgkaOsDtjhUBKhR7FfVIkzCe
8Ha/c5LQN+CILMhxM6JXXzucHHYoKODJ7ziyOUmUFGBofzzWiz8kI4tKxI/N22h5zU/0tK9S3pE3
BFioXql7FTz5PPQS3IgHpLocde2YPSpNXlCMXMxKEQu2YAUsUOHiNGknquGAr+IXeEJM1W8H92Ws
gA+8CujtHJx2EfbP9v5YfLJxXz6hSR2cio8KTkQhOZkyjQcsv4XygpBrOBQkIY1CW01JEP2Onrhx
hOGZIjn/BqaEy/BqcerwtwtESWdGLSd8wp5tQkwZNhSb88bGuv6URPJvmY/U/+kW83NSd8iWPQwt
4SIHHsWy71/GbNr4qqRXzoCi/Z+VxVKXMui8K06UMSXyoT5pD0Lqu7fPRY5AGNGdK0H428XeTqj+
TwivJ1zqfUcsyk9EEXF1W8K/WnQvMlfSJUudN3MMdRFKtY3iYWdxsuBJgoKjffmljQ4i4uUpTFLR
JoVe+UoGfW5hEortDC690SiYfSrZGldfAbjGh3HaWlcSMJBLdOz5S6Xs6Cr3IVou6J20oc2YWikt
oNGBOGFpJhAIRtkhicLFOmy2ZPeb72HvJ+RKBBA0IYjeYf64E1ARNJ6YAF0Jq85o6rxP/fjAQv8S
ityFRToLm30dYHLFE22baydEt8KY8RayRyUqHnw30/+eW1mYTgAnxewQ8fxF64qxe2ixti7L65+5
CdxfJzZkMHFF2JY530qsD2ZL/vAUXv+MkXklssyoiCYPXje9bAUkG8ngBoQ4/xcPY5Lu5JxAHogk
nGv8Vvhsxj5mIGsGDvHgLCx2gQEjS0siv6YPgxeaI4ZHG62Nmrg31Gxh02M4IOASBGI0xBJNDkuB
P4fQb13icvF5DzTapLHmkuEP39N1GPTTcxfGvcd/h/wvdUN59B1/pDE9apvOrxCi3eHVDH8706aH
beTwvjiUxdS/t7Tz2KxOxWyB5c16Z79SECyozQpQubdo8nZWlbCF0tPXRF3Nja6KGC4FcSbRUjJV
amFiqz1/QUD4yz26tBGsmjZB2RSxIygq5Ckt32wyeI7kq1TQgdPlPcAHih/8Wwu+iZc6mRFARkQG
CP02uX3PNcbKC6ncgIL6ZArXLe9Ar35ZsOmCOPrWeejfzymkuxSQR7znNHmiHJPKdQK/UU6+gW+o
VPzRqSqZn32yJCpm3emWwO8ZAT1x87uevUpkdtvGxjtyhFnCt64VpXtTSfYzk4t4ktOZ+YwVYJZ3
kGtQMjkBXY0wQBonAgI3LeexoXqztueBFY7sOW6ujEVFdCDvb2t94luduSfHCGDuFBo8xyMobNay
WloeZnrOtXDuTDdBwI4W/io0XIlBzLSMEaG+zDcCdskRqIN2oGzhKzB+708qf+qTsJzBOtWt8p9d
Wec0gadWoFiPAVPEIQcULLq3U/JoogjHg1+Ym9/T2rBNvLiEusL432b2iVbGQvGGljUYX0z7VU7G
rdYIXl1VxhHh01k0mMcZ+KzFVaVMFu01xrJjT/SX8b0ju6OaP151z0u/q+Uvtg9jtStcvr7RFE+e
ICsvGV53nIRTGlRUwCVv6zlu+K6zxrykSbAwtOCMnGcHczAb1XEEIS+PD2zxI7aFCsQnYJHML26E
DaEl+6r4u2AiBWyX36eo/v37ERcVZHgi1IxffzTUyVOpHF5Z++cte+TKmZo24+GI4aSOhN9gRivZ
eLyyt8n7o5IR6sGug0OgJWYdzw5WwhVpT3YvXGHlw6op5H2D7qB1v7Hdz+hCmpWQXTjE8oMtxnEr
BUaMLFM+euw5rH/SrN7XAOtmIRSdZghv6oMyzTJvjRcO5vjcZ4MaOt8OeGxY6MgUmXR5uD3YDIaz
gYNlQS3hd9+y5B/b+Ddmx5FPlvSA5VB7dNRjazRVbMu542NdAGo68yOB7Qh7irgUFk15HVqZBvSg
CLun3NFzYpvS+eTB1sX/a0ccvbiLJ7OZhu4QXim6QY1k8j/offZAAldtkxt53OdZYPnf+oOgI0qI
0OA0ChTOoITf3bwibMZwYWdS2josbi1jpawCxcklDB2TIs9nLGquzRaoP4HlkngeyuBNV5u71bLX
+ma/cbZq+ElagwCnyOULMS6SNakRPTtp1b+k5zQ5qgYTVVRvkMX5SiCVA0IuBNhHAGClzs/8DViT
MTNAgZe3vh7PQeCERUcSMkk+wW1D9pVstB4VQLMsXF3PcGxjvuCm+f/ge+0IyqukzW8NyzNI0G69
RDjASOF+yUX2uay1xfEo1LnO+78LxdHD+OAvKiemdJQInKrmxrzjxQ3skQA45jHjmlV7DhjQ7khD
UQN5YmD8f0i6YnmhufkMheFNup8gZ5P7WLL2hnIx59BvMN1cnMnjpf4S4RP5CDICCqyhSmfpgC2S
wQxejC2kdPGY9EGQiNCWqfEKR3D+KPAeIJ99hGnATtcehiA8YVDagi+zEysCP7S8+POVJXyIyetS
jWewYo4T6shjyE3vDcfjnFCxQsfQUu6S5Ba8qAK679pvquN+HIba07nQT4rLs0Ht5cJ5+eCCcRc/
j5xDFwKDGTkHuloKnbkQMKxSMtYGMSF17HJMlR5qbjUGbNKSA/U2zVfyAor5QbNw9oZ5OiCuCko2
S4lNv8+ZUME8+haKHyTtwjuKJJvIPV8Pv3o1tbnVijaeMyV6yEkoVSmXbc+kX/HFjj+YcqP8ABdH
Ye9OuuMn4o1lzXWMgvvRoXFNwiR6lDVgq4A5Fw24gUO/Rd3yleMzT91DYK7a+kxjsaMa6a17Qh6S
ypeqr9VT/PcAwk3Kg9lWK0ul6yz6nVPJdGZtxYpdHxAuWexubUMGvNRk/58YnWJrGd1D7FG5prLI
E8kluOOu2vJMKcd7a96N3t9C62AoWyjW46LfNiXk0IdtjJ+m1tgQqj6Lh7VzrqHVeCR0itX8gOvB
fCd+z4dijRtZySefwhtSgDmlibeV+VEnxTNsF0Imow+H16tEPhbQkIQlzKUINf7nKU6sxtUA5i3g
tR32g2kn0mUm2AQGv0ebf0N1fc+CkqngzQPw6oaer0B0VTgMWYUM3sORxL2IceyPwAfFVrKrfXhX
7+zwtukVN8yOL/Pm1SsKYr9+dmLkflDUzExp+tiifjeB4nBWaHCqrEyP54DFWSUsG8v9G1NUM/1v
rzvnUAeL7cBq9XapBMwXnqJZvNwpWet5tWCEJJqjEWrNX5CIABnCPcyGtexcvo+BOtVlFLddSNXS
WTOaImUzhKaE9iwvh395rPbyT2kWxzd4eGEO+Z5UxioVbOb2Cm6I9kRnu0gnZIvRScPlEFwrzfQy
9tL5aijqzs2XkKfGkPBFtMu+SsLP2lTe4ch/nup+/YJREpvChGK63M7ftS7cd1pFnsW6COXjXqLv
MQ0rhZqYIGlrlz6vedemkPdXOaK5TyM3X5bELvkJHpj/bBFsVfJJYp8Z+pK5bVg6jf9YgJWSmnnZ
HO2XGLrMCaEThyfzXaOymBC0RSw6HG7/HRvMA+6QbcFTFms9G6xtkERPA9Bprc8HP+AYTN3/VfeV
/hcjSVtvDgbuhE5AgOofn9efBsqFYi4fQol9aIvnoksmkHR/d3zlII96ytoFm+Etl+HaSoKLxF55
0GT+3TXeAoY4IYnc18ELLUty1BB1gO/H00qrlzEJfAvJmPPpZeHBLBMXX4p4Ws/4xmCT6PeOIWpf
SCaPfFifii0fa6x66I/fhceOZN1yWv6rmzfXD5YGFuVYijsKL2xfH4VjyCLejrkTHWsVgQGnVT7q
tEb+NDm7srq6BZ/+xrgDSmRGsH1WxYGeYMp+Scs47aoSvk1fMZ2l4uAO6lia8aCsHkGhSYuAMWDg
oaOBJXI0LuOOhXCmhrtszhThGkxR+WAVpz46TzmwE8uQYJW3ZcbkGd7TPKvEdiRC1468kxTB/MbE
Ri+6X+74i+5nMXGEf4hdBnAvla3sd0lH0KNR6TMs7BoTfRUUKoInU5W+OQa87catEtpKf/PmlwJt
TzJTCCeyN0nEIlSLRyP+1snmq9VL5/w7eoY25gd0yMybW7M6HFCecZyW/fa3/daDAGub+geE8J/r
p779JsV/cNUjHQ8BO9pARjZiahnapqgrXUJmXIjkVtutVQr5EhO9TDP23nf4DrgrBtYaz3T1l9eV
YniSxVpHSbkqZoBzrW2UGpB7XHLeii6Z+XhN6fHHAs4/PJpS7BE8Lx0mZiOWVdmr38IILPrjRpzY
ZbVxokRrSbrFwl3WD1UjZMhfLW5wGV2z6JBK0MHAntwTTuMhbdH047i5yYsDWV1vhcyPwQmBxV3U
lbBugFg5A1IHzQ2j7vIdKW7HK8g2ddz0hp0Z4UJWBc2JX1ca30kgMIYArCX4zWCqFNy1ASYfW/ai
C4b9V9fLFhEvr6PIn5nFR153quk156Fz9Jua1r+3+fpGaN38xxDs56O1sHx1gedEWQMz376Rjb6s
yKA8FadfxNeAnP/v9otssTYgyddtkJIhHxcv8s1etxze0lC4Leg9UFVU23tRMIo1io+9amc16NjJ
/9LnHN6ZnBLTpjF2z2fQh21nfWG0FZdusGHYCogSkkpbdPOqB4hmJDVBRqV2OFcYZlWhu44b9rKn
kPvZnwqQL4JJxyEcUmgKdaJw5FyON93SVMolIg1Q3uDojyLwB9qu/tmJzp1XO1miONJDeHiQxBhw
wK/IhiB5gA1oPyDtiDOS7pshKHTh2Ncg07eagAiN/mnXGuySxIt8hC8Z29zjsFZI36fVfaBn4Lw7
Wx0g2xc76n3U1nRt2f+gjlQsKd3lzi/0u/jZ9gfW5LkboH3a7Sn0GwBlb8twV8af+YYKASPMRo98
0J7V4Jy0dD80FHZdrmD3+/s2Nu+V0k2jV/T/Dv/3e2+ZNvUMQUX/8Ikv7pm5vFaB9FguRvyrl+06
mT68keixprYJKP8M4xdMLrv4VuLlnhsXGNcA6KPUn8iMlk15lbQZT02FEKWehzhxeOioywItGOuS
8iVtKoIH1InqC50UoqPkZzqEQmFxOJhSp/07PN5EhT/0QqCHGMVWYtmgJn28HwWaPjqnLSG7omXP
Kgj2EPk0k35ja7kSa/2+vWgNBdpuIxRLxvsvJgXs4OWTHZqxMjsKlsRRADCUsz3HdC93mjWeLi2u
dqgFkMjUyJOQFiTDfcrrSc4LdBl1pvNoV7vFvykepwuzRI1DNckOmlBBUVl4n72b1qwIf1o3vsdr
/qlIOP9FkHBZKMvtmlcJ02YWJ6LAy1dMmupEW1AP55l04PYoMIbSV7mKmZrv7xrr7Q/EYo/HKlEl
aJKjUUME4uZec7q3GxZV1Z1gER2mC1y65ncsuYazt7RbIcTwVc46pmm2/fbXvZqunXRq/++Xfs2P
O6S8jlf3XbZA0pKVx8cziaK1AqqR9LrSsmQCN9cfQpW+juEeZjvIUdlTA9E1/kq2cfsBzBZqmKQS
36ERNO1kBU1H+UtfetoeYzesh8hgbt2FsN73am7KmSCUHo2pgtIDC+bmbrWTkv/iT1KMw+gEDt7H
Lj7fMi3Q3TUR0HGvShBZrj4VJoxdIQF/791qkMcwtJc85fwJqcBcU+vVUAYdaFsnS57f9E3hx8Sm
QgEZh7EKMuaojF0hUwk4ZR9LG6O9yAVqkPk1VIcHSugNXB+s4R01u0T5QRtw1JJlLmxuBmUYK3my
WKrCRtX5GP90XjmwjTKXgzffaOLNu21zSYbATs7DoScHz6w7QjrX+RI1CZhB4ZzQLZyKnDhwrcpn
/9qhEWFXzJNm0q0eaVfZpasGoMrmjRF75aiciwEhOwrglNxybs8nwfv9wbfeuaKX+RhecwGnwene
Eg2uQYH/cD+d1pYlxUa3l6ZGhwvWJha8sdAuDC18i+yMUOazjfivNkaYjHcVeCT3HCw3T+PukgyC
IfHqPA21fxYqyA+0ly+XIZAkEn4D+EJqJTagFnmumDYGesNaynuWdyWLqPW/qVOcSQW6OSPZMt0G
BTP6BexgC4GJQWoxla8LkGA58lXAJ06lrxTIqgjwx7uH5+mGFkcN+CmdSQucqIGnuKyrd53D1g5+
eGBEzMaNars2LB4oZP3ga5RjlugzVPp83xhhKq2LUhzHduYOvW/nNPzWNPkbDlI55Uz1/DFNol0F
+PtpCD4A+4HaiRbyjhplH2Uke7Nu2+M/NUf5FG+HsscnRqDmUTdAOfM6iV9XboGoaTpRRI/nV0dQ
Er9MBRcCJHSL76wBTeyqWbnooRz2vLHfzEXkgKfDRYZNFexJbGUumaVMsMxdKtDqRecyvttcJNLu
s5yZyTzewsQp+o5Ry0eh8RX/l6GLrV92M9qap2UtBX++H+WYsDGh+XroqH5wwM+Z6lAh3G9rWtH+
HpYM+/Ceq894eN1lLJtbzsmULRRvp3OEcjSFeCZO4Rb0Y0fIWzDGafXeQrZML/w6JHqU2xMAIqvl
TUQY4iTkh0P902VvrVKn3onLNp2AgnRNL14HBVOYWkGucQunBVod9ruYI8ScSsldIhbQyEKgpm7O
XkSGMG/v3PS97sIbDPciluHceNYHuhvYodhLFhzZl0JHFcZTzNdEm7oV6SJYYo53yYDrcBdKWh6C
mzhEOtZ5jx4LgEzuwCGMerPYHgsriKnL/HMBRxudTbUZhGAAIxuWYwjUkcdy74WqfCFs6GQtp8Ap
ZKAv3n2LUscudBt3gb3k+bMN/v2bgBbzhToyD72w+whKNbZ1IY79ViYtYYungGWEA6J/iVzKbIdQ
lxSujMV+XrduisC7hk86bIiQprMMAHy4WeNoyUBM85kr0BlKMawTF/FLnkrDXINTEZsaK9JDbYBx
LzTjqSdLkeZQtHyDnJQ2It9OkLT2kPMFFob5KYhrhhHHanuXXkacN1HpfcaorrOSd2vGu5SBtd8h
m7c4x1EQfb1UFz316adGo8PQDcHynlAupDIecAQQCfZKy9cR+uIn+xzQO+/mM+/F39UV5hDiWEKB
4riX0kN+TBO0zIEpXp4rqkNGzvfVsCpCpKjxOTn5MpQImaZa1Oo4bE+gEIlq7Id9cgC8q80HX8gA
N9kTRJ61pANbm8DBG9s6C9VI2copfUhjTyCYGvITXx0A7wDmwBv+IkfNmmmLkTcJfEmYI5OPXVlw
0iirS5NL74f2PPYuVkVEwLim8F8SPqGf1qllKHirVvdQ3eOK8PUnur6NoYmIVU3ZOzQAc4ReSUXd
PokcgtS5hXQ8GFOalWJ3mT8QZcu39tvkIlR/q8zmdG0Ayc2R5lxFcb2kYIFNMPzFWBoAv/Tyn/0T
ai6uU8d9g0nnmpGeLix4X+qBe48MASQHG3nuc6ktPZ7P8+KyY/B8zAyKxjR3YlMPqR3fjW74dDl3
pKqECltTeoILONS05uLsPhsBJc99Arcp4GevAMDzE4ZrEsFK2Pc7kI8c2HQGS5S61vyd5U0aTXR4
NRyfJXqrRi6yOFMCMer+9Xu5R0hRK+No8KkFLWMOG+BxWYTNZDYKDqkhO8xPt4/IJIGET0+pHzLi
vl469no10534U1+6br1Lgpi9fmWTUvL9ViBQF2yceGAZeXTkUORnTSOaMmw63pGTCsfoYX4hxSTc
6Dhy8qMTvk7rUavR3qoLFZG3fGABCVE5DZPilzcZeUv05TzrkEsnft0hu4ABUKw8pQUftYTffXq3
vnLxJmBr2joCvkWV/tSVQKf3ehU6b9M9qKC4gwYr4GD6HIrXHoJbH95pMrGr9QSz+JpWrJ+XYMWC
/8bqpB09bCj0NHJyB8vRdyL+xgmxxeP5MbzkVg/OwOaBRLTubFiUuTwfyd6LjTedORnNILKJNaga
0qK3ekplGHTBqr4QB1BITDQseLw4i0unz186f8mFIdTr916ayxwYdaIFLAB2Fo2UIkYYevC1lOee
sECjPNzxYz+Sq+HLYvZSwQ3lvIErv7k345Jf8egWinuCixk3sXYJOVYkzU9vMtxN7HxYh2SVAeOv
V2cpukFunwS2p9GHfUNfsXjd1g5YyoBghhDjvCJ21Q0exNpIRqECDeNoVN6ExdtZNiviM59boHcS
la3VL4OLC9QIDEMyHS/eJeiHvIm6LqX04x0MkU8ZvqBiFLVvnsd5YjeLu++dStyQ/8G+5P+MSWwg
FkG1g3aXdZ/hqALdyN3fLcrQ3UvgU31SeSM0GYj8gzzYbExW3GZoBYd2yXvortc82ClmcTyJozLW
fBVh7/rf6Fl8+L5E+Qj4yZmeQHe1/vD+Nqeb2IErtK9ausLZ5+UPuqkRkS7VX6zgN1s1d3W96BW8
woPcGYwxKagnMQ7FlyZiRgOWRRD0q1yX9273XPuHl6ImoWykjPLqlKQmwZ8nPQ+mI+VGiQw0YQYe
U2K8I5p8uyw62PsYZUjQegA7ZEdDqth413/Xbtc8cEwwpN5yCyvN8I2bxYZB0cGoKgb4JIvZfDAt
pWgkoZLNe+d9kySmMvueRQdvHOLBwwujmQTbcx1565+6soHqsVfiRXP5OXwl2hfMfagstRmrdIii
nF48xHU3SYfM/bXbrEaycUZUCsuhkile1Zu9JUJFee/2zj/SFb/6VGE6xgvGep3mbmIeZid75o0M
KbWn/2tuT0LdNuqkZmXj4275KAEbSAlJ9ethA9lwERukWH0fuuiFCgz40YP6uFbWDaXxz5RPjCaV
K7KNIdReKWJW2EkFd3apW3Yqc9RFOzVvbx4RC3DHxOJ8TsehqSNJ9ky2fc0wYsQ4bo+1z0qEwJtb
uXGyZ9V1vMtWM1Mc4/6qRDtbsy27zstzNXAMrDxW5fbEhAndUJ28B1fVdVvQDhLjUVSoQfSRaIYp
fqqf/Cd9JvGAYHadyKGzoQt+LIGFHfQO6YZKsJYdf/vxrJX6Jr4wAjhrI+MZ5A5lJHi7gmnwCLJs
Q92Uqap4BIUPoRkxtTTwel2zEDUlBe+ONFe2CVo2H810ANo4ll3KLt1xP4rQi7hLVJXt8PhjxpsC
9cKHunlvKexnIn592pjWZU7IThlzbP5uIRs3+j5Pfa6Wwp/f7WztRcp1XPEf0smu9rc9r7Su6FMi
OcvSVLLqf9Iampw64tmkYClIsrjI1e61OK4i265gI9IYFtF00yjfPNtKY9LvFrJ6FDsfiVMWi+oo
jktQ+tHpMC62g7oJIrbqWvKXOwiLqQEvx0FE+krtH+sOHrK6b4zn+2Qpyw9CWSHtrh7zglJTq4Bj
yOEtXfdARdzj45GsUKH3LEPDX70S5LHGUXoXi8/OIm1Bd4N+R1UEfGLpp1B20pr+bn0w9ogHIPxf
WeNF/JFlmtzinVKPDExfyr6NZEDhaRy/u5b0JTRkDgRlqDHHqwFTa0+LRiqQiSOqTCUJzj1G/5U/
YIL0vfeRV8517B6R5PgBEkYzjV69K8qjs72OaQ25OYxcikfQ51fRoJ40XHrKHG2cLA+mDsAh5hqC
SBf5hYTmqEKZPgSqozC6VTmFaK0ZqezgJPG3WsNrwLtnUyVDT/aV0vbzMvM1uG4nvNRpH3/UomL0
OIij8WdI3h4C8VZAHc0rXkPVPDIk1wEfA45s/yO5O7o6FJvt/Kc3be05G/qtlJ8gz0cgMzdrQVpZ
cq7lo3qEdXxBrMkB3X8XpHO1R2povoS1NjbgfrY/sDHqSNVwf684646V9Mk6YFQXHMrXZCWp77xd
Ratpwnutd9TQAfDRvS6BpgfJc8YBVVuanSohynvHncI6E6j0SP2Eg6XjRA9RSaeMmkyNXwUhvExD
CjxD6JTXu+fp5dy9bxWy6ZdPpbbXD3OD9ENb7FklDlrF7u3Ih5q3E9jdaWsQ8P4KzrkZnka00lnN
GANFdAsmzFDmHlzPNXp0pywCX1+xlIql/g7YzZJsItLyJSr1l4k6aHYQbQQLQyJsFC5MOK1kTl42
QFtsQhjXK+468yFMOjIEV8VrOtdX73qne7rBSeDTU4FVGnfF7k6g09YlKb11r3EaBmJjMfpjVSwu
xrbWRJjGHqH9FP4K7Xvn15Vx6hvnE2xwLSExTLvyahk4oU7qplSthowBLswu0kbmRQz+IawPVFHo
5I8/gbNvB1QVayIEB+Lr84P3bfLzFjVtfrHCDWtkR6WpohW7ehtytqlXML2fKlX5w5ukUjCHINLb
3EA8ZIMLgFizXa17quPZr67IL7LrmjxI4B0dlWujyQCtYaFBr0Wfui/NMtvfrWn1D0cY5iDNgevO
oepsaHjiER702tAhEFLaCrPAsvck/Z4TfJb+R3DQCoHJxz3VNFP4dEV48AAM7hPbsKTv/DYLOxed
MIloaQAisUiNHTNWfmnMqEsPJxJvDIt5C9J5CtC0dGKELuco8jHzOHrulnD0C8uzbDUAmB26kExP
cqHXkVBIhD4tuJ3CiPu5zp1635v8pfKtmhe4ap8nfPA525kC2k3K1gGuaXSxupaTFHs4dv+Ij+DH
hS29ibA8k9MA84G24fj/O1fnrcM0eoygJmTnBqfY/WlrPAYr2kIweQtu0dTQzSJlF9VzFsbSQIST
TS8hB1BfbFBMqNhsavTebsjCK/uaVbpU6eu9YBH+4d7/mWzmk/neHXM7teladr17bOhCZWMbvbMh
sujGpNSKTtkLAV0FGybQtexZpuqAk8zxZ+cLhYA6LRcS6JTJ0hmL6WTO0pBN6u/Nvjwotdaf3/1Z
uryErVpEI2GQFlzqc+gQgEAE1+DJx3tWdcOCstTdqy5kTH50NO/C1JmQg0I5ugDUMP3WMZJnii0W
AUc2MOeEQAeqeRZaeDSYeVoVMJvEadrheA1KPPIlMzF8TBf4HB2suG5GW3XsS+LQgGozvNsm25Zt
CuaheNLlbMImZfhN1OWOqig1/KGpi5Evrhlm1PxcLBZ6VwfppSDUBRUE6Z7HEkXAH1zMOAWqfDVi
KcbJi2jGcYKT2EwS4Ayl3g70gzwuAuvU4ZMIbduE3nmfqsPXTuG4finZ2rBH7LrT3+rMQwp7TNTW
QNnaKO/67ZmZlahBz7fdiTYLIiOFpShAOXmNyCiXHrOV255Ppe2vfGKcS7C810O3si6ZqdrXx6FZ
x3WFBvy72hN0vvgDALlHtoCqUnOQ6WgSYVmX1iRnX4j6ZfTRHF3CAAIqN7CNw56q7UJJsXJvkp4W
M4JRQZQ7r67hP9l29rXCZ3EgDHgyhRgwJyczw1KiKT24c/zOMnB5gsAExzGVyktvfaFQEiw0x1vH
qBcrAKbm+893U91I0G+p1DYkU+coR21lUFByEzTcdzMEMbc5iofOGOcfKnmkqjvtfF7yCRuPNRPs
qzfsbXTccDakaz8+UpNJMIqCvrJTGmbhg/7rDiGX0aqUvg7JlyPLam5cULK9+Wq/PzdlHpBAoRjQ
KUOM9oFhwyQOJD0/5r38qOBrqB7XDV88Y/OCAJ8yU981gANQNEFGUUkKPlb/mEoTfJSz9mfdCLqQ
ThLNp/Z4R5AWvwWe3LIz494Ll0dgZ3iXXQg1epNCBGg+SmHZpHtdJXYiMc0ZqKN9wlJ75J+r52Z4
OrMAVgURd4rkLnpgjLSnRhjz5XkmQRgGAJscinZziGTGfyfz6uie3+XO9hbRz/WladehkTgwx3PZ
yezvUt82buLPU07vOH83AqrOXkWQpBw2ficktQXTMCljeaZhiEFgNFRhHjVZAuQ+ija/pC07HUFP
6tRCeXOnpH9jp4KB4J+vPeogPomlaRxn85ywr4//ejWafFxQPH6A0tH1OoyxHEAq9hBe6pt57Xbm
B9Otq4I79WaEkUNAhUhue5+4GPm3vs+tSPE4hiaOyjPJax5ZbPIT67vwKG9rGMLPEHcAst1VRIEC
5xbJK0gYiIRkf7vstN0WcseqT5vmBaGoqbriHm8sA49iY2Bz1hvXCMnsw1PfuzSWXrH0tdAS4axG
fDA/H5sGTUU/72HDA51S5IZLvqag9OK2mhPzErgQaINrtIFDuzAKEsxwThUq2F6IZWgSfYYLYVT+
FjZb+VAiEqlWrJjhkjDKz43yVsxdpt49DK0xmb3zF4f5ukmyzHtf7Cv8Mq2/35phV9dM0yZx910S
U+pUxuPCG3fwV97kCsMH5Qna86CqWDWstx8YdYLUjo1hwyrZSh5jx+F7irMNVyf77DWmijVLeMXy
engJeyqWuir63f+pqN31OMviWvFmZMJRs8vqJ9xBwoB8oEFrv6inULEi9BNKcVl7DcLq1lk1lVG9
SLxL3QNAwb3a/k3fnEDVdaVlp1TB8WdQirTXgUhN75Zk9yfZXRosITNYsvzQzAI3qJ10SuG2w4yr
bXxtb5cPm3Wf8Xnax7QLjZdGeXgAg1l8LB4w5ZNkZiynzC+yYUf4Z9byAtzobYz5rnSOPC5tB9lX
Gs/RHef2DzpKCh5O4jAwK6zFcFu5pRQLhoFiat1XqYB1fKnm2n/btGScNsrrDnia4nhoXiixiifh
qs4OASYRF0G1c7KlVKfyrmq2K0EagGTB+kAaRyciV2InAHk2cDXzAJ0iOT65As1s1GeEcnzqd3Vi
sf8qLAC12Y3ZtA7fluiU/AOxp/NxN6Gk+DwzTu0VecZWQEqk/GG3R+z2p8y8tjAvAWCNC30zH+Yi
kquGPDRFLoDJXta/WZjB5hjKPxsD6jXwVUpubSBJjnyRr/yagdGEMXm2Www2/Hqvc6rK2uTSDy7X
vVjOZbeYgqJLrXr6y1tbfCaF70Uki7n8HrRoMMSqHGsliG3sVBEhjHFuPb1eH4vzf6RJT6BxYp41
qSUAZd5cjxFva/o/4Mhm+dw/QuuJdE/zAJJ5QlnsTyGx8Y7UyzWBiCgh9MAN/mdGHeHL4/VXjNOF
DguXXGMhI0sz6Nb4sH7IW28FsWloK4Z1CdSGlT/yEFrlbf1ac4FjpNnZ6F8AyLG5Q8BHGAul4uos
XulAANQNGGMoappD9VZk0KXdQAHEvZg09QKYzo3Oj0PD8v7gFZ0s2YYLDDhcfncCsKdFxotSaDGt
3GdKu1CWBv8lmMZSonSGNVZvOAb7qGv1AwMtXI9ncHsY/4g3OBjvFuzxlCJEmoUX4kTj4W7Y96rk
Zqb+Qix1Gw0AxjrkbL5MwzkbvL0/FEv7RwS/XuLpUxHPqghzylryBMggpBOjqpxvU9EI/JzDaTA1
JfrBsG0J5jnoeEg333AaNQ8z1obwfkW5FYv0uDG1fSeBuPHPh7W3tQ3flKvDCIXmlNFfcjalBh0T
d2kMp3+dOH9lbaJLYEWlZdGyMTzR3LnO6M/XJRajaAX5CyMC/EWfI1QkFLQ8YEJMFhED+ualw7qV
Xu507HhUq5EchF94ud9Brvf79JHBRV4iXxtyrH8STobYnCbHhTWXLt5gItXWtIgZmKwvfWf0Snx8
K1r49C/miNzPjBs77Ek24PyCmy7OszSUn8DKnNNvbWSgTfHwzc9I7SC7/aNfDgc/i1Ct4XVUClHR
JbGieHRI5VEWMx7aFx3Rfes6WQbphlTnYHh7hvCDdBv4vW1oLDwt47YPVV9WaIEqJfNfq5mH8xmr
/4FmE3h1kRx2C0Y7OJ/WcRyrI0DSFYUqT4+kO6+kjtKK69CV0BlRcXhT6WXR9jDgMiiZXG/UIptD
K6d6+poitAYDEwDBJlI481NGtFQxEeqtgPXd4CnZGbapQiJ6C2egwbgOd675/QJY8oEukclx7Y8M
DmqOW2Z0+JdPtjamq9cjitR+VoteUuWvDDjhWdeYnd6s7gCn+L57Ukm27e8t5PUg614IXcsaSsxz
8MzbQn0amIpVEIR/pPssNQxEkcmOjrWkKZ9jo5M9yBH3NLfPcphbSBwCY88vfRo8SoR9oOHGKn9A
vp+V7MY6Rzpql1MVoZCmDNFjXXo33ADqoYZRVcZdVMGwA/y+pZ+MM7mEn3cV0rmu1+tMhfbRIqxO
M8uSfQ+OnZcnDKNCDypYmr6rLxS3D2bEhuyBQzBwhgqwRTFug5tobd28hFm4Zyre1jLNAoDhANwl
n4GxtmYHkmHUW0kx5YP5ahNEuAEN6G7SRJbzel2qROjb/HQygDnaQ30C32gbeOgwN1uR3FeU3BHz
sk9gRsSz1oDIgAvSUYuFnQPB8vcn0pWoaUorfDXAVLd4P+8SrQEiyoyfg7OTFGmc6axlN07F1TMb
dSjxqWpVumJfauE29wtkt4GZrr6gdLQnTSCPS9oNk7oH9B5rdIYQyZm8FQUIoC3XHdVWUmdKdiso
SngNe+qlasfwDIuBphuH5a1ralrQXPrk8PhKqjVZ/DTxuafX+470PUveXuEC265bsHWvURhtH+vO
6tfFAMuDDW2wGg+zaTakDySEz5he04dRRdLG5gzuBQ8gflRJULu44RtiABhZbYTHeF8FK1ACjJMU
LkBD/LzLBvjxnlluWHwPuA8e/OseNt+Lu29FiuSwEOuoKVlqiM1Wfh3FLqjsmYsCCRruii9X/soQ
r3L5P4u/GGSo8Z2CSUAw02q3wton9PoZ9AUM6RO5cCOVkT6XhvT5xSzffGvMEf9vyu/m7/dTkmNx
UKpo8LLrm2kF9VgvFo7m/s0ed6PRasHh/wHuN6HZB+5cfs/GveKaI17w47AGkcn6lcNF+kDOF2yt
v/0L8G08i+TcNEGaPl6FU7izzLSSVGPL6uW0BpwBFVtkqDu7ajGiDHWbLCXiuteRu2Yes74qg3Ar
JDwzOh0ADqG+RXr5LHHMnLevWeS2as/RLkMJIlMq3URy0N45dK6EGdFFjGECAaflaPn8nxtX5oLk
o/B613k07dMuJPAhT3f6UJqnzxzwHLeonIASWPmjoR2Ajt0MzHqa7w1doSogbkh406SaRYhmtgdv
IrGxnGZ/QWgnpYhisOkb/Zc9s4zdm9EuF/18yshqcSHG1zpIwD1cLvcz++aBJuKZgd9o1WwLQFiu
sxaQT1LQGHVhkWB8kTsgq2XAq0BdOcvEfnPM7nKp4xgRq7i5f8CVS3MpQ72xIoBfJ88KS3ByBa5Q
JK+5bB/r8GLAXVLc2uKcROFRsW7fmWeQkSMeeMV1+57zJcObMaEsEWV3oBMyg97pfRNFduGjfXBi
9jsINWoLUlYBay6R5U2d0N2KhHwtT8Uycmk7nPRshTFqbGPmhtfTFq7vH5thv5W7JL+2HDpfgCCq
oCntdoRBDUcKIxfYf4Ykf4sorzAkjKSqepLOLJO8bD4s3OXwnJzE5anDgJRHeAyNPNgemLdajY+2
D/MdJ6APiRBKv6kWCSkKpPD16Y0WnQF9d6ZPnocOfKzn3n1Vl8FBm04qSDXUIstQ0XjFw5g79nnv
KbSZA2bx6TFCU4Ag6EElEXYsNlzsK3FOhttfSehOzF0oIsrW9lg3d4g0w4m57uD4DrWWnOC4JD7I
a/z4WGJG3q10WwsA/uNnYiDzqmqyz3kXJ2SGtEnq/FnEsPNjsf3inxhXBkZanJcTbdazlZowF+Nq
YOpnjwug0iKfX/B0vSpQ4Yro+ExpOw/EA2A7G2wav4Q+w3q6Ck+gsiAkgLL/bsMNJZk883xxkq3Q
b6xtEJd6g/LmFnwM7pOPbTXrrcuRVTa3hDlzrDKFP+Yg1JBiDVgs5ZgKzX1cF9ICHTIjcyFV/WVN
DMYTeuRRHOZ4HhFePiqvFGR4fAUZgyE9CbClLRD+BpLZeTmcOM9pBj5whdbdWT81awN+H2TqzABx
exCOmxX3Mg6gMAEV0C2hRI+hPFe4vOXhztAfDp+aH8Aqrq807whlO8YrtPCU64vTOwu9GQzaL3jM
pV8xMoS2yiNiOUP7DIu9B4d82szuvpXVNTIc9qq/LsE86uI+VHu672lLmEvg4ARbOrrmBpU09p6g
jtsWruPmzxZDHdM4fXx27s8wkhuXgTCuOxZTsWcrd2VmKMoUaWng7H5FJwggTz9plczQdV2YCZYk
v7p5/ax0LsqMFDK8Hpp42jKU9fY2IYe7eWcKDFTdU6t7krNTwxglstpr/2sU6WA3JVmgbwLW/qcw
PVzp3iMY08wK/tzFrVvrfcveeT0oSxuYx/rCJd9LTsS0HhSVl4ATvywKzVo4QHULkILl0y3lij22
4MenoGi47PdXxoDyVX3fWIA/Bj+7GFd0b/qLkjQbRDaUVZOLfb7/N8Fh5gbaHRu50OGXFJQOYoQl
0jg9ejI8c8F5/TV+2HI60jAdgETA2wHO4qkkXzLt+o0sxh7lYNKL7klAacJd4H55WpHesFzucm4l
Ovl4RfSWLVIfTSxqOArEbI5kj6XfRmhfdTD4csESQtc0AvNWa8a9NQD/ep/K13yacfCnMnl4Moi4
I08dQiJqWirQbYl7TSAYo4yWtK9wcMM3UgDC8jAYcopNherlfLpDMlMXPc/aXBzLwZ8XvYOXdBug
eUGAtfDMXsXaSzRoCq6Nx7x7C8oL+vVHRBJctD1bQwkH0NNVvUyk0ZXa0J8kuiC9pYlxRtouR8tw
rOWjm0KykwD9cT9r+97C59kAoOMexyejz5WEtp0ov9Ij90hB5ba3rS39eBfKlK29kg6JGKKlqFw0
aVx39pOn72SYRBRXYX0Fs8c60OEmXe0GYLBDsCNGgt9iFBvZeeEFuXhdLtDR/wvveSWiRYs+Y0lW
BOl0AbuUhDeHwDKyxyNLhqOtiGXsMlpD7DUGUYtutEaZlIh9pXekpEslQp05bDzppdovKePIwN9f
17/dt0Cs0/RW6W2zkgB2LjfWD1JgE3B3/yNFoUWfxT604DA9S1WqdMWa3XbcOQzGWpA36jl3o5xF
9ZumWOh+ETOic+ZkXuijZmpfLrdSbz/KvDLGXW9xRvCj9hrmSwc6bRbKXj/Ndt01EFmf1Jn1iUdE
AF/zGH+hF1Q09K0MY9XQSdlY8fO0wuIcNLw4lG0PWkr3bCq26qX0AYwQrvwJLaHFEOEQUnTkBQ8q
HaKG5u+g78/1Vd0kpo/sjNRzeqHPcI38fL3TaYOLoqrY6XHvv00x3LJOHpceGcs+/f4VlRlVRDbc
bra8/OCFXEj4WX0Y40n4/b9E7/FTWzyUL1g9ZRkzmWAUglih+KEc9u2qz+Ho16tJK62t+hp4EQuv
wqRG/4/xrf+vSRLRjcC79Vm3syFIh7v8TFM9bIkXgyS1UarQ9UNXgGoJfmJ3mGjlajyEbqr/WMyz
MCd9DoZvLqvNZjwpWIBkAQKet09HLZNFlQGYnYP3VFslLDaz+63/C43kFmMrDPETdGEX9nppQ9Fm
m8w5mvseL+R6m1oEV9uWvARbA+RxjlpxRkODu79jZxKF1jP2M/3eNod2c+qUujknqm5Y+OKiQ25I
EUoutOFSWQgNNLjLabhikMuxPmvIhZPPOTUnlTTDlEBKXkq1pcmKo3VWvvFoROMCtWXUV9tXaLdP
5k0FK1RP7nTamDvR9ubLRZTcuQfsWfb7BjKk4xncrxzl01DUaARZ8LvViX+LXAorF1GXmqDKsLWj
Gs3mE3y91NjKS6A6Lktj514Mq+XjetbRhOMbx/13sXwVcpHdpdHXroeEVpF6XrLzgmKufFfnuJ/H
WsHdxsLlQwesQDtl063j1/icWQn+yvJ+UAk+b6I7vv+iIGBlxypiIm1sDdWqL/oKNlpKddEqV6yE
DTdXiyDs9SV0VYKA7Bx7L6E+jvWJbNKX62cSFpI4l2cHkiMdlJ8K3NRanJ0BB8bOMZEoLvoC7Dwi
KiB+XLJALVnDB6IF7MhJRQKc6hqGOxFdcx/t5aedkpNgawLogty31j4cRC/vMJvOUAq+pKPk9Wtq
A1dys8y63EjE6UsCnDK+17LYvlzBOxZGCPv+94pmUCzOW+8wS6HDnwyMHlowWyBBzaT6CxijdpgV
UN1Fy5sRDeKHnsbmbwh6D4O/sc3AoB8mgbJKmCK5UWzPhQV6yzGpvwWQP3aBeH8qwEz5uWbDeSlS
Tfx454Mn99D6gkvGwM7WUGBNIztNBDqPOAsSYl76tYjtrZ1xjhIyb+SvK6aDBYGTN/+P6ylfNsOb
+zqUlFd+D53QfrTazhQh7VCV7Ydn1qctxrM4DGEc2t/utk2nPzon+DsPzCiu4KVogFtQx7z6xPlF
rLEzipLtfCSjJfD7lYEDoy4CYWYyBn3EKYGI7S0QlZSRNCvtf09v15OmZIUbTeTj0kM9S1JisspF
szzIgC9wXWDFSuAP80W8NGoP7HOtriP00SaebI6F1wUhnV5K5erWVXnEp4MGsU1QgE68a9/z30Ab
jiCefQDpkLcb+Z4c7L1X5GMMsXGTWHs9w/tuBxh3pGxpecnHxbU0gMgjh62WpnwmBSyJocsnRUqz
8BX6X1ILGSIC2sQoI/+SPvwOrfadBYwqe4Y3KEvCtQ/BDHjOA0X8doEMj8IGOeWB7jij/DacGp8i
Yt75WxckQ/oEBFQnVxoTZuZew6aY8//8A8dqtLzB2yBAOopPICJQ55L/3iuCgavwY7J8L1WZqEv7
fktR2hrRjePc7W07MhlMIJ1lY0CmMLa8P5KK9SHvUn+s/+8c4BaXOWxGLPMH4SX0mYc0yCCtSu78
MPqOo/1lbnFWgC6Pr/IgtkdZVZsWk6yAyJdbOXeBoOZMO6QwxAIRKIIKvvMIBmv2aSUNN48KUfut
He2RHbl11C7Wyx1e26EooHlez9EuXW9lSQCSyjzkzsSfzAgdF0c9/pHiyOE9RnOBibOgU2qkcjql
xBO/SBQCK1mWnRVA/VIe7bqOy2UpkyRKpcvYBcUj7XOAZgJ0N20clXr5qCIFb6f7FhldGFO8CMt5
HzFLHqe58h1N658ZFThVXZfat6RSPtXVJ04mT2JzdR5jDlS+4Hj2l3kfW/NJ8GkRdRBxndcJescU
AW5cRpdHQHTPZJUO+xFBxBPXPvVYOMrKf93Eto0wWMKBieevADIp3W64qQ0N4OjkfMzzRr6Y7P99
lm8H11Rnav5zoC9ziB8f5KtkfNcoY9yHjZrVlB/28eEyjdgFxtyNhvBHykBMW+urNkF490hJ1wO7
Lqnk3MXDTvjX1xKkYWgKJscURYWryoGjFJiydLoUeaPD2vKCSHtGhklbsqAQPNefbITesD5GCZly
p/kmBlRvdyROf/IMqdP93kFt5Iiqb5xzxAp1Mm+ZyP+ykQKCTqdD9FvJ0i2V+AVnHAsHhNuyBgtV
kDp6XaHrxUupQasBkoZgbNcy1JGGN6LySK6jkDGRRWZBUaW2oPhDRCwlJjNA1qqH3HCtURv1L3g2
rGwgvg6h8MsYWJAJFCx2tnyv5bNm6fQHHepGKy3BT70V1tnKhi9nId0ssXeq9ALD+eez8U4E7Ifh
+7H+s1+zhG2ggGZb0+PTCppSzQHnpOSHb7tpv97vXH0esGy3gDBFBTdqzcfYvh12EfTo/qMb47AB
7Gul9xd96yBTuBJpL6LkspbYfLP8j9MLNiDSJ3kP49uHq5PODXMlqn6f4OafVAbaOIvAatD6f0yx
5WGKbvZtsX0RbXQTXDmRjsiVXBu8hZ09DV5uoPFA+lmApOlngsvyDkEXvg28ZL3kU7L89fjffIsN
sV3U/fA0iJkutTlVvcGsI/sOWNRjL3BwpkrXJZ5AHY0Lb4BZpyObprWZuwYWJ4FP/M6eiEewJWUN
ogtdOH9mN2QhwUA2nt/SPcjkP3rJO/v3ICHIQfvxawhllMOxlItFbSvbPblojGIsVNvYt+Tk2bi+
GMY//nf+lmdr1ft72iu/RptMUluv/IzL2ynQcoLPxH2r8efEfH+Ly3DyOBofdXXFNOrE7pLeVG2N
x2ZXWyCW4fjctheyBSFSGtCpFOFKc8Wt8h2bgxE4/NlT+5QvGvQW7W+zxyE5yJoghSEQ6k1tHcc6
uXCDUG/V93YcxgZx1T8fXq9WFkypnU+RClcEd77gwrt3dzqbFUFlo5ntWF3XYAhujoXciJfgy5gp
LIes9cNd7OdChQYiN4WVZdhtjVg1hgDQeC0g46laRDqrvY5Ymd3m7HFqWFg0W6q56IH4XY+HKYGH
2xaBJiYHBr61S53pdcCAozPiHyqsvLXHQ5qBbMsPGBHxR68jY8cdT0Px7Xa7PY3yfUWkAqdaRyzJ
FB33NpxaMUN3xdQNt4B4D0mdJAq3TSHecld26k4J6c/W4SeUP7bEJIeXTHF5oF3Ca9AI354+SUpt
nBt2JnZJJpNuaz3BtBjLJU+0k0xzIsZ03DRcojrOlLhBepb8rM6GLBKQrhuYBMGNhpV8Ybgqn+4n
axyO1CBLcC+3jI2T+n9PI1zS6ySZrJMD7uyh04Tmh8CJcS40LvN59bIhQOr17xbsEUG8Yv5E4Jmv
LAGbjNDwFy8tmvHpOBRf+AQBWX7jdj4o0sJbrf23fTv17O+bt5I977d+1kcLHfxNx70ob0MtVi1s
zEO4I0nBtuJs5lWvksu2kD7Ewao/D0HKHI6JbwGics8tc8FRJ0lK+npwFqjVO2BwGubJzGhmXnG/
0JRJSWbfPDGc4ZateAzPNxoTULg3Xvx/cvXxFyo19aAED5s2qYisOc/NPayyosyelSKn8p6qRPkJ
5mzEOEb0yzCchEaEwiOiwwgzzDFTLMqmzty7jwKgEqyP09+cYU98LKxU7jEpY5CLVpbjnUPwVE7b
Git6uEQkCJ2eMPAxmtYplXGEd7LMyoXVxRo2DZP8ggmE+ncpQ8e4CglAFOrA/0hIm72OD9bcM0vS
HibRUfOlGilf8MZ+FuYrwYq/yKhTX1iMn+DD6wEpkSGxeuJuYawi0O+gBHxBxOnP3PYooqpo81+f
j1EXSp9r2iEF3yUwWXpQKtA21XbP9zduZGQGb22kytZRRL4K4GXbjAYOz/PCJiPFKjgGEifew2IV
5kQZIq9ilpV9VkeWICPiNCjdKCl4ChT858KCO7H8RU1qwJ4r85scbwtnQcEjwcHEgTXVdggS/aFg
FTuKAW1eRlBld8h4zwmWux7IUFZHUP7PrKIpqZg5o15sp1b8IE40jcxdpbWr44ZXHrhTUfSobms5
+dMLHFpJTIDLkyK8TnJpK6n2QhGEyiTKJYf0r5ghHZtOT4d+xu6zxotycpN2t0X1K0cPnEpsjmvb
uublj56TwEG0ylkwcEZTf0+7SCsHqzsp+Zoa7xTo+5gyYOBxsY3i0fy2ryTQQhocop0m7HllGoBC
q/4qKB3VRgMqT1SDCVoQkzA+p+a7F9VWP0lI0NDu1EKX69OuF5Msh01hwK4mABYkaPEd8EI0UlR/
mpZpvA7a7yMHaXjmK7Zx6rZqg5s+3qR9RzaSiQQp4db9Y20wbPLKUHmBXAFAl1oS/53Gz5oToZ9d
boh9BsAcDtuV/3k1BCbmkmLmmzU9YzAL38NleZaoRgW5vosoHxWYKJRzXArZwPWL1igdrMIqo3rC
rTmYsOkmnhWqsLGPVPEFWEX1EjPmUR3PsjTxixP+bIOQ+U/W7lklMq02tkg4FcTz0grOM47udSCq
Jevdh5ZBnpS/ZvRIc4P4gJjcPRujWPAV9V8ouPGwvm4TlI++fl187tQ+dyxz+GZiGLlj/yh5ny5P
cv6YGaeJBAve+q/7wJUtNuoouOflUpJgdxafXNWViCbCe9QVwx7FxXrgZr4q8qhtF8PYho3MDkqh
GoFnbHQMtSFWuZuj1RJ32ex+lh0JleaBRlKGe8/fZyUioBfc81jYomwUaa0GlIMNd70tzQibpxSl
p+eYcHUmMuSxwmf2stL18K6WuUkT1KW75TFiWsS1e2qHIF3x3yPepRRquNIBkN/ysInJLbjDsur7
cyPhd2hVOvh9pzLMQVPVUqqP0s9rzbJUTP5Vp1dma1Z5sUvt6MwH6elGW2HHM1kEB6BwtRY9NztX
WJsDQIk1Xc6tMOjF6T9bFraU0LR4EjY60Gw9B004IB6aHyInhVq8a7Fj4M3S27j3oZV48UJ8dkhO
iRIWffBpUEHKkUHnQ7XAl5nYmvPzXGVRO5dRA6UYVtCkugjVr9WA2WtHFqx/rB14LhBiQPbIfq3r
1n/UcQs0v+mnYte4SDf2ic5ybQOeVtvt43dz4EydcDmfMr7dgzD/VI0oyne6Dn9w25+be4+by+0S
uqwhQ3LRrZKloKKGVFEQ7XHjMryReTwfZ4t8Mf82p0IcdlOC0q2O9BX42pMGdBFBR1szggmvmuZJ
MS3+QLvjbJ+LAID/A5tjiIK8FAFLOdZS/mwIJjEQJ0wl1/d19biSLxncixglK5WE25yGZwvEFSH0
noOafKgTW4hC47t1G31ngvzaGWgD3Fu6SDmuhdz+lVvZQYUd4DYoG1t9CWzogn6yb4Zrkj6nmjxk
mcEXfel/7aRCA/QeV6FUaFGKs5n+oqzelaD+TNwIbUClUPEFMlDuTTQiLGp6IodHPmHRMlQ9p8eU
hIrViAwKNh9qHw1EDmBfe/PSdq1yU8SRtoP/q9CR9yumQqgxK8IwRGL7GAAg9GIUenv/3aZ6Ya+r
+YOygMiMEGOUczfjpf/z7uhBcvHeBUxKCYOVK3ytiDQ7gw1JxNN2iEtjWE4ZikQTHAlycF2Hve8n
zYho13v0TL8zi+k1XJmSg/luqfs64eF3znQqymQUgsL+kmPYmQE51br8FZIuJ9B1DhJgn1g2UPf6
YAKj+6rD4dxv4aKovLm6wk2FyFgVJmVtRsOSpuSP915+GGOtPii0wO2pKa8Nwxs6Wud8av/meNOq
I8WMFFONVSrcpEAPtGEuopQh5YNMWI7536S58efzQzBAro25/wHggFD89u4poZjjtOtV5iDoTGdN
34efyLXs+R2M5U2Y9BF4v3Rfg2nrQnJh7Fk/+7yaFEwOk4bU1tq41GTmN8beJQgy4UJ/nqb/H8kF
Tk+rTUVbx7waYXMRWGPlSmzeKw4/GmyfOgI30BQv667l7WcAFwh6wCUBBLSfr3gG8fgV2WQqmLR8
ooGIfl4AWyvb+lmWpjoglDBNip07gw9+VZby4MtsabLvQptqP6ykC1EQ8bcxh/SuBgtSMbW22u7H
CMS6upCccP0PeJbrutoLYQbMaRsEClUNDfd/Po419/WK4zSUjkWCOGbVFmpWntIAedOcNek8mo/N
Yyn6BAjWuqmCTl+pa0xTC6qsjmmt0FCKYdEY2CmHgQYHVUEv81JFaOzlHSl0F+0LLsRVyP10FEkD
ngb5GhDDJVh0ur1XE/0JrD6jBuwl7wO5n1CMdbKIk9anMI/Mj6ZfsMs2YY1gKu3iosAXJNelmAk8
QbLdBZj8qjD9fbNccA1i48qHNh8KqOIJGjVKYi0Vi801LkVz/+Ho25MdC7A44eK1pWc4DAerz42q
lmExxf9q47ahFAg9d2CoDRPcuuMCu6xnEnqisPaqYK/JzVGt8XpK93oihcv62gNeIVYpQON5ILIS
n4sIo4z3/O3U34O0H3+F7UjYULAG1w04/2BDujhJbBVcJrA6vbTk1zSVQPo6mZSXb3QlUYLc7w1/
ibd58sNbTmSpZNPaAVEPW7YXWDNmgukomgZup2O5Y90nqBAPVPzTx1bd7pw9zzHQnJ0/1JN30gU8
4J8Rbm/qmG0rD2ff7aem6x9alJjPK2tELruNefVYHWbJucNBg/x2miyqvGVOcT4onn5lwrux/aHM
J5Z/WsK0gdoPFUMm2Q0Kb0gCvnq4aeo0tkwZL0gvYMqfpFNmriJP2a5slvLdrWtCKt7LIWAet3V6
XYE46HLIJk4TVxvzjesW6PvJd5ZSbaNu21AFb/VPOp+9YjqtcgK1Jv+eBUTdLkFaobrBfnb862gC
rhcEU443P8EPpdJ9UZn3YI235qY9A7QuJMy4Xd07Q4lB7y33aAQ8ect5QyXSVMdU3H6Bf+ovx6i8
moFw2Ax8ht/N/s/+U0aQ0DoEDssloYXjsVOYHQeETjvZcfy2w7gMBKu3BxtCn+bl6DYhsH7BHfGr
uG8RIvPRVW0utmbBH2u223IZPf68Hogu+Dox8fD+d4rX0e/Ew21UG0VO9FRk4pPhweLRzZU9yUQ+
dJzlJ2qurZ1FDcktWVnZ4g3HlWsDcPHMxEoBsbJJqYmE3IQNCXAz696ElBZK7Zk9vC7qbye3Bf2C
hgTTItWFcnab4IjVeGwHlI7Wsk4GsSbWeciCo9/GHiX901z27aXKuP3R4ELAyu7v0Umqfq4LYNZM
M3QMkRecfdOtBtKGg4bHAdi3gjgZ+N/6VryvsNaSPXIxIRPRrjJpuo/qcKqYIrCJ+i2OFEN9kgOG
wOAli0m9ZifIAPhTtBFahCxD4iD2lpSonMMyHhIM6vBFzB9bvOYGkSpUxyR2ESXxZftd5kzHWnnF
iA86j0ksBfNvW8X0VibmzyzEPe16etp1g343rYfnGrOIJzxsP7nFn9EHR4vRGnhYt9o9pwoWNUHD
SlTfGHXkjFAqwFPDylszYZvga9V179Q6alHR4gxwQ9SvezrWewTjm/Pu9SvPdl/KBRelu9+h8AIc
0Wm9JiSyr5DHTghnOB/JIV3ax80fyblOhSAzRvNJ4ZrbXsi23Yy7moZRu+/kug+JIXv6DxVybcBc
PDP4/2aoMt7n1TTu4digPrJgAcepqp9cyMIW0NBph0MD3zuDSkgyk+ROUEMUuPSDPh0e0EtK3k0O
c5cvHBCrqxrHg74z1YtGLVrmcrULV8v5YCnU99zMbqXX/iqzNW7t3DZjXsn10gshg+jHQRXJLNky
YAmjCqJ3JJDDQ9e2D/wxTJs6CfQesG1+bf5bCos38paXN/kjvoZo/MqFmNY4ITUu84Zc1J/ehNMk
ooZXfilZ2yJYDaMKIA5gLiF0sdiQdQG0XjCF/KOOW/9wX+9e9Tc6t8itx/42letb42rGRcotIxSp
q+7EuObB1pXlEpputFWkDNbmNY9VQXEeDzk4kEDQiKpgH/H5MZc3fApZlDk3mQI6uHo0CpiHxc8a
TuSPDFQtcpMot7Nze4BzlX3gFzk35c7hN/YCN46L9nkRitpA0AD4ZGAG6DK5xEcaU4sai3bPhf1y
1ZVAcxWqKQcGGMoTcKsxenAwTtfAxb8T8Tz3OcXsKMTkwK6SX4B6J80Kb9Rd1D7v8H+/LaT1vvie
cXg8mnQNSSgarxod2Ap0mYqg7+HRjoueIIPe0uOb6Rd2XG69qc+RVUZZqYBeaHuJtk2Zb33smvc9
mEFLve8//FiXAzGMFyyEp58bn3nQWcjPAd2p5IxmTayLt0aIAhQN2E5eAk97GFd8MGgwnaHHDVJz
5wJme75XcqanOft5AD67vdxJq5X99eTbZFyE9XUPt728yRRWG3QCS3lc0tetFu+Wj60nZgfwVHNR
jsaQgX7L4V0yctmPRvseatDl3HbuZZRmzh5Pho+YbQGtKwDgAZPGFq+EqZVW0V2UZw/x0LODKj5G
LPocbYKhQCB8OOYjl+ee0N3UJMiW6pLv9p9bhyxqIPVPatqSu9uOUFnCkl9s44QO/rJpJVwgOq6c
agroIoHgLHoo+PTe1LzledDmdZdVQKhW2BL3Sse3b8tExLHgJ83KthAXaqgKOAEugstfYiI8QE9S
/+IUbXP6+Zw+0ApmupGQd7poXcMnorlP2VDxQh0nRAp51e+CkBke6c2TUhQVfPIjlCCB+bO6mAkg
YOgaM2kTRNB0HgscrtAElfgjc+d07fEi5PVjGZWn9fzclIgM1d7mYuZAKCoghb9kK/v1hlz8qM/Y
ztAJJfAXTJDfYgrhMPnh+tUEEm0a8PuqJ4YQmMo0OfT0bhPSbjOkCPMlZmADYzw1U9EZ3+iz6g9v
jWJE2zBFn3OyEkaAusLNkGlvK/xEiaircUQ1eWqsxdkF4RDgHj9868RLRgSIUu4648mkv10Re9+O
zVncfTb5pUjbiyXjZKThNYPGdV4oJhpwoHsmwl9/bVWAwvRdQfuYVb5fy3h2FJazNz2oN7Kww7nA
Z16qHfu3IIidqKAK6ZuPr3VTj7i/akMQdTZos2jxLMbcbC+wRxqloMzpE1TrWdukwumWOd/sTZWY
3walwvKnlaPzMsxxsnCR771SiyP+AQyRYaOLabY6aMcudSGdIuD9FMAoVH3Sa23oTYAppOKa/BVf
azTqMal0V9XhdOjo1OnE57oGNtxqfAmRXfHcPE89Y/TZXk3lBpAXVYTiEa1+ad9pAi5aF77v8Far
NRnH+wkXWPx71ySOunpUbr246GnttvPEuRpAmMDyQ4owoajYRRlXXvkRZ2g2u03EmQ9TPlJsD7TB
HnlTrlUTTad77MEhviwRJSOWPL2Q1LQT8Lk1iahrVhsec548I6R+0fs24hAJrCWlf3b2O+87VuI/
Et1YkIJH5JhamjGDq86YjKHHdLNodruJaYoGXMdF7pAlibCCMlZ63kCNZ+CTl5yU0U0e+i8tgCPl
1JiAZr2lPmnVdCBQ0XrwGdo0BmLyLKDRYOuvi5pgTxvRhV18d0gxp6n2di23WUanuFPB8XCkG8Nn
qj6YDz/fJvZg4hBYWiOodXMycWX7A02hw6oezXTkoRV4RYBDstNmToAwkiKR9PtEi/VV8w+5ANoC
QhWUhV1IKH5M/lLEf/unIYp7Jd1IkY/1v0JDMBM4yf7JWT9FiLA1KZaIiyV00GwvZZ5Bfd7HI4Dh
J1hNFrdoPqFA0r+6XVojQ91s/vudvgUAkR5gHQV8LZb957t2austOkAdJacHJXcUc/HIF4LSYJkq
kHwx/DANzP4FJLxzuFcQnQrX8AEFw807MsC9x2wFnfbuxWO5P/MM7dmNTdfpUUoPbHmc7JmwnGxj
cYVCjrUgXmW29cS3E1NXFrmeXEHLj4oDrkwgdUXe8WKUVkg1DHAG6GBmxX0H7dFV6yX9UsyFcav/
AOQvGix/hnnbVqyTbVXCSywSobPGBlvqRBkh9VZ2EkIZwJZGCtKiAty2qXGS208QkS90hx91kRhq
LyIKmdlyTWzHUiMzufomxavOKqRsc1AGvQFCotkHihTk+h8+mB2avfLtePfy8zekBvxEOY+NiRY5
l7MhFX1HzMvDqIVJWmu6tEI7d52g3vUSZJ6+kNByH54u6d1ddQFUJxj+ybA2vT4JeynCc27O/dSj
Rwobwzi7c9oPzQ+18UF1BuscU0IWtswrr/RuZLddpk2uKsxxZSM1wEJg4eX78Yjk8mKZqFF6VqMc
awt5zSPeNT8HWisSipYHOmc8pJ7nbaDl3tSF+HYM5tXrEV+aVyxhrgtpplJ+3ta/9Ri4TYZawbBQ
ZnVEKL5JOocVppzD2B8/l9cIyMXF8XYe/HGFu/aFgEoTQyF30wMn4kUe7G7qP28A2YzXHEeg8MED
Avavogof+OTOTvby4QL5HXzwprhrtFzRLbZ0mfqDCAm/AZ0tINcCG4gYShQTLmp77nNCRJn8rzdn
S0BPuAL0mL4wH8US89Qdid2SeTRv0wZ6Dcm+icAD0vdc+AgoM4E0n0x9vpUIYJQ32Y8t+8KdL+GO
ltKxwvhgdM4DM5OTTl1qMwTZzB/MSPpc/n2Mn0PrbNhGC9sQNHyr4YM+olwXCA5kCSgwOtCoKDeY
y8733XmwiSR0Zmlo1zkhAtofDbVvio72RNnAkTP9kT3TfoUDgUIDlDiBfPAuG9z9L571ILlgenlx
Y/QHPOQ6HOQA3sBICmkqulKBUR0b5W9D2XhLH2EdDDGz0F3JWRw0KUY4guSPxmqq5Dhz9AMasiWu
vW/KAFR5BnW1I6fprm+gx+ugdJOwwYu+SsQFxQQYJQ1WIrmlHL4XfVxqVk7/C0zdRnR02zE6q32x
pIU4Fh3numH/UCA4edOmdGAGqOj4cEyExlu9OeWh1yw7lsSxS7yP5mtOYCaXVaG2lno5rkFu3S8G
czBsr8EcN0+NHONLnL9PjJyWqTofhfiksAIaPtymISJZJ7onmYjHMSK878ecVayIf5nVn36JYW1+
rX9lDWSFaf4HZ0xLLZsGCcBnyl4wUhY9Eu9623U3pIIRWA32zUVgR/0dNnE1mlrSHM2xtvewRHy/
90N8DQOqw+VhhdQY/zu3yRK4D3cOazcNthThqlLEPEdfGO1/RmfjFg35xJSuQM3FQJM7MsWYiUW5
d2itYk2R9eK9gXmyNouf2uMIBb1D3g1+xsSi4/MLFJQ6BzJ1xKcAgzzb5H+TIk5MrY0SknNmWTu4
/BtICRHSE5fNr6j7voQaDmHu1v0cppDZNwMk06dNpqR/Gq1444UvqYrxQVbFAsgZhRjq/UEt7Okf
2xCc5PSJHaA163Q/9iYQe2lux6PkQhKlY7AXvRHJXbXxa8Pvr9uHnf7exQM+lUl9hxlBUpwKM+eQ
f9/cw1ko7b9pQR4YEpmQnORKhwj1lcMCZkkkVP31ccLpTMkFd1cJX0Bljvy29pdu7ynL75mjJwwZ
DZqOOvGr861+z+dNDxXHOmNCEAXPi2r01GZyXxW8ZAwJeUKdDEV2Ds01PSgvkymq1d98HROzTfw+
65hEplIdgIMN9Qy6gs5iQKzwB/SOP3j6ce98H9z0kSvWu6HMEUD85AAJnYcxF0HauB2k8azuqpOM
4oooueGgtTQrLg1q/EVY+AJWdMcQt60zco1VN3ZxS51nqLIkRasTCW3AI9Kg2e69AsonbzIVjexZ
5SntiitSHWY0XdI3becM42DP5e7d9Rp05+WLvg7NJSzDrdNaM7iO9pjqLLPnxYPfLsBZXPh8/6vK
O0z+vQJQZjn88Q/KczxhWmZTEvYh1uqeAAy2W1jZq8xfsveK461gmMFI9iw1rfXYRTtAU1qlXunR
yRTqV9erN13nfKMI4deT2vPtzKcSCa9J5wo50spUG8Z3iSgg6M5pRHKxXQMOie4p1O9PXNYX25XG
M6kdE224g4z8/Ps2jssj4h+YVwE54CGJD4sPGqTafiy79wd/TLxUgMBBDW7tngt4aOzqvEt489tv
puHLN4jyffk4KhU0/UEIW7sQOkIj0QcnWzgnxVy+bJbP+2YZlrJFqNFT20xkItPRONa4rUTJXhKs
d7icteZt29/wrQy7DJTup0ZP+1CXz53zVYLlymLm66RnE4swQcvziV2PszioM98sk1TvpCN/TpPV
BI/nJL5Y2S1mWWypSDoUNJbhAdFH0s85PGB7806cC10fZucQShkALPkBjJJs9sjo2UI5qzBMoaWG
C4Ra9633JuQl//pnE79FmJceR/mP0nILiJevVnLEDaPIokt48ABK2z0I3QLCcJG6LtLh97fYCstU
p+t+rrR3UFdTID1BbLCWPlWQ9rnX6JO3G1OUiWw4huxKciUaq5djGN9X/bY85uhk8qSvMSw9woeD
QyHvD7V1wcuOQTaBQNtXgIsAXO5gOMybCyNEAluxvRHvzfcZaOI4yAHHOuRiEzJr78hgaz/NUjDi
aAUDTFBdiG3dsektwrXZ3KA/6RE76ifGRFIAb6sv1dT024E/19U9DblubEGcdPBM3EWTEo3i5GNh
lfpyLflcozBXFKHItgqK0DoMRyR2/AJHx703fH8M2AVM5qKSzkymHWUwj83MFd7oa/81jY9p55La
usGDcCHMrXvP9nlVMp29GJFOvxr4esUgbGprfqN0OzC/5DOvgnO0NDLLL/deFnYW3BBiu7Xgn4Eh
r5o21D/Y2I65stpkQL9rY01+pkNoE2C+mTrd4SeP+qt9njODuto4jFb8R61/zElvE0Wl8s1jcX13
sYDZm3zIO/CbZSne7nqOiSOYukWgEG2NbSPuK24NDPag5gBtVwCR27f0ko5onPYyM1acR1XB+q1X
B3ozdRlXd7UKxOD+ZW4dIjo5ak/7aqFzsSwTC6nd33PyRj2mfVOcQpPVSJYuPHIRZYv7GFmXs9BC
jjjg29NExZ90UpJSpWEPd9MiTTg/q9WTLb0bChFpxfqn+XNtR2UIC4y9wGQeWJRZF7cBIrsArNFt
gH6aqwnqdwwlPBO3oiWiqP5tgyy9wsIwTFR99khZAKIth/8ppDJODvtf8PuNp/ZDET5DAAHf9pmq
Bz/Cbc9wK+DN7eMPCFR4D8wqW2QxCFxLLt5BrHP2KV16AIeiAMhAOZHN6RfiQybbNmrqcxqiBraL
LOY4POXCdMxBKGxe/wi+t4EQ+wjdi9L5OaMaF2OYuPtG3o7d0XbENMS1/XkVAjqc3K/UP9gD1e0P
B/9bSowOv6NOGz0YHqQI5eNUPcEQkcgElCtf7nFJRupmlInSBJznvQBJqV7nUgJ2cjcqu9QTYtur
8KHGk1BpuxA2tatCt2LjVel4cgFHBCc1h0r2LQHPT7nyTKlSkJNbrakJzQ1gzYGraSUvRPNHKyXE
kZYwonfC72LdBzs5tM/h2sNXcLJZWKb8fegK6dg3qK/UMfudDsBk9RUUG8NXvzN55iR0OHx828dJ
7Dbtn+R06Pdbn8+goGNqtQhk/0nwJapKcN0eEXsDblxMBwQFP4zlPOt3rsfmN27wqvWFXxoTjt4a
DcGQ76jHXE5HVwjdXYtcZsnYExXGvR1eC4XqXEThnI6rqrY58G6skqKdo2v+mJDErNT5S0DACZjY
ZxQoUlo/fiy5C7Ve5OOP8XbmZrcx8FcodYlc/rLhDyTBJxS1yRafCS1rgE/QtcyTJvBuHntchNi9
zPOd71Pul+QInwMEwd3Ki93WnD1jqiQiCjcGGSEpe40SiPGBw5YCexBa8QfVUbLCyAppochBbWC4
xTUZSos2DRvl+kbB2lAO4Xqdd8rYUgAbs6YMMho3k9DnJHLHEntQq9sBgktLxrFWbkjNUQ+2B388
9iPZ0iaow5K66b8FuwPPVjoE8G5PvpREDqcopOI6tFtJ8yjbUuJUkg+exENLOtnNRNN7L9J8hdiq
0Ke0MY0ujv2L6//2rXDrzxVvR/cNIbZagwgbtx5oL/nOofQhaLrOCmzw1eDdqzxPSZwvAKBi2F0O
HAKHm8Kld4nf5dgeQoF/pKwvN7cbmGb+0H7IdM95kJ2Qol/yBAXYj4mo/yu+hS35Vs3BrftW05PG
B60/m/DS6KpceNnfAA3bzAFRyoQYKmLzaYRTmk5XdUP51Z4OxQ6dN2BrGIgLDHYUJP6sgJcP4c5X
Zf0CU8cnsJNnr/UkB236e1YKErkw3GvYPii6NiI9KVloq8tIMz3v6SJGg+cJ7uD1a7TOwAR4eir4
zHBYQ3Q3F03do8jKEEgnhqFyCfQev3blar+7TpsJaGGL4s/pofIQoPhpHvnhs5RFSmGrRHlxKesp
wqQH6qHW0bSTsdoF2DnxBUpKwQlOM5mv39s/9+oT6hCIIft0pyU2rz02ThwT4/h+2jvPjTrR4FKL
jtfwExnw2vgykohwzdBx/yLfN5EDzFeQI0HLS0PVpJTo/BzhGfhqOMi8atI7FZ8Y+4dMWDb91fRz
FkFaR1HMbcJT+OHSD3GKq6tzbGSQoEMZ6vO5BJXLn7MbBxM8gT5dKOvRBcnEHTiRCMgJ1MDyBn0o
W404g5a1lTHfh7jLccJVdzNXIU/1+Opcf2+fd4FHrLuSiZviiLzSCICnlvra0tqY/joLeYIaySrk
phNgqrvKJ4SIJvgwpeTUA/kMG+TEuvUKFlYaIq5/E/NV8L66s7CcyMg91wTlvqn/Dc3RlAWpt4CW
7+i8CdLUEnEm/H7OzcUtD0T3sjxxItCjrU37wRf1+7BnNv1xgRrry7P32JZJhYHTpOenN47eYyc/
L5uAufmoxevAdSsg3rG6PSdveptnfR07IxOvNmuLZEWFN+Emu0UlaZlF1QX0dQkGspxqnSd0PSVM
+5M3e/sG5FWS3VMGBaEVHeJtiq4lPiybRSLez1ydkflWemEUIMzrYxVhe3VyVLE1bPjAk64bBRt8
fA1Eu/xvoerkpyhvo5G54pif2qTOq7/R0XkcNaUP2+OqIpVa/PTQL2k1tsoYcrr9Z34vDQoCkgU4
4u5dYBBF4zzgYJDuWkn+SorLR6bdfQn0WjBOat90sb0LGK5kf2QOF3XepUaiom86+ojJpZ0wGS8o
Eb/BwvaSgaZ1CQQgedeelHfIK+CZiomueVj51TJhRXxflplF+6zp0ZuW97E/CbFSLAA0SvaKS+gp
/Kt0FmySM2MLroSaAlu/FY9adLvNtHRAs7pmXsm9TEm3bIiea8EQB+cHXcBCedigcjGJnLc11FDq
36+OvHbz1ULITM9e1waP5oOso4j256YpDzxt75XZFa2OfezaBYK72YFgLeTXsBWy02pSWw2zfo+o
2yYTgtsqAaHLo6xsCa9Q2xj+q3vZtmSq0efkokD8ri6LiiA/4d53b0Dir8d6dw5aDtmQnU2pxG45
rjmswBOy6+/VBmJqaB0lVnQOmjU58q9exxmKJCoDPJ3aNwG1qc/VQiE+Qo2WwThBD1HKldFBjZKq
JvHMlI0pAJsFgrl+AF6vZDqYaxXqrsrviUQp7+6HyDI3NI8X2DKUOj0BAZfb6UsY5rBOZV5ezTRf
GKdp1SifxdQJtkrwR4yxh6AHSZI1LUletnm2m26j3MLjU+YeHheNMt/j4dX+s5rn2mr1os/Gl731
od9tywTnqLIwB39H428xaPmvf7BonRwVrn89985bTWeqtz8uUIXWvkhXLPVBKUPP6zV7iS5yANpD
gvwr6EQQX+dmk5n7jKqSlSCNOYNDMU/1xluhuNKhJvw7zw/m77DGDlzHjCp+172eyiYMNUyitulu
ZgW+4VBzqYPPhTy2oOilTsBaBgmz3ni6qYyoRqIUSpL55btpMR1blJrga8mHCB5ymLdoo/I41PO1
xR4JIf/xraf1EnO8ujCmJXKgfuRbaJByX8i1JhgffmrrA/wNR+l360lnzqAjlKROmHBbzzXAVJ++
0BmPzTSGU8iOFvePV/Azrloo+ek06IOTsEORbMZy0h001rEwGOUVzalxjPhEljqXxEsSFVwq6rXa
gbbRUmaJBSgJ8NHWjeQ1elnaYrx7qrdC2focQwz4rTm7bFu9Vl1BN+AB214WRIc0nMaqS8ryCdpK
1Tvgy7VI1Q+ZnxgPVkCewyvMtrm74Vk8REOHrjzwWD+hICbUcrWdUBg9iPbs4nDHsINJ9VDHFjK/
VfiiNPVp7EAeZ0asTJ6axZnNfEg79akNay/efqz2jLCdvBS0vCUSFhv9Am9mRU3Njck66HSzb8AZ
vke2b1OcX0OF0OFSXRW+jW8HWwIRZyJs1IEemSlRnqanaDUnPjQJpmsUzK5TCsPYQXr0sSQVz9Ls
RjviK1DWUbdJ376VY3nk/clQ+IDlxRDu4hBDw0ZKtJO18wYk/bQgxEVivOThlruMNmZ2w4WhlQg3
D7X+/sbVTb5jXK4pZjzYLjoKUtviuOYloaIjvrUT51MOBv8dT6ivmRpufABxM9KL0tAF2jy/S4zv
VNjXfTvuPv0xBUadCO/xTRMBI6+bHfcamlA5LDfkm5TsmU0yvXOUrI9fI+sWEY04hUX1epZ7WGSR
iexBuYBr+PQs6Eo9kQ5xQvZv33aIsx3G7T0AWaJseMkS6NZLBW1Bw/0AcCEtPVcuPqjP+129iH6J
8eE37P5FLRNBR7ufSZgMVyFOpZpPK/PfHiOyb2eWamUAxe3knCK8tX+dg2rfkZQW+M3Fp8JIj0GD
HezUeMMGX9Ge33cBua2pww4VgPzDJ+QuJ2qS+1amWA/tOC9Z9a7wqMgbQBDvctBhE7ztfSXhkm/h
fMokrLQnD4Mghv05P/K2T2E/nh0a4xWNvRfYZngU+8cCgly5xM9FbubTHhZ5SxGrICUKYHJ8Wup/
yv3IUJprU3HwrH7WJ/FdcZEpDj4incOejuJNE8wuj3aKg5g3cxO1+4aD5WfXGPTdyXFX8onAAY/8
AxCK69oDoVGqcwRF2+NP8zLBf9Eq6Inyj3MyRvK7za8/hppWMsVPvb0+HfFdhjQ41ev4OYRJZdSH
XZVTtzmBNKD9QbkVnckLFgTXHuVzVFDjmYbFyYQBw5WAr6ydNw2WqYW/cwldD21KF1N06n93gE/W
ZjT+pDAUmKQclt0NV257jMTOFw5crbUCI40hfyneAEKOYMjdCUyMJhHkIGCd5AIanfpQBmhe+jR6
C14ccs8nxFMQXnoDu8M6/vOABCqdTsREeAZc2aEwFe+FUzXfzSOZkwTHLC76Ki5305sH5rIhqE8F
dq5x8r9mkpIkb4x5IyyewgapHPNwr0NbCHrMmiKa2dk+BjcedsrKnSDjarYmhe94M7y6epAs3Ue2
MPzBcEUfX/pCSrM64ZSpqa9Po7IgU+d1AJYCcQr5xtaV8vzlVgr646ormbEMWgTU8k29pOA1E4IK
nUbmC9AuHMYEwXBSP0tkc3NIuMSExrC01TJOYnUE4SbhEgzgyT5/Xr6UMS1ndV+3ofGVRDz6y8cy
axiZi1QBLF0WA9uuE1fkfq4Db9ExFQ6lr5Cyrr3gQftBwL0ZpGc/UQ0B7Uv0Z4WZ90YsEyHJWepQ
aC7E6elgqBMR7CZUhKPDmPE/YBZ+jC7VsYIWLBwr14oxKnTN+ubPhkUnuKyCFiJvtBBT7SqxwtR+
QzvuaRaD+fOlcqFrJFVoV890kNs41cYgAQhhGTDpDCnTohBmRgnGGLnHN3mjakNcb5lwzjwyDq5N
pj+cPI0m3wVhBhj60mvdaJbsGqZm/KEBmvIL88ISf6ll+MFGfAIDQk5EYDCg4+cM/nq1KN2UcXps
DsgkxfFJ0a8psXO3KOqnKA+ooo0DCEXqRt+Oj25hvmcKhWnH9Z5wDkVEe7GuP3TL4yddwG0ssNgJ
hI5+xUwtWXTOFL29biJlvwBPEPI/H2EkkfWZse3GXX3/sin9bycMql2fE1p6QskO+4Rt42A4dL9j
ZLvXAFQXl3DjIUWcTOHa6w+IH7hC6tM0CoiYjHSwV++zIZLJSdBPzi/9RWE4liNbfkyJQDm/48Vi
2Fpc70rjOhSX/yI4yqjlCrQ9rrTNnHs/Ai9IQNvXHnlnbhU2xintXBW2R4/fNJu+Ul3Zpya1ZJSM
8k/meLOTrW9xFkwA3So6mIoz55kcQWw4Q0qlLovCYfy3L/ZjD2fbp6t5e8JeLiCkAKbtZFmj60X8
MwE6Q3Eu8jT2qafFFYXA6B9CwS0mejq0AaC8H3vI5L0aFOynBniyK9U2FGvVeYe3aFeHMHMVARWq
xwomF0r1Br7r8o1oRKAe/OL9fsnCXtPYv3jmFxBax38hgXJFq9eCsDdHWGhptZXNxnL+Nq9JXcsh
q7UmqFt9xe860dAPdluAcdncIJ5S1FD1cpTEhcdtz0Yx84guh06SA9trJjS5mvmXi4fubZOVowei
AYR71dorqJJQb/8JK8KbZjbVypzQOwAdC6XSDmX+DoCxXbmnfyj6Ctiq4qyyhpGCVIXYxVJ5xhMg
JcapjmU1GTdRCkMKR+x4f0934LQchUXGqedi3rtFYcuTd2e5vlFdmEtEVZUNM188LErWhgXH2isF
ac4Qjow/822jgoU55OMJBPh9vDquFhSd35mf1t7anphSWy7cKZdxjtT7Zs2Srmp4qrNRpayOaQNi
s63TApOM3ovV7hXNzt3K3cF1U60jdxMkIvf0UUdTUSzIBHDrjZdUfnyy85FjNE0c+EJ+1TpfhLtK
goiaY+xn6RXqXXamq+bYvOIxt6BkCxYArF5glRVuH5qKJWw04r+/s81o7VLHnuijL04PE9akr0Id
Ovdnjif9FlzqdVAih97P1FAFZYE2SZ671orbrIGUe0LUs7ftkNDEx2L49SzwUDr8nZ3awMsIXWpZ
1v+IgheXjSCgbxqXlo3NsvTDjut2gJmRLqafIuDDpFRbKbXZ5ZUQ2998i7cwsxNSLmchGDfhrY5X
HmzFr9Fg/QRAezx35GtRVunOqozrpLITMmjYC1Ilvgl3tLk0GBTp9/595t18DYq2oXjJmmF9RtF7
3D0t+Y+gar4vL4chOdIw0AHO69FxYb39QMP9mTO0MyE3YT4P14St+1qdtyyey+oSIjYWnck0mAar
tDrLBGTQMvh9ecV9IFKLTYpgMQApSn1rwMurYpaqdtzgTD1BdRaETKLY+aQbNJyouzR1qXDt7oo3
0k2qQE1ThTHK424lT/8TA2QmPtTwDjabteRuRZK+8CLAogiTqZIY8W1C1sLOAgAV2p8LKMoTJw2L
T7NBHKc+vmEfgk5uP626qelGA+KNfXrR9QHvs9jAx52rIkzhpMRFGld6nUAT6BWdmqsuoXh4Kz/Y
t1bHsezUV27UhpQT+O2Hkuo9EoWCaA4EO0e+GUY9Z9MzvV5JHWkcVX+EjJj5+VaSviuHHIYS63wU
PHAjAf4oDjqF7ZOFOZM8ZAvbPasEAEs9tyjM1Jjfjk3gtaTgcfNpsZMshOZoflLLSVrbT/J8ZWyo
HVZbYys6GqwZRhCwWu4CcvZ8JtnFnvKAMc3N9+OHkN7T+JBn8wqZVCoERVkOqoyYKwSlCVqp/g8f
taL9eaNVIgYqgU4m+gTcc8t8TVTnHEhjar91nOWUJHcbpyaLhXIJh9DY2oc6c5qMl08M66oWQ6WC
zNs3ySvYXFojx9Zo24s3aXRUmqKu7otjIuIgl8dCb3B02b4uCDkMDGcu66NrNRBh8xvVLEJCVnRi
d1/wAV+Il83YLsTx5N6bhkKy9ktJDj/MyhFhggiYEokmD7lh65EoCijZ0DEQN1wf+xhZkS8S4310
2FE+NmQ5fyQWAMx7bCtP3Du8pUfDHtUfXs4cE1Sd06/JoWEVqBow2vuZ/PZ9htOy8BnVlEOjnkxf
V8r9xRjbnY4XHfcpuD6czTDvumOcHYYYsdHhmin/4V4QHldN4ZyIdqknjAzY/hnBwI/EBjXfpepi
gQ+LMuEJ8HvdTbwX+N6AebNAge2glsYTcf2EHdW3EGPa5/okLT9A7HPXdwWwyTVQpSabHW99jLku
6jD0RTjdyExn+VjknxTadbN8UNH0cKV65Y6f3K/c4Wd4E/9fNbkj+oHfaVi6tjm0qJunYoh02E60
+R71uPUw5xagw5o5N6KXJDBQkjpnj2PkIe0eVmH8nLNWLs45/8KZj00qyITx2zw+1UjZvP3us533
uZXuUn1smkj8hMPU0eylF6n3A8fnWNK9Xx/YEeNqCNRK/f9JjMvUlTRdYcds4UdpdbIiXnb/PLaX
RL7LMHv2k5UCc61z1F8fyz7s4JdQ6f4C7HpRqq3B+cogucImiS/knRwvfYruaK5mGhoW2LJC4SOE
Pfdu1jfuYFgIKRhYHIhAjwSXdRlMq8NJt26VgU41MB3NyhwfE+brR/6yfNNzxoJ+Rp8U0WLTN/Nw
vNj4zuUhHAvaGDZP0EKhcoI0b5RmBIG0rodS+QKyvmKmBdhyF8XBGZmyL9DnwMJwNTVjZkwzEZBo
kj7jxAQaI1z2/O6s9WqnsuRgDGHVR9KVfwOzRslmwIkyVmcuCrWPuAI3oz4cFBnY49SOgSiEQBlC
T1xoapkd17mC31zQJ5HbRm/Le/yFB1PELAWP3Zgu/yNk7gLj3zn7CX7OApqi3qTlDY56HgDLTjSY
x0zn70nFf34N3nMTXXAp7eL2ZokX2g6qnF37/FJV4QvM+OEbFA9oMbzTWd4MVqrhQ7dqRqDWyGuu
f0B8+FHVvtxu1T3rHYDSvxxnk/cC+Hj5RvuUxGxGLIBHlIKshvjLsI55xx3L1qvswqUpmeNbWTqp
2QkHrVpqqnqcZAUpnguIMSbdmxHTskw8OUx6N+YcKJIfYISjdV2voVVIexbTtDT+RNGQdnJiEAiH
3wCpX/I9RUJU8F10wlipp2qk6DSp68neCIrXlSJp+r3CZ/REhooBNgkvEkLK06hoiIqHhz+atbWZ
QIynIJf+RiUWQC9ihA0L2gwFKQc99TFxnWmlfFLDiFY+x8JEkwvY6PcJFI75MbLL4VgSxqgqS83E
IaD75Jn6NxmCKtpVx7PyKLtVmzV4vtAxd9AfR6xAx67gf+Xco5IXeUWtu5aUVSwk1WPVhNqcxR7+
64QZv5sOUOXBWoTCmHzHPVmhHYVcp294VR9TYDbwS5h8bxqun2ENphea10G/lYCSWd9EEeAF4gHt
fWmm8IfZoGtzutaLOmzkVgJKBXfMFnpx8SCtNkmHLbdd6jjkBYez4otxqrgATXeJHkvJsWVWuZOT
gUlcggjEDqOeWFebBy4S2UoDiG8j6Udga/c2ji9P9klCP7VGApuHFLr+h83Ho25/hI+B9K+pTWzp
NhdcVZY3tfHHIE+2MpFxP6yB32mWfrXkDXy3bB38HIxlGWRm/XXJ+7OrlE3uLYYElYCHSPScKU+U
tKZOvk68GrBsbnmaNeUXbiGn6062xaQS7y7XG+79mI1R8/sU5yYdkS9HksvGnTtJCR9A1kizG+pS
zF9QEOmfomWa08hZ7bfvjhhVt5OwQQdFmHNBFbsjygm5AJHh1hginWq3CA4urHcOYR85s0zUaO/X
kL7MuwFXWQydjQhqCDCJusfyka8E620ahkC/K/1N0ZJ0qK6XBemW6ikc9/j1uugHJRd9pV44MnOh
CtB6mITh1eG1xII7PaFUgCxAIrhxB6Bm1CV4gstjEO45cyaxdtCKceQImv202/B+RI6RFJpq4d/e
Ad3Qh9yREKhqOUcXsQLadNILJFNzqn/t5atAro/wMrDupFBuBqdWHyo2qgNn46gStSoasBuffg9g
n/udPD1gkoWp4448Y662v2/0r7jcpzs/7VgXjoTVqlg0VYd1PGoQ5wq1Yf3qcRg7vtTXG0mfJN8j
bgZgSzQKbg1IBwrzGNnE+yaiTjWajSaC3y+PiKMccNodrpnm1wlrF+RkiNulhmoGmjWqmyL5BVwq
4n+LWH1sfsGFRiRbhgxjQjK1+VQXksPYwngOJ7ifxRS61cfpHijQTnXyTTdiNHZlyfemPhzuRka8
hoLPii3JgVcjuC5Ccp0PvvcRMMo1WdiVNE+KwnB6TIH2bwK0yKEjIofEgXN9HBgn6TJODyMXf9kb
1jcqmENfanMP7qaXtQb+JLSNoVCL2PCV4jJuVRylXFn4zz04a+TN801MPaWs7j73cR6FE9WZ+qak
Ebti1ldikleF1mNywdD276dm1w69iA3ulIOAjPEvwR0/AWcNefBGcXPVJkhwVreDehujAy8EBVak
p0SwLzZCZtO6Xe+kbGEYrPFY7zz3lBjNAAt2/fI1kJ+a4HVkHjAxVEAmq4LmsV0c+V0q/MWB8zoB
rGIdsN7NNL3uKMaOVIYAdmw3yY1P7KKXxgxx1Ymh3Uj7G2r1jolAACtTDSZf6xSy4WxkpYMW9z8q
LDxjv17PSaowKjdIYKoLH/NITbB7g+3wT+QfVXt8wU6JUDcYe+X2ymh+EXnRDbARNXRFv04KpY2C
dEMefDI0q72TrkIHmNY9DMVW0ZA80CPWQkOMBv3Yow8VA8qlzCRykMpfQSkwX54M9CT2b2m53XAD
DNJdWsHoeRj0jlG7IRYuB70G/KN2sFWD3/DRVC78X/V0vdR82XHeGdgYb1hDTt0xoGscognfmYec
HGPu2TVZg/9xcy4UOnd3cJxt+tsBtphtOaeBJZcA9MzZ/LnCGOdUD1bM4yKUKsXepTN+ieT6bV61
Gv0z9KecRBly0jyjXmZJjmlGp5oc5ZnT9eilQEWybj58US5EO2ifZloKyilFX3oeSU8HHfT8+uVE
H5hsIbn4c5DMYwjhLbQzkHbIXuhgw9tSH90CvxF+UBtA8kWdp0T0Bdnszc0Ii9Rera2/a+6C83As
Tag+VpabbRKObKy0BF9eBxBIQimV9WG+qx9tUdWJJOF13ILgSyCzTa/0Sn7eiVJT5Yz0D9kANvvo
f8sgY74kj0NZYx5f4uf9HNQVTnEHdRs/kIMomY+moqzemh5e9nu7u8vdXzUz4k08PqgaLBcuq0iX
b5apc4o/NE5FUFQsPiq9y7vtLGrJ3RyCSibM2t0++4cFrCERX6eN974KQv1OXPgK4i/7royCIeUB
AzK7LNyA+GgpfJUROlEHXP7EOP4YZIYT5EDOt572Oh0wWoOafjJAoG2k0tHdjdz8PtLDza2s2x+V
LPU4PqZUBgwaxPkn9g85f0CR6wBViS04MMr8ve8W05Noh0HBzpy9Xg3syq2uAQcUPHKW/YTpLJme
YDdgOmmARuaW97KHd2HnECt+8Y7pNJIGCePwxW00McS4L6U0hDpqecnRZ/BIi2kej0EkISkXcelJ
lbJygjq8iK6avGzTWYMkE8hlKaaqndaXi9gIL72ROnVbn/E3a053yN2boCAYiiVx+RSa81ZQqepG
Ls7p9cWJNybD46SEGzQSLpRm0nwSdPTBqr0M7soYt4szD8y0dTUkzVKi2ENlb2/WdSnkQTEL+a21
MrCrkeUL6BPRTZdovZwd3OlTs2U15VYD7RO9xYw4AZoE5ajnWAP/HJNXU52M+JsvD/LTAREsdrzo
m3ROV+YmwFd0GZPkmt8hjWPhTW5CQXtTHIPtM4oHfGvu+7Z4cC7Z3axFARI1Hx4whkpoRl1R7xid
XVXDVl4dhfjD3oUA7YT4Ox15vEd/hFQMVoiTB8cYB8Odcn2JWH2hGm3EcBXKR/MqNTeskyWOg+Vq
YKrmQb/XuhA4tzvUr0N/IJMG9BdCpYFzgyldwQi5aBXtyhKzlxl/gbToVFCavTAqqJMba9JmcTeZ
NWxT2s8UjRnqgj4fSTxempuBL9w2J6aWgvUy0d9aisjBq+3XgQr7CsJrG7IG5I5xbGAnW0Iulf4g
GiF/EvjH3+gu4d9QBeSUUhnaTpjW/XwWFmThQu3qseKAvp0sngsrZTYDg5ZUo+C4Km6Gdon6r70w
8l3vF8rbgwIKIkqXxtKWcpSNVvH272T1Q/7nUuzxAtD/PEABvTuZ0kkvHMDMhQGUBHPjWNFAo6i9
/fru1Dv3sinG70NlqzMFfSeVW9HMDs5CB6T7IcSsHAhZkxva+BrRkXQDG5Cmf1zrroj9kluFc40b
FFivfddHYTQWINoMTumc8nU7idx07NN2NbmA9YubFpM0i+uXsAaCRdVx8tD7UFsZDzZsglmG6RBO
VfHODRBsCE8q+pDaOEmA6kA7o9HIyEHhsTLZTvsqGSykyht0fgU8tbs/Bu/rDEjrF+WzsS0Az1uz
rW9Hkbr3ba2YWgWI37pJRHOcImsgYdvDipxCVnqJmSUVnNpT04p89+yHIkixWRjkdLHGl2AAq4k1
KPFYUaHFT5HXbf1mBKqkkQOl43pjV/rZv8iQVaozHU7RBZYWs/Th6dvlWlwdIZpia/SsZcpGr8//
AhZPic1A2NiNzah0AsLubYJqCpU85anMuwdJGagi776jQSgW1NIdosapF+rPtVaOhzqYJLy9b5DY
6lHWNVTmq5KBwFjTkJzUSxlPp0a3Ip3SSJBE8kpQuz2/Gjrl6fzfKEc8T31s62HnAfadrS+kZUTn
znVkzNB14RL6UksBFTnAfmhfbU6DWGS0CjaRmsi7b2V+gvOQafsug1haVCcoFayp4XjMyMyTz1ko
1GJOeYJg4Knh4KtBPogsY/ElsS6tqn8RQU7hr0X3AqHZEac3otsPnU+LxQcg2wfC0orr0yznz0Fx
LNyFXmiFJB1u8acRyu3dNCzkuF4mPqJlPPYYnncVINkUnGhNBVIMDqeP+PeSLrgtPf4RWg7crTHD
DTnQubTu4SXtgDe753nvVnap3xJ27UTJr41sftJxPM2f/JvHr3RW6nCcHDctlB3oOfvIY+3lk/rs
oJZU5tOyt1A9XctzTXwYj+zJHl7kiJxOIVJdkDfJdp9zkzjsHrJ7swt43CN2dPPikCdgBbXXFbDk
G5M2nseHxYE6JfQGAZJUg0YBIkMF/mY0gE5l1alOF1MfD9gMnrg4dRD3529JOAnvaqqhvcwcGC1P
0f/qQnpdBAwCv1YFYJ2tOaSEhuc7/PMoWhS82xCCkN/ztmeupE0tRmoKE0hgD0nmyjmx0VyNYLbb
14ZEIoS8A9pDdkgj+20xFjci8PswKvSmny60yD04XaA33T4I7hUXfSwx9ufwZHg5M1XeeyH497xv
nVhzIZiWhTT2iNcmqRbXB5Jk5Dimxsm3XewOZSjMmKfVCq/QfN9No4iuHyhu5ONjNuHgtkHw2Z3M
f/ocRONFM5P/bkPzO99pQh1mhrQPChW/SN0CXX5fiNgwclzqjn9t/BObpfbo/1UxiKdKtiXq1hOy
7oa5/QHrlPvBakH6foBs/9xAghpVIz7VeZe56tp95zfY8jFc8/kG6e/03FEP58VijlUDoek4Awmb
/JxZyiQk1ck2R0XBZ6lZ2qXQPoLIzc0mub7/WpJchIyPdiwx44W/RxFkBJh+j48RMHYd1f0g7KZC
aW7lmN+Jpn0+7LZq/cujDj7Mu5d017dzsQTa+/Tf5roGh2fMuXc+YqVGZB1VhPXcgH1S4PYZ7ocW
1+RLyvdZdp6eRiICmt8DP4l4SK+6i/re8BaExGVN3N92OEFA6xMCVw5Klq5qxRhG3HSvXPRLwThd
MJb7lKP6r26HHiPFC0muuBkfkoQgHwaKyPmArSjr23o3CxlLs4oB96z/4RWLAmSjZkMF5AsHUEfj
ttar13cHFh5qN7211oqTItqRi5cR9saQyAe1FlPJsXfDOjrU0CD9xlRvRuMB6j7azfJNa42l4ym0
s7cd9jWO9HwEGZJ+KL6LkkhqjOh0EM9cpV9u8IKNd0qac3w/CNijK2P0TwpzYkDtSNs4MBdsGJYp
SYyW1wj/CH0ztOD4Nh5l7inEpcDenFL8PXQQ6KkFUHgGwvh2LcmGnEK6ULdjN47feftD/EvetJiZ
2M6AOeSKaeN5Z1fIIDXpkYd2cfg57OC3DgZu8h46BHtFkLSffQTFigxy+LdmCpYJBlifgbH//vhN
sJD3F+O559i31SmTeGGKD780wE5+KF+Fa/AqgmMdOXe+Y7llJpF+qAv/3geN8SzDGMGqJ19GEof3
9hZe5k3cxnDxnc1WvpimTCjEB2yicJzFo5SVRMeQUjzaowbUp8U07WutGrFNQlQv0u+w8Lxo7dQe
ZczFxbtQL4LSHHS/pvizAjH8cBtSoEgS/fDK4nU/6jOYV3M9KoYZQFXQGjtgtBrioeWQttAvITfj
EtQZSjojZEgixiofrgQ4UWNkd7ZM+6RF8S4bE19D7gNB+AAkxpn1/mipgszDYtPs9qWecp6C6CRt
+UD/PHLpwVgbq/xHOtIqfOowOtCxziVXbwqMozHd+TSGFKJTefQkL4lsj3/ovJfwAHQO3vdw+UHs
lJ4AfLT1q3FzdsX31vjBg6e6E5C1SpFsD40VKRVtjnd4GIn8zzCfRqEMAJrZT8etMYDaFBnSWv65
ds/M6NPrf4ifi1oo852jo95p0WdAfYBZV7pdgMIB74FQyxh2DNBaSSNNa91iJCfkaIfMz9ZVj/tc
OD8N6RKGyK9TYOIUihCdyAZWpf6K86ho+wX5+Qh3C+uzy5Re1buVxPaA+fmipq5LoK0Mg7J7LP9H
9UVH6LPu1fLsxrK1NYI3mrLAhadxkIP/S0wGYgATQDLZq7LsNyHg0h4RfN1hE8QXOJCFblM/YVAr
AUqLfs2JQCgcnZV8BuEW9IlOPf65pmLjtqdILNajs/fF0ofUzCm1735oFmpsAD1TEtzZXrkwBnW8
AShMxyQr425dgihYov0P5hHZt2D8vnjrb5AmVOKRxLYWvnhC+Phz0nrqD6ekAQfsR2k6uWAMxjCl
KXYaAwg1aEnV83iDof2ZeXd9mdv1twywtsq+ZoXTh9LWWEPPsS1/hqXEEkvkyAjUzm0xAWPRSZMN
TxOonjME/Ctjh/hU2AKB39iLEtztQYcF4Az1KlJ1P2Be6NRfagkz4LcCvP/gJKdjqNIlQkuA6RTt
55b9bCKxM++Xpd7V0Eh+nyQFcbsqR9tu9DEBpDnyfvbh9LB1LCxkkAUEFzfl8cHGj4FzxNeY/waP
VN8pb8JM0yy+ACMBRZBrG3FFTqI2IF24Zrs6QuZD8OwQbTkxdgvMQjute6194sOXrpb+lUfEhhbK
PJDcc6gyfHHbXQlA08dL2/jFN9FbEjXhoy4bIugpw0Zv5pFD1NwEUL44LMusIEdbRmd+t35cXK4p
5s+mQHLwStzX049UbfRsjCE+wZPXdGqa+DmfouqVMkUbYA4tyk/R7u8RAwTrQn2MBm36XKUIYg5p
Cof23WKYuIG75gz7MF2PLrxfnZW4sv0stFY5bKMJ5UUpMkZ75Mb5+r1VEgHYGPFfwH240bk7UnvD
H8MFCruTt1R52WFPFsa60zdqMuatXDtM8x24PGXgww8SabwB5giEWOMUC1uoeEKeXGl7/WDNr8m3
z642s8eDlYL8n1DEaZfcnOR3TsYO9m7ry+3P8AAyidWqk7/3QNvX4/3PGBEoVemFyjqZhikkTJgD
NoQQ5G2hoIZtFibwiqPoRkwf80uj7joVsjyVv2KJhFqZwBR7UA0NvERr5+LuI4gtqRSSOLX0RJgA
FI45yRQAPXk98E5SwTt9ypIYopomgLKvl29HmdOoS205mF3XhleJcKYhgHP3cR761dL1kWXFrCB3
tNC8FNVQmKnJTjhGT76yzZtq+N7HfH5lrEO/oiijWaM1TId1omxn5wwJ7I6hf37blqOMJlDI/BYA
CNrMocuUIAN0AOh45CGtjAlGs3AuiGgf41S48vyKOU1l/KqBYvwGD8P1vry+6DcoJCKP1sGGFd3t
NRBapdRazCMwQqDFDr7/HXJMl3O0PV3iRgqJK6ixJ2w5+AFppvOtpEicaGYViNCr2H8pThCFN0jJ
QnulYIwmTIgCgBoPUTlYWL3MTyrq/MyejIt1V+We+abUCXhZmSeJgRd1gvxl19otnXYO00ULXArh
JTmTuA+MP1FbW06HjPLC+9qfRKs+0XxeJC50K6pBvgio0ip60V1ekZGP2fYvVDVUgKckFW9Xmpfw
002meiMV3Ifc9wZuTkn+Z1cvnzxOH9STd91U+KlOg8bcWbpK6txhgqaXFL9MznnsWGADlmmhKAIN
Oox2+zmwxsJFa7OWMvKJxWFX03JRtIIYSFSfApt/z3xU4sEPShGtQyLDHtWagRELHnWAr7rx+hmr
3nLfa2gmtOO5vnrP0ZJ/Oy3s3ZEw+VxlBI86TGVoiGYJVniJYeDHbV9FUF1fI60+5U9H20nBELsG
X0bZVuC0Q8IyrvCiyvvz3RCeCoGEQwRSSuewGZnTw3bJDMuSQ5Q0COO/EhFzGLQHo/Xlb7xMW4by
SjTj2QDiRQq/foOl9fdT9z4HF2dsmV1piDdS/wvSRBG4D/t82d4oM1vjoYWH7iQ9Y0lIlf5bvDi7
g+cfyVVLiL/Ug0Ml5EH6uGe71mvgrVyGT8eZUbjsiwingkeWJSlcT5c76nx6G1sC9aC82oeVU5LU
m6GYZdhsieFJQfcQq5zyMfZJ65cuUzW5Fcuixpgr4GynKxwRWd0uzo+0/iVSH0JxXM/dBiz19NPO
R5LXp/ssGKC0bg1GeZrvNoeYWC1MbtDa2wsaWCuKSq/fuV1ZUk0WEAmRAb/4S5Ok2xHZUl4k4a6I
TyCFj/LEjzXjQ3uCq/G35HQwM9IXm9qA9eijVtA9U8flcMTe345Ed5cEkrKp9Ob4SEY3UmRM6hC9
D9mlXHVOg1X+mg31t2zlJLzRGSvWnWq9zLAk43KTW+19RCnCe30Oq5sLvTFd+zla9FT+IRoXYeVP
kYZ49shuOALtd92qitgYSHIvmKRo9OB3NF1mvFO81XGq8MgYSEfuPUwY/UrbcftNxgfKBmm/apiA
TVznkW8kESMpwKjMW4mN4s0m7Nj/jRC9MYqiNW5oYly8nbjrEtToWILRjzYgWslIvbUfHxwojp+1
5wECI9XLRDC7MWnGans7yTPsjGnfi0PL4tz88eNFqgjNtjQIUi5fWluHK4a4iyI+KgaV3J9Sx6w1
OBx8/PuDYsPltnGNz/lWEpek0RM/JkBC3lTofozs1M8+7K5yqJdv7yoKsuvpW9zzTJMfKUB/dXIh
1bDozFDFPAagILq1bYlxztp/Vu3WjBm76+RNYlQ40XjfPrT/agQp/RAqg3trrROWzDWwf+zygEcp
Aso0TXtoHd4VfAM/czYp0BJ9UyAhbVa/MLxU5wBdw4zKA9XbU62n3nKuOUxYZWMAbntRtlUW3J7f
JlK4vx4OWOTpNkpb6iI3TBM52RaczU6VEPh606bcvPngglbH8hb4Ra2hp30JIOTue9b+Fd/ya9x0
GFojLMhzQBDxwXEpecGomfIwmkzei5rb7cyB6a9bz2c5GaMvVPfx64uzEQnhOv4pYReJmw7mUzWb
/DmBdVRyD+2K7gy2NTWLU1hEQmIu5LeeHi8rCIV9lClEvpHcDml/Lu76Kr5ZMRhm3sE87D5NrU3G
ei4K8ur8dSKyRA6wJUyZT9K+dt+EfrbOHIT7qtwv7s9Bft/B3GCCRMoOOyQ6VqzRzvuTo73Mm/u4
FrxMEYraY3LDdeSDVj+9QRi1UH/VTcf6ZhglXkNIM9V/IFQVceXya4/ADWmdduL9B+dPckLUXt75
be9d/sdtfMRlGXLIwrVoY7oyNdHmvE0VAVBUZHSQWGeFAPP7VD17Nb0eY3IfhYBxS9mnOMFypB+S
gaa6LzqQ8snpZ6eK2r65ThFZ3mMrLDnwxO0dsyjdw7jeoP1mQlAmcp1cGaNNoPLfuQGhdMgBDJmB
Qmk1HFuJ9/rR1KbZTFq1hWJn0u1cFB+iBoKySSvQIj8WKI6+K4QLXCSDJvS3sXS1ZfUHjIrH0BCY
7arR925+NH1F6fzlJKSsPQgtMSbnz5kLw38t/RShryWn+6Q3V1l+klJ02lNo1MBftgIfnoz8wS2S
kBYg7jY8QIiqj4uok6B1vekNq3NaqCLE3enBHwstdcAZQhnjOCsC4YQptVcIz96YjmNW8xAdjF2w
ecMBFYIH5A6ZOlzsAK43q3CgIQSVCqQbHBdoNiSeN6dcETvGcbBdcn2sfdhRi3hcyKASEmIQe1yT
2Tm9IVbfLR5xGKKwU8XxZbSHw0P2cadO7ub4VeoJ+3h23SEleXBnZUaitmu/RaBqJRYZtUmg6MyC
juAUs3xAwQfGSBdOjWFEr4Wlgf14Bw9wm7SXEiHIBPQWq3rXhdI/QedQq6HG5Bq0gAOhXCnnXojS
aAYH/b7M9RAFi3TUIlJmg9LHAKSjxX8cdSgV6edavrZ94ldC0Jvs3e8AZuJEWwnAPSTRE9G/0ALW
MaUGtzHVvCfvkHJiR5XpKGOSjdde0CCKBHLjUyzh7UTwTH1b5CLpN2DWpU9ED5zHfEZ8r8lhrjTF
2hkzsNruEX9s1P8PpUcPyLD3Za++RBP8+g3GL//lfWFgxhYsotJpQ+z9Xb62MfybMM3b1A7/UeZq
1lFqjJUoWCi6/0tdBzjsdhgV5WPv4tA/dDrj97Ss74efj1JmlhOntiYUzk5eOQERS71HZ5WovTWF
It3MARxxRUdcM2xnCLFbZ63yvBIiwIDt+HIroUwOk5tHdoSBxEQGTDFTK9YwsjRtkdJe7wgjA2kV
i0kT7uK7xprChJ6V7VJEXTIoo1hPpQ4c8QXWUg0C/iZ1t+NhJKFfevnMnjLFsMGAu6c9EE2v66wI
jeMIcbiqOxDxPg0NwwjarsYiLoQoY9eNNw+PhxieY3elB0k0GLEZENPyW4btlsyEmebbdTd2JmNA
pZy28uxstJTbJR+XbowfqNl5YS2+Q9JYvnXD1huB/5HKat76wx9DrYU5XpFQQwuICOAas580+KM0
guYV04E5PQHhv+kUdLK0sV/0rkmERQNFeq6M/zZIme+Cdb0AjJgO+TKxt/4tVNDhSbXNStqaP2g1
A2HjvN8h+6evE6sq7VQZ2KZuRSGba3lpKfToMdigGZfRbLBmhicgmr+qFYTMtx0ipQb1vnLZ4tDG
Ka7LygRPFhEg9+q91YueX55WO+sL8jaIuEQ7+iwtP4425+97mafMzqOyQ15lgCiTIvrJ/wqBDv/d
+UMHtkhhKvP/EAdQilkPY0HPW0kxz0F8yINI5ap1LPah6eyi7JSVvb6lSNs4pPzxFmGpqIV20OdF
9aXr7rS6bmWMq3tVQC/Pe8t3PRBQDN4WHOL2SDqTQ9qkzRkbsu2PW5FEJj9nhKgGWIvQsqK6Nmij
ztYR88og2gdWDzGu5UP51aLXVkEtmoNQ5ENXJ+m32I1A9Hx+6FDA6XFHvDE0s++kdKCG6Db7IdlJ
uDkwBgMih4Mpf6Be0zO3O1nkCms2Mu66dtWU8jx/TkivPWbgQjgNlrxL0cA8sEVsRYDeIE8okjRJ
l/QqBQskuULear/z88BdOBY48lsIl+N2Xbsc9nuuEfmkRzRchLvnZxqIFwqqTdV+jasQy/f54vtI
rzbjzy+XCTythvnWXYIAptDN2R2eyp9X4bW4JFZWXYgqKlHWad3elF/Quu93igsnAifzf0gscdfl
pWobfh1BPREJSUSYSYvAMz/qJHhZIYoehaZ4BTrGHNnSbYPKUEAGin+OK+jK8hixGf2G57nzpSV2
rr/E2rjdx6+TdDJf6TNFV5f19MN0LjLtHzAavUgruxNMcn1bbMU5fvdtaio9lfU4Owm+Cg+RnG6o
zOyVRyYD9kv93NWT+DG1w7up15PzPZOxf9FEsS9T6f8biyF4OYMzRb51qAB5qhbp9mCNxcw8TQIn
QE6w9Q6dSQzHwMgNQR+iH/54j5hQ5T+XCBnB7FhnArLOvhqNE1V30kr/1zPyeC0cWIP0Ijbr2JSf
ymDnn/cK/iJq0b+o+67Oz365jGBMv6EKHCLk/Q2ryKEthiK5FMho9GYqddMILbb/Xc9tx4U2gOXQ
tYtDBOImC6efmJawLTTb6pNyPA6kEFUjfncJHtMw6CCXrcv2a3OrzywYuioS7Q46PUtIlmg6PiYi
aKJ0d4M/AyF3dASQbFNtDCEz8yzJoqRRW02Zg8bZHlZmHqzETDEkwTMChn/NeP/W0m0hS3oTTfsF
CTpeJGuPe00oS+lvkE5Gf5ruSwvxHyW/RJU0MN234/dXaLmZYWhJMg/ihAxXGiMz7io46OzcbY/1
/Vq1lh0l1oQU7JWiIus+JyiwKEXyDXvmnzzZDzrUDdKTcgJHRyVAGN6CU7ZfjGtjJPrHdDguNdUb
DrB65HGNYDtnwQt0G1zZpRbPVg6z5p/K6bIaX+ETG0ipjLySaYvzT0qjVZJPcCPGx/cl/taNMwEx
tr+59cwe0O4ObXZO5K+w2vod2BlPqYcC6QOHmi+qSeS0oMRKR4ZBm4iVgjEk23uNSdRSfYpKSOdh
2d+ebg4EoT4ybOyFE8UoSdwzztsEtZ5LB7UKMUKWoY3PsUuapcx7vK2kbFqWVay0kHj9QTtty9pZ
bAKOjH5c7PqP/jjNFGYbp4OlHcjZzueSRTxCP0QfUMbLJlSQ/eSqwEZrteBrQQ9iBhXd5nJj+ryo
2cbWDxVmL7TH+oC8PAlUFzaMzwqXVPYuEzKdN9/mFl1M+dhxxYi7AXjLWNXg8ZxLCCX51XIH0vDv
YKwtKcIMV6TQlSA/+Iumh3nDsOyWpW7z0VS9WcxCebaz1ib2bSUINkMhtfpioK+Um8gzowAZprAt
1I8ObvcM7Fq+3yfFBaRW1fb9Z/R3ntfE0AhsfiuSPuU+/Lmu8NJdbo9wqSfCsOMSkW35Ipz/BHu+
chxJPfRqVMR2ThRoflkOBfuMJuRLkIqggwG4dsDXnBvuNRszrSkNLIBdqm04H0JrRcja4CPBogwm
4XN1MA0YAe875qlx0vtIPnycQFz5hzlyoTbskM4f0cT+bmU+yjnRGsFSjOgBxGJwvU6mpZteJa3+
QjVb51MVSPPfFSt894Q6TUHfGbTlWJpctaTvDbLgacqogEegHgAhYcgt45mzceDqhCH9rzgCUTAR
V3TSywz7E9Y5+NjF9u3WDHcNNlHz09WAFQMgkPqKrvuPB0r9U1DA4wKe2VqoDmqFEyD5KifDVMB7
0VQ4uQJDAGEW6H//lP5lKiqWuQpGgTqSwpjVx8ZZtpWeAFd+8+pZu2IjR9BjXPz564UZ69LY+6++
4Zxob+p76NlQ+8ZtrrG6JAdpCizztEOO7YkjDtNyAqZDoEGuTDUJVJ6N8s5ECEN4n602RR1uswXa
yflRnaK/DcLUCmjFXw2QdL5ErwokzHlhlaJ8gZWGI1iQwVvro0vICub1t5j2GB28rpb0vzFr9uQ1
B7LZk4nXkm5ogY1pemIa6dygK9Ly9nDYmVKwcaAt+2bj2A7gI5LjlBVpYr7Rh1xG2J2pZ6fBa0pY
xYbe2M8BN1SUojhJwIUPn92uLk1M2FqVGvhPOBAe8HganBelnBJpnWa1WMyI7uSaRlhCditMcDm2
2+kaVxIJ7/3Fx0jwfDIhGR9KTwXFAyR0IIEl2z4OUueZX4gqJ9pECUSoe+CFD3gkiB5z9ThvNlXR
Pnj2O+8VXTd/vR9Odx9KmwgIa7hdY9CNv9Kwr4Kwv9gVcHZXTOPXu1q9DR2eoZ7ormEJ5wsriZ/r
WuDrtv0f84KKssgtvY5fWNy8Hd0QCYhxQj6ElM69TYZC9m76Cq47cdXWzafNQf+qiFGuBZxwZBOV
wShRkifTKlK593O7sY+IzW09nMA9ZAQz+aFFShveT00BnEAofI6BtC0HY61NY1RHI2OhJqJcAN28
5VeoU2i/r/knPSAhV5w7gUJIV+Hql3vCqPcofKKXUfo1jDqVlRmjwBqdwG26Salj9dZ09w/FSoa9
LJ3PC3pbbBkapoFogxCCBd4gO0STyxnqkDCbPpLLpKXDkEged/xkjRwfrwfHUwF2aAn8kaLEIERB
bI2VoBf2K6GmQjWqonIlVj2Zb1FJeIOQ3xJm4A9smbKBW2Txg51SDVV+1B58DgiXXXhQV4dM7CPY
RIofwat3JQYVNNy2iRXD2xUVB2sT3EsIo2EB+rrCxtIPI+tKBxczsBP7bDpXpMUd4hkZwstb9nyN
JF+PX3Vs3IeBvptdkY0ZOBKcGxnC6QbY+cxdn5c7avkhvw69btij4oF+2Jh6PcQDQe6m7X0PEsH6
xjrjJQ+SZPbSPmPdNvfAs/ZHm5RaLxFobdJupLLIFOkRgMgBKwiThJj7bV+HFtl5c71vxv4+yyrR
jTRdUNrpY8yds+LhQQ7+8UhqO60hYnjFdLsHvbvTatwc3n3f34trH0T+WSt6/1cnIqxGuCcwj6WY
9XhSWRnUe5uCZY2zJEcjMTt1X60/HDAcmd3eeRGGCUcAwsjrYdvQxm+yxIq8aRXsVbaNhzuBjY/B
uC3FB2zVZMgdpbOWD725pDWU7FrKA/tpwLeDR7ZAQl7+jYzEd3aujjqk03QMWu5DK4PE80X37kKj
60fQMWOmC8MS3IU9oLUPgB/FIwhcRmtMbVsyZ0QN6+ldeG7rczJIhcZQvRSIMD2h4AAoeG6p4LjR
gKr2tsvkjJvLN1ffusleWmZGHDhlXqLdw/oxfBVUbqaYZim9/8NknClR1lMCCTeFTCr21NrmxVRO
NmpRvOZ534OKueDt57soWh5Cjn2Iz6L7j1V1qIN5q+RcaIqGvQGcAfpkBym+ckG7EPwdxrhHwx/g
PLIr6XTxita8MyiPyehOlLo1UmgBPAKqHqN/2P8lMw7KrW7j7YMsyslvf3akVYrppBmUy2SdhDPN
DmN0YJ2vlxDL0C03gCpeV8br8aa9r1yvpPQtD/2bBRBdxBxhoPywcsrkhCDjSltHRHr1HNE5SibI
sbzU1aFaWi2qEvrUvxnrg3RfU+Ew4JjS159jlJjhfEaYm7BQ+Y2Z+poReLYl/7uVUnw4j4ouvA9J
PFYmxxCcq0hqKdrKeaJBEaiBpvxJFPWs3Bkyc77qrFramCpmVbZJD3lkH4awVUg59ANKo000elGB
ANtwjbblm7IkabixA0qh6U+UTfXG8WSIipA+ynM0yc87s/DOgdCjKosN92cIpqWftrWibl3RU2UY
zfe4o0Lk/1e2neppc9X9kpmMg/1lrESFZUcQvVm48SngzTsVJWKteTCEepxTMSY6s69h4ORsHdGY
N0NUfXuKTDNYWKvuIhFtKffiMmxdgyMxRO//fK8NHsIk6voBVAtjCeVlMBWW2m5M/tIyBdPExIDI
/ZTs6hu3gxjHw9egaF7IkcDVXDMTILlBOGJinu11xoLA0ESz7NsAfpVUzcvNLtr2MQ+XQSFDFXsU
fuWahSXuEL1xyEEbCbljohIP6f+qPOOWLT555yPvmDJ1BATuc99/Aim2Ow5GBWnmU+Dyq459vOwU
dB1dCYRZcCphHFN0A85QwSjEEJoEmUeJI4IUp8chxTWP+0skxL4ZaNLQsNsbiTElnP5IPyyiSpy8
iDwDOU1qhxldedIEMYkdYGZmzeqTFjv2DLjhz7qZ7vrHGJHhHqVsz2BeD1JXvQzh3ym1seXYK06M
blnG2mYDt9donohFIoEoDA1K9+NT6BaLZdLNI9vn9knn+yHc69O5f49OPmYxln3bbybIf/YvXBUx
t229Pth0jXkjfHaayiacTP7bNXMO/G7rS36qRFcnnB9z0ARFzscyn+5wjpM4H8EgfnwSqqdq8wCq
dLDUm0kRQM/Nnz9YzNSzqtV8YtiD/kGDQVCELeejBmcrLTze0B2rnbg3Cx3l6bjQFLHDgMR2slP+
j/3uMjT+hRbime6IU2M4N8ui+m1vGM5hV5dXAOEAZxv6PfeBM0PMNAE/u1Lv3qZ9fr/l3G7LGXLz
VlDVTGbpmbykYaC271n1Zb0n1WbMIddJj7gaxZJRF2EIw61FvL/1YdFmyvZBamwHVRzsGHUHsgPV
/u7ehXQN3DONhf5tCT4zAbM6FUyAdJwQdlyC7WKBFDQA9ch8veR7XbtCOnZbhVDnGNmGHf3zFBLP
evAVuyLKbRmYjO6QZ403Bjoj/SdO0V2Fra95Go2VOg726/9ruNrqQpfIRISztc2P9xoGLUU4Y4m7
ShyonvVemq5p/SUwiNPt9hGpwgVSpNtqYhHcFCN0qNPXpA6A3nXgwDeMRd6Yj9r4DxiaJqVtenzG
yeb1tuADqAf0V7vHv6ftZ+EdJCnKK2ySDC+4moktuscjz1Yqa8pF0qJ8s8xwcgNZRYknczExUdw7
LGSGnQU8V5mvxpsfZ0ZMSufV67ox2M/9ZbIv0i4jYN08X3ck6lvWJA9gFCxk2K78Kdd9kZMc3VMw
PkkwWzSMIuJj/RbCAHXVH2HEPa/hYWh+FlpcNVtAnTCogZaIDvOsAzAt4MMEuTyABRcyl/rhoj0D
C5c69iCbubNrPt6Unm/gpFpXc/CKzG7/slEXQMaV7pawUdBYx/RTFhP7xmiGPfo7IjHgt6N/Fv5u
+gmkJI8WZSJM84XMYhdpRBOjTwjXp6NffCrXg30iNSVdzFL9i7Y4E8SGpFwk2D+6l0pWEtkaNfCr
Dnyx6juuyXx8PwlfrAKJdHGUSeNNvLwqu8LIDq0thS8lhgdkU1iEAxFz0ZmuCoWBp+I+whFe5HhA
/jEI2vkHpADbPtYv4MWLtdM9HeiWUzhIUoPQxMlIDcf8vGARJ4yvsa3Pjjju8cBUm36ZWqsWXdgp
kO9tDxS2nDAMVQ4L0LOUGch7MS6xJS0s7916UlJBbXOJUKpZf5WGSiLjRxKBrd/h59qv7/JHGjp4
Z0XDygFZ0LRXiXGS9rlS57NA+eQbPKIRFdPKdwpjatfqPeMwc/nct+8cYUVlkvHGuKRSOVh6heAA
rD6Jeat0GVQ+9Ubyp641Sz958NBDWayer5GQxlj/howomi6u3y4tyF8KaJRDlfTbLXvVuO7Uxdv1
j8jZpppvmfyP7e73nyit7Ow5nX6/Ly28dMjp8wvGuKlFj0S8n7RFY+NuItsMUyTgW4T3eLiXzyTx
yUOc0mu9D3uSFU5dGnbHcnYK+68nGJ/2zwxNtK/UjzDGH9RqZbbEf20uJg+6Kl1G5YBIqCxTu7PB
hJfmIXWlzkCsDjjL0mkqBi8LMS8G2qsXy3widIE9oZ+2u995ufdPU7i5s50M4xZEwoxGBYYIxltS
MZFIt8QZy/2r102hWLbYLkjkLRwgyl6X1Gr2xw+3l8FbwBU15I7Jic6vNXCCL6vFiMtQjyuIaEWv
JIK2fZw6iZbMn7CjcFxezcEk8wjTAq86aJhRjvF9nNyextDV89Sa++5cgysfNcxXs5xbGwpdxhcK
AyO14TYc8EDvpSULu0l0XBsCF6m9G+X03Qum2ndV5viWk43tl4rP5q/RwaAk3DtUqukDVx3uHgf7
5gL9xx/japXiuVXIMI7IjCFaRD4atWwlc9tbUJjwhZLU8HhoHtuMjx3ErAtBjPP1HxT2xwUA5wdP
uxR+9HFkiH13y2yRrXmhANVK4Mk7y6gh0wLSfg5ais3oWYyECmLcYMHHBGF8F2lwlb0yjdhuWMRz
KLX62XuKaS834l4TJamDiLvZ8dfq/PM38CM32v/Xw9BT0j8KKwirDlJBNedY8dQDubMaK/nzecFj
R3j0KSx/gfYVUlLecdjN9I83uW/77+jr2LBgd8FLYinEu2EjZR/o0Cbq4H70CLjDDs/9DR0ojK7W
73MlCMeLrq+QaS2/J72qYoffgHakvBClK/ShAYeD+H1VoNDodZkyWtxKnmfEGTRJ6aL3ZkcH4YZM
9RGBQPkNqKtjtm5bGFyvKdqMK8HVdiwmfh8yZ6m73OfVBm/hW2RGFjLFrRp5DIwlNGyou86cD+Mw
QidmHM0ZzUcwKPRoo/7/i7f2gxytEIfFCe+I2UfIWjaGq018gNPBhg+0WI86lBhoI/yc7yPlN0hP
V5Sbvj4LY3tHecDnKG8Cvfg3Q56aBshKmf+XEMRbBeGBZ5UtC6gqNrKJl3ceCO/TpEAqeQn1dZPY
YKyX3FHvP2/OPhM/PYISSsnA5g6tdhuRfoVqAZAj/hb3k8wmbq1eYUCT8nNBtY7dKrBJNkeGbx4P
M+lzllBhsrd3Q94hGNOhOwWFMN1T2lwYRRkhOTyBysM1bSL/mOpctIM/TC1qOW+FVxmR/i9ghOjd
n0TmcYjRxtWPG1OglliQ5DnmqIlxXQUAIveXyxercdS6QL2qUBzkTtiOXYzgC47C4S7OmtGC25Gt
NxaRccLT4E5Zn58e6t2lhCeiFp5lOYyWCLwCHGoYDkFYcWokv2Qg9XO5fkYLLaYi1uyQvb+lZYny
Pmifaz44/JESwGnc9aXqMgtpIAazdP9HWuFSiv62S1CEkHMDtZT/bNmrbMSfZTHxt3esxskHMR18
Um2h8HCOobm52cBhgr5dJIX/phmr9nsd07VxK64MBGYlcDs6oPw/LIU499kz+E3gyDrpCM2pFOO3
JFapGelPxxLdPdI3HICPLZ+AWANBLiarMLSQIUQjRZgrmNmYus1RygksusKPIJJGWStcScWX643U
wJdwXOBTS7c/zNgzfn8nuSho8NBpQn1L8/b7fBAVRAFqu31lVy9TXW1gshbl69V56KR3kTdYFMlB
pdhKqeLTvTJiqzLKmtWP4u3s462Z0pSXGA9HRawxoX0PQZoqREGjg/8OM8r93wWd2TLtFbjwWYEJ
fmf5jBBW+UOGtZ8VdaWDWbDd54SspmF5EJhObL2fTLen97fmosaM9r+mptEip0aVhyNEfffCCcj5
Q3mWP+yWJir3AYQAlykgYmAsBjxemQguZ0CveH7c/N3sd+oFgwQ2LteEs8Jb9B1ZAYB5q+MgXlV5
0BIG2QTFcZ5xRDaMjwqXeUR7rOqQEl/s9EQmUrSjgzTsIpopcglVnjcK+tfoWcMxAa8au+YFC6tz
v89OFkvd03pYP4q+JVi4x4zOTTZtdg4Y3b9xrUgjkTQRbaBRCQhHCMHTBZ66eRGwQzQKhytndVgd
q7cMQ4ZQKWnB4dZrSqTcXDY91TvVoc8nQgd5+MKnXFLMU4EDTAJNjUAnFILDye3+lMvn+1PBCB78
Jgs5RqUh25m1dWteo6fpYj4YO5LSMdnrsMZvBi57GbhWh5RWCGg6/iuhcWJg3YSiBkTaYm5SVJun
nxyMPdU8YSoYPIF717N3GuGzvePU8NHLTrpP8+JPapZmYLs0nctYRdcryKQpMLZ8Um9dpTHOyRKl
n0DqtVp0yfN6T6GOaRb+mADdtmWq8/VQKnMlDDkI+dtcce+kA0JPRGg69PTr2KzJWXSp7utf8oop
T5NqOUkDjjQVINv6XrRRdue2HglTCnNWTyDwCsDfqpDvLYIqx5WY/Pjjdi/0CQaYHCu+N0wM9rb0
Cz2ntJ5gtFqeArotUbd0wHm8UB5e57B0mnOk8d0FxjjoR0CgTlC19/gcp6VJdIxOSucQ7pAxh3VO
r3mSJFTfTnfRd0pE2kBziT3THN3yj0vPUlMZPFzECGu1ejCBR/0bAq7lAHI39b0+8XPsplU73xMV
MsOdsuwv918ZFAUBPQCt7z8FghbkUUifFqcrottSOZyu3o9I/5rJkczUvpiZS5/XyZGcbCYbCtGl
EIyf1xB7MgJxYB6c3sewXK5wKzCCAFEDYbzEXRg/9sSxUY5JXi5HgxyHSp+uoSUIwW+A240af3mx
pjNSHlSQMOz66TPqNWKIh0fy6lvOU0iXcdpmfaMZrUk0w7lwrCIhDJnVAqfKlXORxdptiDA5XbeP
ydTZC9NVJswnWo2M90fKrcQCyl3YBRElEzlIMYe5T3/2yRkq+mAbXYCOnDXpunFEj3Pskh71KiFE
tbx3sbHF07hkvssyRru3yy4Yg8k7Je7LFs+c8w1gUDVCtlbZc/EcUanA7xcw/VDZsJVYu0uN7JA5
2ye0iCBSeReKe695N+HGGe2B5fE31Vvr76yxmGNIay5SmbqHRrEtAJyJDDo1QpgK8So7ot3lSNSk
6pGsYsxd4mTilPYT7sN6tCpurFirKDeYJG/eIDH/allfXKlgWvJEC9WUyWqeuFyTr4E/NwXmP2Gm
0mec6Dn1p3OVRe5CKx18RQbtfTWFqK0x5ZupFU9k6appcqT3PKANjJJCfR8noryPZLRtnVfd3Ohl
qphqUQzHSQ8gLjk1nkwQCg5pZP5FH/kf4SqW/3b3wTYib7FoGs/GB4LlZjzQrkrla7bHppUdenUv
0NAIR5qSddty3MC1dtFYbRPHUVZ4RjJU4H/uFoV07Zy9VeI/6bPEOKF51DqDRByHTY41mg18FZpc
ScJauJUlHbLJ8HKhHaLhjedGo62lnVSCA+eTdOvD9jTJUQcpAoSpzy89KmMA967JryvGbES6G8+L
c6dXf7RbnzB2QImYQvV3VdwYOmb9lWLKRl+N8Ud/Cmkc94kTiHZIkNDs8Rddlcc6XZ/A2RgbSIIj
Z3vovR+HklcfiMk6Z2c7S1zfW2zxHbQPoWszIHN2oKZmzeYcLGEUXtPO/w8HG0Hnynvpnw87/VVb
3OWQ7yM9ncywc28D3INtfUX/P46Ut2MYkZzC+A0LmzAWR/MjGrz+ZFXUAcYsR+gUWkFPvcn7cJj6
XMfY2ivSiL83i+ki6yio45hY/AlUSyOnZVRuUNuykZWi2N/1/OgaVYZIcFc/evrOrdenDzsmdfHM
dmqNNQo2OpocFStP+lZSM7UMlAg5B56CPcUcDQM9GCzeXNgyw2vW7eknReS8GGvc4RZdDucMvFn7
RDVmKWbJv/PdEsZv/wlmxn1M32dyU5ppy4B6f6XugiWwoFjbxtJsaAHDZ07cd8xDWLlLB/v8kIsr
0cR1tPDDx/9goKM47ORjkw5ka6lwvQv32rt8HA7SIjiegakKgrTqDH65jk0gF4MyG0M6ZnNRCKAB
pxBsd0A1DPQ08DRho1R1/NO3lCpKSNoeTIVXf/9vJGlMOMC6hBR77SmLJUjzSch7gK0f3m9vtMOi
VsLkt7c4RtfR+IUpNhMIoFFh/vK6Yi5UgQAs42c2r37BWuhyXKhy4GV3kYMcb7bGEDSa+gaWoXE8
GLRpjMcnjT6AUAZcY9LZQZVqN2P2fJIcsmYPynorcpfv5w6YH4OCTRfbhRXYCUYyZhQwzw+eVklG
Q4IdOZYkzuXiC4hj2+kTmCRw8cLpd0FE8HKkGpweAfSP+M5+DhIv5XnFCehRuf3QvvQcZO5Nn1zq
plrAoi/d90FBTLLhxfEcs48W6+jZMNdkw1W1o+PcKVS/E0E6iTr67jb+YCGu1g644HdEWkVRO4XC
ibfNNH03XyTrBiwHH/bNAqAOun9eveTvaP9CspOkKXQMIub6B6rbllWz3VVicut+qoYybjH5dZ4N
dUXUwh95wLS5I8RQgBI389ZlApqyUaDTFpDuE2vO3i5FKtEJ0ioiQk4QfDl/7xvXH2SQzPgnKtYv
pklu7oLqR3G0a2a+osVFGCzNgiKFfJVsgI2T6CPZs7avpTmMmCUcAJThvqrq5joRiwZTY5gBZluW
c5kfJrTyQGVJ0YeueQfUgdTZXgKLxeKTrG6L8m00U3c9+Yp7LmN6FEqCPawaclRHF2CKG5NLG6Gg
DDBIEIfyWrKv61wLCDA5cXqCE6b9/p2LeXGJ2RFn7ubnSbPd9gA7wRqfbJ1juF+1eY9SKN+wqxOz
dLsiboxtYNDucSSE3qug7iPo3AZMSZ2mnVnKlvs7sHrIoPuaNT2QJ9NzdEke1c1DXdCpgtU980Fj
bm3XS4ShFlhaXt3AvNyCH6ffHNanUOBuo5Iba1YJuLc5mOn6OcoJRTiLmeAT2d5nQ5BQNPcsRJii
4jW1voHbX8qApNWeE6bIYxgxK6a06THMBJJsLpXHFSIqMV9Ho+onw7Ca+QlP72iv9/e4Dsck0lSM
QWcf9SX6GB7XxvPxV5fn0zqul2PTw8Qx6qeV5zfPC4N3ZD86QT2JtjNjbfmb7jQW2IIF7Y3TYCm3
sHSlQKcsocL8T6juTYfDpNzCEfWRtvuT5r3tTnP/kUNcDiB7drSNfLuRpiEj71lDwqdsl/6WSfAH
BeOZ/cMezh/WomXrD0dQ3Lv0bXCwSHh6kBng4TPBZ+J4FWO/6d4A22b/9QQfdONmSOamWRbKAnrE
Xuo+o33xb3RXh0lTWUOKfYLWHV79HDhh/lIPaHIDcNLQHcq9wZkunC4s5Nl8kn/pE5asmIfR3SGY
Ih6JcRk0mC0NlGR+uu62VYx757zgw2PP3Ic2DYVyqy6Q6dJoLVPDCltKRNN3lOz58VdxtkT1LXkQ
k4M0P5XG6ybGl1g2s7GvJzYcDOLAa1H48WbMBWxNnNhO8p6D5NNwNB3cIQlQZmlTjyE8Orh9oU4p
J7ypdUkZnsg107KAxTJTQSqu/lEapaTfTTKL71bsw1YzoxBX5lBvqoc/EXiRnPxWCCfXCprFLFD1
bJ2Kaatnwi/WIgqa2mn4KaUWtXDE8DJuGUf+TdQxnZCKG1lxT1AgsKhbrPNxtqJZwErNerv7nr3Y
ivI90HlHOeik26V3OxBLATNTuzlcRkACRZNu+DAdRKF+wR3gpsoeF2/SOFx61xs7sUobyZUJ8noX
fHgD5+We8kidp5Xvy5Bxw0cGjU+I0cHvj6WR1wSY2UXALpW0l0eeyyxuyKpbS7VKltezVkWf8mBu
aznZ/A5Y6znqzXxm8CiLo0/4+HiJrAv4zF3oQ5kEf0Rl+/EeWsz4hwmqFn4JDldiJAQbJ1p9Jwo/
Ax4PdA9JHKhcKn/S8dyOtWjl+hkXbKadOEPACYDQKsg853zGI2SreJRoSbVwPrv9u4/PxXzMXKuh
v0GYwIwy1BlTK6r/naF39r/XdtQoW3DsN1Q5GSx4P5m2ALFr7zfKOBh55UvQorHDrpc+QsU+eIym
XIsz09fA3LG6a3x27UsKyEYO12+PM4fOd+mUaiNOzvHR7Et63kE/YhsoReJ9+pJGyF6vCczKt+1X
Uge4S2AGlUxUug2dDJ7rqWCKITgOii6WS2kc6uFeCcP05Kx7C7RJu6JI6vk3/auSUfLR/VKNwcj7
ysNrns+bMe1jfwU2/HTQeo2PYJZ8XJpaIcA1xzBNkWU9aXB8XgQxbIFcNa2LGZxNngAq81iDwEqx
tUWhy4WLybgMvRcOjivYI4q2Ws474ho+019JX+BXTvQbGhclwtrRLFbuJNAoQJr0sqBTpOGyaC0t
tDpWnO6l0hFB3N3x5uCvlZzG7PCMkLioJykothNm+xIIEmXof9QoGs5LUP4Piirss7wp0rbQmMCs
V3F+L3js2EmWwEdFsJ2IZk3ts5l8kmY4EKozR/cooTu52flE8MiAui/pczQ6wTIw44MkAq7Yw9l9
v/yxPmKKrK+oDseMgNoYwKWQNXgdnXAIlxR/lUJdwKj0ocYAaS2a59VIDhevHKIP42LQq45kdkmZ
Q2I4ZeRR0tPu0bSLYI1a/vFN5VjfFmkaDIMcu8s3+hcpONknrP1nZWbDMihi3wrI69b/VUpgaC9P
uypvDonf4O7QCd54fORmCUQjzeTg5UivyS7l33j0x2ftoOjvEZxa4nKkq3Njug9piWY5gGwEaVPF
OxZQvvxu6Ep0aN8MrPQp49NWwjhsYfwB3TzrqsHpmKCWXWuvnCpWEDbsJr0Mkz/ZUpyEMybGG8nt
zsxcSbpj+qxQPz3aWPESVOjhxMr6/V7RCngjfvApHmpuh0egF/l4sMpWjrZqYqgY8/WDIiDu+wsi
zJVlmMqMAryc1EPp+Sjjb9Td1zBOnXJPOrAFUhEo86xdBks6Hb9Gf1H0sku6QXDdgKwFS98DrWrm
Y0jALPnYQUDNW1ftuoCls+rkENPITEjxRo9Ghriej+yFxmekyhr4u/D4dWYHL3zCJefcJeHr8uFR
WXdqlz4i6ypu3S6Ooqh+E1w//fW11Emram4/wy4dvzeGgxmSDCF/j7BJtTmEkHbXH6qtILwbmxVq
10BZ77gE0E2uzrt9J7LT6ZGO16zGnq1TYCKZoEgaaKRZhgb1lSnkpYXrZn71fZv9LaVBRXyXSkuJ
A4vzrnP3klBzwPjLPIKdZJ0hVzjwPGgjkhcVMGDo0XG07hcZ10Jnhs5biJtu/AKX7mNCK4BHe1Wu
6jrsJfRC2Dbria35KFGy2tXOxZhrwi02Bz6NkcWD6hxc2UoTi70nFMo48Bvfv4ujSaG5v3iXKH3e
eIFjQj9rnpu+SeaaBW58CCCG1+EGTnnlZ1iW0HUSUey/4a4+eZDeowgMN+u6TMhosF94rebYI3I7
4uenbqOE7/8feTsBWJOB+9zs/R9BEK8ScdueM9P1tDWhsOkkdMf9SzZaEmydgdfw5zoo9nc4qkt7
I36zXuOu5lB2eBRavNKr88CvwatbKPu3407jtW6px0sDPYYfzVrr9tq4DDv2LM3YbI6tax1uTKo5
gmUApsjbB4jSmCSgzNL9UR6a4LPis0IrcgO+Bb5KxYbqOD+DY3QxjHN8Y3itWwwSAz4elFuIdR1F
iLiaqwbFQOWLaymQ1WmRWmwhkP5VN6sj22LJZNLJLUKu68BblB8LiRJt5YD/mQiqCkpzztSvHCJo
QEzeurMvi3v7EUUTiXwU8uOdDEhCOhpCO2tB7i3mIW/wvufuHo3t6n5kr0zhHXiiHeisFBhASeW8
hzld6t8MpibscIYUoEtblQTIbBx2NPX7E6rqUk3pRBTBd2mz8I1azim+/1wtLcUKxeq773YHTbIN
p3IPcIJDWvF8NzuKHEWKckqKeMrGPBqie2Z4PJQIINqwxu25MPSP1FlgFlC9CNA9Ebn3oZu5PYaF
oHBEa/+5cEqSdyyLRpq5r0uBeEpQzy3XNjRk+fHsf4KpPbvXIRR6JqpVuKrrAH5Ic4vVhJ/CU7oB
2+xs/JGn38lPk/gBUMEZKhPxKmvkdjD52Vp7V/GnJTn+VBHHhH5HXFWY98FvrTf+VZsjSYvitKxD
Uv6Vvs7Hyh/yIiinENA0afOv3dodoKWOnzS3KRPvwyeYuQkHkPX/WFK16R7TH3chQCgIT0dribXN
vcn3nJiqvq4hpDyIwf8vQDPV19pHjxI1N2UHhiIScc9P6Sq+6yx7smQdOP/HJbDYAWVqNi0eUTkw
9qqxkRte/pHtBsg76AeFJ8huw9uCwyXvsc/Kw4K6xqm+hkRmVs8UjhvdhH2b+ZLBvSIcYTyDOj8v
RnMT11CIYo0avp37x4Ki79TM/FZhp2XdtRt5VQaQwkWUYhU0kM+zmz83mHB7mxqtr6quhg9WQSlf
6PLJ+OPCd+IPi1j3V8VPNVeUPbHD9Lcd05NKFS1qLaMfV7Oz98qoJcaqyefvn8+rNlwk9ninJCoB
YZ9qBCtXOvGphMMkKza2aJkI7ZaJRalpPoOEM7af6jjwOF6vqUMW5XRFcYl8ibaIOY68whvI0ZZB
LuE21hqEqPikkfFTAxl0ft2tT/poV4HwmzbqB9wJmHKdDaEeI4naUAVt7jLZ50M3isLHg+zMjmq/
IFxC7qCfj8NVxjHOrtGrU2Cn5iedntx8HVIHVnGNOu70MQBtFLCpXO9TSIsazlqe31R4VjYfP60r
Jgr/b4gjbcgTbug7vy35JTYrdHWhrpsFIBwvsARaLKwhs75vipoipy+ekqx2JaZZKOEIyzSipPTf
xxy8wfTMaoKsAHtd15rNy46N2dMR3oOZGQ3k1Ip3v9AGDXq/M3/svvT+pvhRdzndPKw4a9lB8TF4
/fV6CtOiRZl6UGJ4/U1CU41jQ13mwCyK/X4YHLQiuQX6Gy0HLN77GduTo9qYCoxgunb/QUxrKbSc
BlN9fzaFvxkyR0gF8xJsCPFOjaUkNYUNOPGrzuNQJZ6pmOysoQ3hGi2rP8FpOUzbB/DSwUFHr0WS
x+wcWUTYKHQl5eYC5ocEyjuPwRIHvANcCpFoY0JrYL750m8bCBJtBlRVXLi3ahHdJI672e5qQPEI
LTWKHWK05zhyTm0wUKjDU9klvv1JkVYKE9XJkNnw//XNBXqQnQW1ZDbP9nNw98PuVmf/CrkVUYbZ
k+ON+rwRuUwx/XHP1lz2Kvmkt2hjrAKuEs858dHzel8PS4n33PtU+QvqzImAEUbk/Ej0+uwSLByb
etYGaS97LB0/omb+J/JnDOPWuz7Lx3+E7asDSB3ecmwRjaSFFUz5UcbR9LD5UMNnxmFHKEER+ZaX
aB/458aX06aiJCerdBW4dNRWfldRIY7PvuoOHYBxILzdxNc6NmhZ7A80NFHaTlaAMz5G4y6HEr76
gZu+8WCw5+Od1BbpLBtdmO8RbIR7IHqavHhqniHXf5nJ/M5PqU2esE2zvaxcYr8wW70tSVUH6X/I
1nVTeCAXw8npYX37Edd6JDtYyMaoabY5Cm7eJdMifE1DY28gMuIN8vByAuhwyhD3PtBVBG1/+oR/
QoTJjvCW0733T72XRAGO6+QKu7L1zxvA6aVKI5pt5zGQ+Yn+IJPJ6ROKfl6vylJRZaRqjCxtT8nK
TyPUvaz94v5OoVMM948Gt4rmv0tj3Ji6/CvHX3vN/9Y93iO1XAblHLLtXwMueKmsnhPhwJKqpcnG
DvTnMqlmZGOV74OOEUhD2B98DlltX7dr7d8ksv5c4b+BKagtjEayZ94IDLrH/7u6PlcoZbAcbVRS
TScURZUh0um07eqLr9YpoeaOe/TLc3OlHiyPyv4wkxWTGJ02Ec7AW3fxWDC1EyxIBCAYC5Nw1CN1
cyhkK25qA4Myj8bxzCkboCuCcUP+ojIRoJztcKi+tXgBjP1ZQLkO/xoFZHlpy/dDfjYBHzxatAqt
qsY5dmEkl63jgj1CuDh29oqULJxkmM7fzT7wg3lPF7dSpYcyzwaHk0j8whX+W6l51Mh0v/EVNDv1
FCDD9CmQZ0yhhZL+6zbbKrsmKhaO0dNnZKJy1Ywf4i6bLc1HfBziFlf3G1Qe+ospSeu0Fb1b9vhZ
ZxjtNGtF+9R23v8faD8OgJcDaKqvlQ0x5PjJmjKIzE4o2Ks5NW1damAlaLV+KdoIu1dAXRmgx/rM
qEr6/r5hZLz1UMP1zEQ0k2zFNuKiacI9EfIRdNMRNClAjSB9mcjOe1ZGAC0lbzSIRIaf1Z9+zNIm
j4P+wPT5DGz96kTVDoSPcNhrei17WY9KKILUBD9+dlpLSlzVVtgpRJ5tQRNOAKZW9x6SJ8BbLrzi
4CziRXzTvGhC7Sq0/np9uxC67y3yro5/1IE5nuMLTmf8fQ1L5/JSks4O7MUZx1QmJgyDNa4exXbN
x/Rg3iLnQA5w8BmocH++ZiBRngx9fT2cJKUyyfa2sl6yKsfUFuvL3Gzp7Hlmo9OKMkhX44p6XroM
Z5k9zZMBncHzbDURRRtDO22QW0Tb+kTM4Sir2tc5FT8gMJ0T/xPdQzdKFFxY5GoAcFDSsvCf/CQp
BtsPdJ9XrOH4w64aLbOqSG9jp4Bn3APcbNFhalzMJ7jUl2jSmbV/ITtdBdQFd4Zrbu22TvFx9S6I
bNzVieVR+DmnG4A3+GzeD7aXwGijCEa/cMxK17vRCAp56e+u/yRQVAP0lea44lmCv6ACDPy9o8m3
IL2n9yFxTlUK4vni3mRoPwHwyeS8WiKPcwrD0sja3xtTNEZao/EKyZAdrwco25nmACE3P65isyWS
ycqm9Va+KnGQx4tdNpbb4l0Xskst6B8lZiOyxKvjUQJBQz6jb2fpkfcNvSEg8ElnTgM+NzRj70BE
LERnFYYdR3fUEXnoXA1A8dH+e9Sp0JnKF37Gcm2vh40Gtl5fXuC3BhkXKD8QB1mORXE9cAAxPpv+
mtKi1uNbEVapnv/zOyrj2oPdQogBlVPvW+OlXqTcpACQ/jn64ASgrTrAaWGkxHDOvwjOJ9+jyeX6
BjUe4Z22AwT8dl8DnyEgVd5ueepIAoP72bKSFzlg9CGSJaBIVTNfpWvNJSslvWHUaBPXdq7Ebsex
2aTa1inbfyYc1fqZuwVlZgv6uMMp1UNxtR3ENRHo1COjU09ajQcr/2F6FLhvOF1oSDfLRNp9A4gx
e4jydFJFN34DicwClgXMUuEwYijzEQOppiKvTgibYYUcVsDq8HI0X8Me6cP0zWVyY3Wr26YcPMcS
CmwSPh+ghOdMh3vLw6s9DXpNxh2QYhraKQWZxYcP4qsqatKB70RqClZHYQgacoFqG/GeK75PV6LO
Q74k1z8FUmj8SWHi0F7DTnZDrVIY1BQ4kNYxfwxqdSRDk+8HkGfNE8I77Dvyg5juCKFeucJtWrlH
aGYpuTslfZ5lwh3IJUU33Yy3as2263x/x68GxZ5w05ot/4H3e58FQNZPisaezS8MspeAwI8CvMFc
u3Z+r/tceP2XkCWzVaHS19cn9mjSTZvF/RmL4vHMoMkKGT9gm8voY29fMBCxMT0Cz9RzfLc3izzV
SXk73l+sBU6RfSkE1BprWhKPsb9oowg/b+Iza18zZ18lMJ0+IGgEtbSSLJGB2ybteovBsxiggH+t
xBQu2cRtQVdl6jzoYwVwCS8mNNYJDbmgtY4KNkWpty3M/uX0ztwRQZm1ARcAV6mgY3267dUn0H5D
C7MWpiY64Lao8XT8OKQrSmBLcXLca0Osco7uBq830FVvYR7MOg48kkphaFZvhKvZSpdPuXQ/u7Fi
SRd+66MBlVFf09waaMETCAXRb8mFM4g9lpUc6efsw9+IEBLllIvyWnqse002ddOJq/Ge3B1IwYBW
yFFaJBlzmFhxFf7TmVT4R5kPSfXteWVLLNzF3aV8I/Dfi+0Mz/QTG1kDyejyvyJQVkrKYob+FD5s
3Qo+u+KxwH2aKrJ+jPDw1hqG1W8EiwXwkvDaJAcZk2pQGp0wKpEUEK3oGEGo/WuagPKdmhJE88ry
PUmEzMgfKheKpph6gdxjWaWK1z1VwCXTKtNychFjHqiyCuyAb8cWl111/B8IlPdTXQUYsmir8FdF
O8FbzOyr49Q8C/pKZY/oeDQqbS9Q9llqUKARYrYCpEBIM3D1zkQ9T98ilLMzFpadUO7HU4vxqQDq
PmhNfLqbtSBdmi48QucsJ903JiXLO8plThxT3b2LpqAkHhDh/9LwviL7efVrZGIaZVHH9f1szVVF
3wbR2N6m2sPHrywJupIi6l8NFZ3Ftg/Z6CrUYulPIFUYYy7LRkEvQEmlmLVFR1O+bW/1/Qa/jiyl
2M0tm1VWt9Cazc1LwKdZGqh2ze/ETtilc9k/TWz4KayR/9epvVY9dddNYNJMu5Ytt746TPU42Kwy
b+A3I4PIPlC4stpwZQMIPSltuzNQoUr2t71BaXaX6BfINAQY95I2uW23uD7yqklXbrAliUkdMf+Y
jr/sQEzQ63ypNdnqhD77LAh8631vDcV2M+CEmUUVQwglEuRbb9a3QDgQQQWPtJgl1wayeqU19BDJ
nUyK3zg7ogNSApxGUN5JyQBW99McWL8JS0kFDOB7o4SBZT7uE6F3W2IiXVE6Hh5nZnhsr8oVxlDS
sIoLSWdrn9MeYMsCFY1uUV8nXS+YIXCDemhpuNMU/0twv5mrPsKxMWL+ZIPAU5gRecTqzpMbaMlU
tsE7WX0v6B3szxQd0wexvNRtz/tgJvcOdAUVld2qhI54+NngmT0kLTgJ8jpWwxqsPL9tLD9ChuL9
054EDJscPwJaQZCqfY7hnhBQZovI7fzS5i0VUZw8I8ODY7oDlJMrb1XgVNeFbE7tsZp8qxsSwvmE
YLL1uBWEbdM2YBO1Zn2JnC6fzJTWwgkcoiHT2ZXyQUP1kWUxJD/ZGXbEh3j8CNLwj46GFcz8cXCs
TwFRzWtvup6WVUWBZzv5kicj805zDbFAz0l7SA69poA0hQ15KYvtMAIlNBn7Aq3IJzP3CT3rjpTG
JsESC1V39V0uK3tqAcej5Mzrf0TLVZlnNnjxP4GK5aC/Gs/PTGqmm4fp79P2r+X1fMc4wV1d468A
qWEuvD9Z/pBj2nA29HXvBs45JbWbnC4NQyuHe+geLskJFe9kBLCBOh3/QMCCVSs0t/YH/3ZQVNg1
ge2aYekkpSjFqBewE2XqSET05hT2qb68XzhZUNT4UKGUeguVYcHL09kgqrb8GzohWJDKePVfX+/j
r9ZzL6XOnOomOQG/al1ueKzOMHkh5CxGebp0Rhj4rXJuLLP/7Wrnsges0JO65B4L8xGKGRP9kNN4
PBewdak6fgFdnYIju8BwXPnkJ/PJ/LUmotC0OoQK45nspFOE04ZQTWbwFu6/Q9YLm2Nazc8uBI6H
sUhT4FGgg7ySPrMl7KoXMTjkKxsR6qAqVDkEZs8NMQCam1pe9OBdlHGOI2Qfl9nfxMdyUS5EBdM9
ENuUIKeR06/U3RYGqze5A7WhC+/6vY02syohqh1aHrRo+5F1HzpxhJZ2MtdyeG/KSv5T0AO8zzAq
ngBVXrDooQNZIwJLOCUrIr1FVRyNsXu1x3QHHcyPzHmYlD773gtrgqQ81MG/0S/EpEkAaoDncy4/
fZ3PsjyD1R0NyT8uMKGm37YNNR3u5Hm4LEAOa+67CrtGLuZZf5c1Zl/EqJjdJ5/rG2Y5+rRAub9k
I+qdX9vBashhQg+493WMLUumJ2R6onhcWKIXILvhXlrmlErBNVjlbunnCxeMSE4sQu/yYCIL5Arh
wHXNXC+S9mJH+Bf65lbFy0M7Non9SdmmeFiNXvRSl85ZJkQrAEry4ySHIxDzaSfpoVLgJI1SVYhB
5uDeDhm2SttshjlMcLvNi49WkdqRZy7C1a5s1mpAwJ4NlpDRTbLaf1VJaGWFWL8zKbTCU2f9E1Fz
KV7mk4payUsKXFRaxTE+V4aW+OG0NF24px6OvES3Kh+VaNfNDC0nwgEnCSpD5BKCVtFMjH89GtO7
wOVowgwokH7PTdUbbEQorI7EghnZJXonBdi4pVkJZr6LcRhxRHtlm029zGXP5ViRM85SiqXJCdyc
UO5LPsEhQWrq+NkqEBHls1ZGXwVMSVGQdEzUOLfCO3S7LjxDvG9lgzA6vA2pmVmCRpdbC4U9vFSw
8xNM64UNs0/hs1RodRZBStC4UU5kCicedHO/HumAmawr+3ZlK9PCjhS8VCbtvEdgJHg2RDULXjqp
AgdI7gzUzqJB/8GY1TySupq/LIyUgFGhw3buoKQ/tMuFcTP35/59aaoONcStHwtWz+jNDpkBHKaS
hBYCnfE/QAp4kpZeuaBiLPSC1/KtJXOjB2GioBRKNZMhG6liogHKRkz6eElg+Cvl5ghMBRMNt97D
XPfxJQEty+nX9dbDnAEVBvfHGDt8sC59TuVVfDO8O6tDQ8f3PpeYwGWlSfMdB9owj6e33dSjKSEB
Zp9iOFcJY4HMzQPibyL2a0Ajnx4AjaPXd/5H3248p8Mg5dCaNf7Aw2rvqsp0cnKtFsiToS2B5oQs
Yl4Y2p3Xrm9w5wQKgbqncFGBwldZwoglU+Hm/yFaOjisgKIux167EEfvroLai5EBJ2ewL8gyZFGf
ZDgMwW9ZLkYgiLIcTX8zJtSenuJOIMoUhovEo4fFdlIilG7LmbRR6Ztb8dHQxuIvsQ7lV2GOtVx2
UXJFtKulm+KNAbVmQDHDt3sgqXdD8mF+Bxhsm0BJKCk41AZ+nANld9oRXYCmhELaQxCRQrJ+Ph2H
PZqZprV7UcOSlNpnEeTvKs8IaEV5ndSsOuob0xSRVZKfR8m0L7mK9gydpqO06N9RaVRxZu7Pc5dU
PccLJJ2NShuUAUVh612BzqbTH1itjGW7p8zTqrGyitsTKDukyY3VNJbjGJMPQtH60NtS+ATrOwyp
fM/PSbaMcKtEiQHGqSjEzJZOYYz7B5X2iL6kdFjNowK9hvCiIjdGfz0aho2ihYWh7zMOwlFUxGEX
Yi5VV8wRXIpNjPzMFDHxysDUNFcvx+iB2nqNQMQQIGnqJUXbNfziJi8wMJxdEr+dBRAIe0j5ltwY
lCEBSU4aUoWuQ+cSEuSNtYvb5SIyPfZuybUNWD/DhjU/VjBjn5TMQq6HHdnMvNMK74I3UXI32SWz
AGZDf1D8OOWVK+guujff4KT/txe7bRQer8nvA91AI+Ok6CF6tCAK53Ms61A2gdlFlG6oDC+v38Ru
ss6995BNPfo5ncmfRbq5uf5ImULMDraQBlW8w03ZzM2w0SaC5tQILLLYbM3Rl+NaG2ppfULznMmv
975sdALh36b7+jfkYkVQLDRWXq9bWjJUarquwg5fKjBjOyhVRMuyTngF04dikSljvFuBVojb6wSm
Fe/w/XEwPbHUKP/T9/59GksAl+52fKKrP+HKKK+P15Zb+fE3cpdWbsGZ3c9AGKX8eHYuWIkfByMJ
R81Jd0OAAh0zwhn0HBEdWRky1xlf2D36i2wZPxEp4V0m7hTy5YI19tJhc/UUoTA4bVQEcTpD06qd
X1x1C0qFkDLTKWyQxbuoKywj/wYGDQngLPZVI/kmoQD1lZjLGt/MJe+EsHMwaW9zgAwujp0wzgIu
Mz4yvR7MzWpf1TQMK/z/4KGVLtyNMcFdgOf3DiEZo8cd74q9zMAxKPIcmybxhkFFx/9X1/7SMdc9
41gVpc9pBgP4FVinDdmOi+jxmYQ06daYbFxNaXuBo4EX07SJzu1ZUSgnrN2N240XSeixzCoCUgHB
vChE9woJ+C5fXeVqyEaA1/d1Mq9B5Z6c/CiGzHW2d2BwftDV6qbtFSblqFT9M72H/yercn04l0f8
apJcvogqiqRxhiE01JNrxTJaAReWcDw1dGb2DJtGXarGquOF4EB1EW59VvOIoQ9YUr7wRXmL/w0O
WJbfE11Ol662of0kLnWJS/bA9Ed9CQ6U0NJpDpoLexkZ9Et7w+0SNewQJWK6t0CdNkEvdLtSBH+K
H9fFRTk89pVDLWMpAVo7djLT2k1B3OJR+JO/EFwCimugsdWJ6sU4o9p+ht4pLA8xDPrDbqls9Hwp
mhUBacBU/JCVpoj8wxAg4l4E86uq2XSM4fC6ZE0XU7Xq5E9Ke2LVCMvCKkIgNccbcHYRvX2Cv60l
FWwhm4V7QPNf1Xlm9JK2KxB+X3M9BCyQ4LFPFf6+jsuAeDtik3gLzxfcrbtQqBBRCAbuRT6U6dUQ
cZsQhXoZSFLgT7cZhJhcco1N676XCsiquQTb45gkLJCOU0PYlJ7WCNZ/23PCm5EJ0m0xGVfNUcPM
zCs3Cg8zjq3hQ/p5lpmX+0/FiFcimEA0RkzX0/GdH6eIvKx7wrCmoC+IY8Kz1NRUUWX6fWNIyqju
5In4GKh2xttEYeD2nanJsdltTYPdEnMp4BYrlxLXRGkEzi+EBXK+eAIZlguBImg7YlvS5ib5LQj/
WHMTuKU4srzV/SqJNN9F/v8z0fQOlwxUe3gCcabMW8IpjbBHOK9W0gIt/VGyizhM0vNKQEFk7yLF
jVKzsKev8mz+pjA9UQUCe4IGILvkN3GibU0sMRAp3tVEWlhRnr7khlegoohWN8DarLE8nGUxNbdM
DCxtxEpO3id85N6G8Rml1Jrzlr8B3BfzGcDS45HmSch+F6oFurBkkoEBxlfNCgRJgrc7cC+KI4oh
vtML6nA2OYKIVLmL+ciqef2yYzVxSiVm9ZHHVPKkYjltewCnnCE1VA1WUoD4Q/2mTClt04O8UEkB
CaiMCNK3Hf9Z1LRQrJQsT7xxQ5zucBNkAnZWGob9Yr8XTngmVo2b3z0UDKofVBiqaLkxZ6VH9uy5
gMCr1a4HwscWKIaSU80X8nsSQ61Nr2tFxjrfZSoszIAJPTPVriwc04JVgge5y/5OZ26nhpvcQTUR
9I31FQKQhBdia07YtD9oPL4MjxVFW7Pg1K43zq7YPBkqBmJa0ogLNCEqn4eXCO9+jMB3GfsZ/PUd
FStkByGba5JuwUkuRQ9R5Fi3X5qSMcqPMpWPJtBFX7xGd2DLA84OgcRdtTWb+7+boxGFZlvi6dTK
cthzHgzwTDp1B4KhZ+Mst9RJDLdRXRDj+CNjDxyI2Z2x3ItOpGS6MqFGxP1U0SsYJR6LWWFY0dw3
LX/PWKB87+kXPjH0geg67WxK4InshNdgjJCYXYHRZJYG3KVlEWpckVJkfLT5g0os7hx77UVUYir2
n1WhPZJW8tAdKy63owR2vLz+7uOglYAAt/S+Jk+uszP5v8zmMhGBWasbWwdWByz+SaKTjTQOeQS/
HDy+Nby1HW2TmRJGr2JnPfhrxkg/3PCLdm7yCc5MhBBvYcm7to8Jqaz0iWMSqJr7G7Q7yTwfpcT3
d/Uz8HG8B9whDRhRXjG7jjw1ty0JUOd1yf1Q9zVgDgnumVzHmmIpEHijDGtkGiDyMxWtRQ11JvQ5
3SfpfFfiBoybJ3Vfbcae9XdZ85niOrO5D0IURt5JL8OE/zvpqBuHXHtAjQObyaAYAAIGp9VgQ1jC
nTKzOzV4wGlIdCEg+XS5uvGFh8Yp+6KSK1O40ovMAQHjsHjPp6/7YsnQ3QqNjCk6hzxo8baGMzgw
grNVbnuHnG8oSPZgAQKSFPUM8gqo0OvtZIzGnPQqhkkhis16lwTNHeQvSW9X9mUh4cCcw3pgOUKx
AVPbGmDGy/5njh3hhifJte8kONPM3FZ2tR91VZW3OJYIFvKoEoiUFXqyPzLXjb+79HDv51jEtF0T
c4F3ei0zfW4F9piedEtgzH5TckbKi6p4vYB+i1IfsBS6KZs57YiRtPIhlaKxPAZv4nzc5bMz10q5
Mg1/xGPGEO6uHrvUs2Yq8BlsDPc/+7OgMiPTcwWdJCke7o7DUDo1n/eMs3RXvJNO6KXVEuV6GJYl
Hu7bA1gewQey/5LQBLeu1Uhov188FDR26vKA6J0UHbGwpYl13mkTXIEozX7ut8tnx39a9aPx3K7F
jCM9hmCictWJQlgSasO50JxqayjLHwK31Wh1/6F5anLxhrYb7/csoxLUxEn25Cryw8Jra8L82byK
mseorReMYCDGNtnBBmy1Hczui+FT3mhCZN5ALsQBXWCpeMJpVNM7Dy3M8Cm0JcDxgkWD/5l+/Q6T
xwgARlXH0xWihVmNZZM9qfimftL3hCgPxe3Go469w4KzKvD0ZwGUl+jZmIUqae08zkrLCVH7KzDs
qhjQPenoS/z7VxETrSqRK+FD/Xzkdvcsgz2lF9eUyvymZxFZMHzMKpHMVg8lPeRWt2TWPGMaY0b4
8vJlTVfPSFbxTJYXi0sYaMLU5l3pPMJs5rRvc1twuEaftwdu+la9aZncV7s4joYK2v2nqgKLGK0V
aYq/YEnJstJeL6tOZp+ae3kaNHv6YUfRroBAybscPh8zMqDeyMNV181dckfw3QZ425Qm9VG95lzg
jWsAp6UpDeDpe1bZNkx4PQ8DG0JLg/PXcb6HOMSgjd2nRCGzVBATWngPLk8qZLpAqzzEFKVAd2Iz
vBRV9oRG/zzQ++F2ZAydT96+Nh33njHebl7gvnOSJmTaKEjXRdozhOaKzg90WlYxq5mmcaMt7wet
L6+LyVs1wSRl0k9xOr1DsTe1mLFJz4lEAOI8+BtaQhnZUxwqn++2tKU69w72J+hAjFRBDREiR3pz
6LBTb1KJseaoh7phcYqsmCWAPhrgss/nB5DdupPfi6h+F1JhX9VN4n2MgZYCn8dzMXsfosfj66ep
lL/WFl+DXckj+PA9WHfljGNXeeGhNXoYZnzFb3Zjjjjt77QBoTqHUAfUoO7RAyuTn8Hz7h+2Hlsl
MrhUxgCrfBi6NZasPQm1eU7DpAmKEgdfa7QBjshpKsgVJDXmzTZgGaEJVSBw/fa/iF7/3Wqf8yAg
cyx2IwyrLh/z5KWNkp1z41xfq6gl2IRfT3TJhQ/e/w1IJSL/6L7JP3i1ZW5tEhPsUTPAf8c/FNGj
dXpq/xcinlqzPrjJiui98tg7/veg4rS0N4xNoTuj8/nBRj1qiBaJBbVab/bi5XIUWRP+rLRTzFxC
9I1S2nr+QfPssKPgT4H9jCADngZSHiSJs6VPuI8dnAsgct24m+kpwumT1tT7NWwUyPSczyOOAji+
W3q1h02R+dKgXxaMUVwa7oK0erRASoh4FHtdmH3299vukJW0ps1msXDrjepKqwIMTD9m2e4+h1wy
Z5OI+yGIHJV+FMCQlLWKCr6FmoJAHpFB4gX62LTnjrsxhOQPJu0NGfoWlpUz33jOY3MgVuK4ZNiN
6ZGoDWkaYRcHh3jPvDdFBxW4XpWZ9JC1dWSvnzCmbpQOIcVMP48LwEJ031/QvAH78lGJZPPrRBxa
Eu/Q2rdAW1g8VaWjT685aGpOUZZly0dBs8xSXBrCRYGQsr4R7BPknxKd3v3I413zcO9x9TFiTNBN
1q+uX/UJNOJRrKjZNOMg6o+78R834WEr7Wp3sXAzFjlJcCOPS5wM9KoPzkhZQnzcXP3PLr8bty7n
zycpKZxUgBDnvP74rgAjrXsw3M6VY9x6IKaQZ/BA3VR+Pjdh5Fclbka1zuU9BKiWIblxzCwWnP7p
X+MFgk4svzj/BuC1VmrftzlL9RCni2BAGmqGfvPgbnWEW5weINluejZF7o4bzhU3/6ez8XWPw73M
Ua45ka69g6qxGQJg1i/THbFwOA5DrZ/IOWLTDgcyHa/iPsGK/VnK5Rgpcr44FyNDoXo9S2Z2Y83f
PdUsCiTkzz9PwTCk0F8xIrykkusZVr5Q38R4BSkOQsuCfjDqi+MtDciUraymkiwyG727xILxfFPn
t/uqwbklJsFAZg6JThCVTz+Y5ePsBXLRnIidGbqcFikMdCUx33GvxmOHVJxCHRidvht7rXYpllfM
FzpLuJX+YaONEnrdLqD4Eo7vIwxmiT8eoGv0fV9JuEN+oD0rWMhMNqbp8qpFsjo8oifXNeF7CiwW
9P5EtbTFnyc7by186tCeemu8bBDAWYQUGdqBYz/GM2DFos5o8WzMs0GVVNzqXLNT8qI2c+B0aqXJ
VcG89akkehXqlfLQsudRI6/ngFiRoJljWJZptfdx1RHNEZnERpyxM7yXq2CmZOaSQed2oQ/qrRXi
NaJc4ZxHHX8VJfc3ug13o7qOImfFjEAFlBotEnl9WV3rAMOGqv0qUHgTMA6oDBAP7Lht/6IaZNoP
knn5cDoWqW1fbTaUJSTZpvjn+bSna3rxMq4LHq0mFXxTdo8DKhy/1sJ/JPzqpvNOakZ2gXguMPzj
K2LwA9Q2392qpgpOlFj+3HUCllxwywyAFaqjI9eMoGDKDRKyOf4kezuzS5vgGw0UXUCIy1ooJ5BY
ztgZOoF23F1RQohCauTfQPLmojW0l3eFePLAlr967M4XzOT+XBDb69bD0JndPH0ePzvfDScXqxop
za6rm+1L31XIdL/iyYkwMCqA4w6RI3548KKE+jc6Ad5SZOHMQhqcMIrLbjBacSuZP2K+ZI5+61FE
o26+2xhUHlAxssXrXz0ba4mtx/8/98EMqdNKEcB80wjRLgqXcvpGqgbSc93euHiTwZ6XP5ifznNs
AohUhSC4gkwIW7BU3kXs3uNJjrEcJkLypWB15XH6/CmPExkILXvDrMeik/Mzx6T8VO/Tn2TOzLX9
cBWFhd2aXU5ESz1e+USxOKQL6+wzmRGWgdsOxB/YfwNIC0DDi+FS1lHXUxj7difSphjNYQ3jCpWO
JEMp6qzLJ4tn5ueF3dLZteUEmq9YxC/Bl+ZBgm5jp71NEDxhUcLpefVInxmC5rSvfPcXEm6BaU3K
/YlsREE0dYDnI3fcWFx5miOQbTUPH1v5Ps3JUgHqC8+jOPlM4Nc+o2fH02J2gKlpyVjIKQFQGzG0
UzA/2MKA20ut1J7sgiruhFRkZmwElQgk6hDIeZbvViuYrsW81leXt7sMIX4cCi7M4/1++gUnmOKF
NrEsY+swz8zVcS93J7JA0f6r3rYeAf0SWyh5rv4Nub8rs6UuoXFbCEvOXqrPHB2heKlMyUy92aU0
xosZ2qgtANm3baRxtYFq+cf97p8huV51u9EODzV5prl6bKwuSrVHefCujie4mo6wtk7a+BBThL2p
5N4m4jlv6XdJe6NWZ6bwKLYKjQsSqb3OmKJif+0KqWLgAlsiIRlH5jUO0LkzYgjlKI7oJ0pHP5kh
hkrYBifYBt36F18SC1PAVWhJmADCOZQUVHGTXHh5bJnWpDVujyy9rkaZ53mHJydBbHL5+W0nQfV4
TtKbuVQBMplcfK/XRs3PTtNFvfB34jYxwCu5+IJX81BZ2EPugUXxd5cS96mduwHXs6vGdWplZOZv
XCirXaGotkoGnvwh8mMhEd0RI9APW51QDfXXB3zv/KaUju+cil+3N4bEscbW4SaPsVR+oSA9HO4J
ycnMVmZ3FJPHwNvIFiY062qWbFL1z8b4XYWCxy98Rxm/ZRQqDwB2HNA+m/gUyW+w5DfQnPeoyUk8
CWH5Vr9/elgVItCIbQe5Gq9Lb4j3EUnd5vK+/nXro/WMdxeo28mpvFaAbFasF1vOZe/CohMyknh/
zietNhKE6R6PGY//W4xhfOX9Dnupi0BHg9vnVfkWpMU8NWBo6Pni0UqdVtDXg/q9aaghvMdzHZMv
ORZWgAN+5DVOKxn8dZcCDqkkaD2jn/Kx44OTHHj5k0YqisnX4W06gSTt158y3dCvcLzKyID0J6cc
ZpPBf47Ix5AXP370OC/gKcFj4F4acqWyS+Eg5YMZk1hX2reJtroVFTzhWPSUwwaTkdpF2nGh/uAw
fX42lF5YDe4bmaqpkFVTs/hm8Hy9zDlBVmkS8UjrS8YcEO8Lz9v98debmziFzeQGA8DNGr5TPP04
ltXiufKmes6mHKUGzxSdcKPFd5xYMtYuxXLIQSVLdiTJV7eRI/htn4nhBf/3GPsl34zRWH3MKqxP
hK8vnNa6OtKtBhp3JGxLvAHC5ssXHekW1troNYVB/GSPlqlwoAS3hElTwSKbljmo27LqIru7CvEm
9ey+A1HLHS58m6/g4DSsNlXvQt3zi5jEY6BY3g6I1xIPlMtBPJJt7PImEv31csrXKhteagTW3ymk
155kehlhcqLIpPVeKMWLG7s56lOMs8jQFHpgRRo7OY6+KE8Ukp8MEmIMGi85pQVQTMSxZQnk6vl0
ReOQyddOhnHWdJb445+t7pOCk2FBAYePL3GYjHge8zkJZjCxMkps+Z8ov7BnrDjgzQRUxSd16zbO
bBESSjOTNr7kGRaSfj7R82N/dqrMlSaaS0/HM89OhE9IXYdTe55gc0MuC6JUW971zeZHe7Z+oqrd
QoTiHp/s74nqNmtV0j2mmwUUUvhowPU3CROWbiOZmzBHLu+Jzpy6pbPHpz3cawZR/cAk203pzA0h
vFOeHem6WnKrIq8i1/pqfvv8BYWLjMI8KzmHBBmrtMIUVfDOzNbEbnTc6ppXAcFFXA2fgkyhvVY/
S7jtZ/ApdQdVkI/Otlwo7RcGHOD+XhDIJ/6Hq+jBPRsep4wueQo18JL5Z/p/ERp/5k2nD9jJPoMs
XuK+HvNkRJ7C+1Y7kD86AF4P9hCpn62MXydUOcy2VggPYKQ3akZWdaQIAbTRiPbX/d6OL1LQ00zW
TElWp46ioP9VAbvNypKwQ7WsyeqD2FJ8IAd2vQJKBCk8lfD3GDMddjiUmoXQBu0rViqr5V6XIrq5
p/aJ91HmIHZZJRxGmGIAyWDf3qqExkDvYpXvvsUlkhwzwFDb8C8GCXyN12tCGAYr5yfv3jUm1Ik2
w8n/d6GHZEblxjpMFNZQWSsfr3VA1/iNkggYhFQq7BRjso0qg1O5boZoEBlkU0FmwYZxGG0PsahH
wwr0doulRr/p85nPmEzqPJ68Q8iRuIZGB9sUG36ExgtcuM6sAL86hD0jCwSnLyDG+i9MfX5qG0sw
wT5DS8LAAI39IjWD0tF2Na2pM3ISM/Yrxvei6yG8BuMMltrhIKd9hCpmS47c1HL3OW7cF9pyWGlO
6Vrx+lsaYbfB3DfRgJh/uj4c09+Fraa5BiFLPLmdiT77vwq6IzrXDb9H0ouTkiZlt8nfYcKG3kU7
x0bN1u2/tXHrGJSbclyuc6ZT/1e+yQHUTfs5A3RnFjTx9ngXwyyKeV7AUQh2A7qjp0HjTTpLXcqa
AGMvm9fDkb1COGcGWLGW0M09WBZ++WKLoRceq+6iQYMuRc6+NTXXIADq4C5v75WL6lG+S3tsduUK
Yu88d3JHfMEvdVAyt+YiyS3wbtzUMv867LJBs3EN010KI9YbzsC1mqnvKChEqT2zvnmpAa31N/Gh
2nXNEVF0DnYB+BRjNm7TTXD3qFTEiXHd5foXOcPg9xwXwTHFTa0i3m41QdZOSU50QgAEfK6AApzm
3OAT93BYDHVPMpWVEKXjHPdWADhE341UueQ6SFLSU03b+BlzougmzrOlYmNE/VOa31IRE6FAglGB
3eAZVcMOnFIMGW/JbL4fmwvYLICtWHrwRq5gq/5pKTUdbb+cmfzBGibFt0nPo+Bpju+zdZZe8SD2
JEF/PKV126UdB1JIK/IacM2uuUBlN4q33+wKjhIi+VTQCmPwoF7+6VO0xSiifZMGJDQ8ORzy+M6u
6ZuStw/wCpW6X7oc11f3WOpxA3+v+GVEsDJJzUGKHDp7L6b12C7UdWitU6xjpYosRsac2+casaab
phD13CI5rPMPUwiko19f9QSOQfhM9EIaC1bi5CeYpqIPo6vqM/OQ1kN18gXaFEJTZ4onrAuOf+y2
qnLIKSJQpG8vMfEav9bdjp543MJmMaPxD6IgTWSK04glRt6ilGydWluMVq6oqJcyEhYsPK3Car+c
LnMfWfNtopIRUtzBDxPV5MDN4uCHgwNlOla+cSRzOUtDSkT24am7PlQv29z0wQ6l9oiHIzfMKKFD
zyigF+OwlFIHbFxCC9aebj4uiCYr02SsYTRyQi8zXqJW0LMqRadREBPz05RZfk+LWnPjd/9EmPFM
yk7jCzjH4ShnuJ7yXPfUhBJHJUoPSE+sCNT+N5zPO9T8IcckYqGUiXA/FottQzt48lTVy0npCdlz
jcdroX0y4W+He9OdDXqk/J0sMh4d8jfpYLxn+WGHzUTpTZAKMGykE1ZPvcXmZ0PvrYVzUMdlQ6sa
FdXWD5iiiFfexHl7NXWLkkdjuAGv+ZqlrKpuxcFLy61XSIZIxBZgwSlSOAeKXyavkQo3bhMS6YTD
788ZzDDV0dvSYFXemoGVj8hyDTVCOeKJGYH/zs1TC9+jW0DqL6CkMn/TRZrd5Qj/Pk9orZQ84DG7
+Xg/YTCNpBh89bcTJFUQGzhrMAHHRoEj+2Wlt9rCmh46t4eoJa4toVavEhyQMP7IKPkyXJZc0V3V
EPpbu24rip+dy25+76YEtO/jDyzr0iJtnLVRfPH5Oe/Rk5bjL03pJlOO4rmiHTmM/xaDf8aOr2BB
QGfQx/cQuW5pau0CrpeVHesJFgETqqVafSb7j1CHUMwwzk0mjffxFt2MRRXLyeIdnVYs1YMbKE6s
UtGonOfaoWhNyiURHLl5yibuBdenM+m8vfp645XeS7g5IIwb/TqetJGy2q5tlNUtrluHdhAXonBY
wGh+LWqWubHUvsUpKqLd+FVTOcdNhknagPkIhOJDGn7Fo5wfxiPoN1sm1wHohZ9p0DCkqGKERpl5
aWYAZHVnRzCj+AYQzBljbrAO2bDTJ7gXO8XWOrLU1bDGKjkUz1XpPYcchad+p7ZdVKQqOmdRDfAe
OkVeSX0EeoxxeYBrZdV8a0psBzSETEs9/fbe90L9nFAa+0oeoTo6r3m0M1TYc99khUgb3y/kHWWA
CXZxf57c7K9xeXfYUxgzZ3mbbBi+BNq0E6ltm4NSrm9TYB36KdI4o0vueVTVrUI/UCTcsNmO5R83
8RLXHyMDRl3wtn/nhOUx9iTrgP6wOuMH+2t4FHOnR20/nxa5Ak9LzW1HEPIYBk6og7QiET/kvIRO
op4Wgefd5JI6Ka2Aff45tl/zmx8KzgwugE4yLOG6/95WamI8T0p+8ExbQ06RYvJSQs29isqKOz1A
ocwpQ5MPTcg2hfXfTGETzuoTRbvoivoJ66PM3lJ+Jmw/v6DfmZScK3W6X4XXBsD/ev6Zfwb7a88c
bv7AG3rbshg1p2Xz66ZhzkuJq4qo1h3xKvV5eBKTqB8nilo9aSmjiu4pjqIvvsh8i1M9FHZQNv0j
i+Mwz1lhXiMSuwvR03+s5OPAa5EzUd4qVLSCnkOO09pUdrxFU36lTetdtxp1rCizf44icFu04p2I
6CsYr0CWH+L57nV88fuy72CBMpBFPDUmVdVmmP9TAlvUvi/8dQACvayHY3qDgeKy+ouyv7qY7QIu
kpojQ2CMfo/273aUR/Zjim10DPurhYdmOuAk5YMaJwXkFXjuwz4ZekMyoR3/RgGt2CNLB2DL/0MW
K90BbJTTPGjpuEdPKZ1SC/cgPxNskywpzphbGYw2A+LWHcLall+fdWs7wEKKijiBE49N+dum7XoJ
9cjmHhmEwzDwG/m3/K1dboJH9+Whe/SPKR0gMAl31c6qOTrGMiuSPi4pkGqvKp/yZgMy/7nOsyg1
W8pkQFa3l75wmUE/gdOTJnApuOeOfLeXjdjqpuNHtdphbwuVa0zo8L16QKyuhzCyMQGAcGkNEU2O
kGeNXCC6YagWUBessf+bfHOF7YRkQ2BZjamp02c7t0Sb6xeS/7nP3KbEO7UYgU97CO4Z9gw6FAUg
11po1KqSV24nZzmOROVLFWHnba5tfd9FeLP9flM+6eKh1jv4ytmtCowDeC8dfZVG2tQihl6IM/cd
qr+PqhH4HCLwU5x9A4no+pukWRiHpPB8b4QxWYznLlGJHW6xiSGPdEA/DOb8BSZ6+bpw7EOZ0wAS
2D3aiEmtucyyjDTCO94Nl08TU4jozeo2YqNw5g/A3SPjkm1A+kZ5wOyONGMCcPxKi0vbTPMUFRRI
pSJ68OacH9ifBKMdzAZ5OV0UPPS2Oi/x4Ou89Uq3U4bTN5Mv/ofntpM9GefpBQLoixHfciFPXsgO
yaBkA/fuIUfB/2hHA84jBUyPMXx8jv3UXt0AuFnbN2L+pG6Fu2Qgg48MOhGS2WOt3g6KlqEciT+X
7vDBWx1Q7SCpfyp7g8k2XGlWdzBIdAQGznufaiuD+EpVBuaBTSwXamOfNKiUm/wIrMmyw3FOUsY8
aJ75ahjFPWHHs55J96fuQ5E6Q8RNqnGfhxeJ06X6zEs7wX/hrwW6Hwl+qy6og29LPgUVjawm3MR/
WZfE9KxOAA6KS2TO1DQPGM0lo1mR/Z9Hh/CLJyWsfAihPmvDDuduJciH3EXFZUG2KTjweMxseD6Y
J0JswTctu0r8MfLIjxUbD5MDWZ8hrnWHMLUHbiaf8nxDXLgY+U40ayJXV+UoQv50DWpPHW8DDFlt
Ey1QMNy+kifplWTGq/5RNezeerRtdUaTRy/e2yyVSpcvs1U6Hs9m8yoFhmUCmx4W8J9HyejvRbse
vYFHnC7S9NgGEt0Tftxz9PcR8vPOt6gYrxMQTU6uT2k46YON+9X2ecDcGXyT/85YOdIhfwi5+90U
HnBC/TtIeSHLazlWgeXbML6Fzwo8MhKZDEVPrsW+QBPcliaQf9U4A/mrxq9H/Orry/34rM2+7tOV
kQaCMcwYitCKUfmWnOexEIB9F4mNhcwNfwiu/vahQ4ytcKUJjnDnBZeVaetIJ23vJ7k75hSLFf6Q
CW+o52uzZ5atMuHy3Qy24UMbUpNTyz7aCS7wUK+oXY9hJI3Gh5BqDZrMWi9PEnrzawOsxjhkV9Uy
xqLTtInALclkp7RfOeFU+RgkQh0a3LwLTw3Rxrr2x8Mgz3tIGSKA6cm8f4464Wb7zHirIda8+2Qx
oPSXwnpOys/UIHWXyUewLTG+QVmoofwGJImMh+rhJ8NQOx6xteebqoeEaz5pctebiCqktKa0b7Pd
N6BGRM8AWo+hNoQL8miVpGrGsF4pS65v3Hff4SkChvHYhPmdporM3yWSBnlaSccFlROfu+w4yjXx
wcFZ/S7m3u0LDFtMjn0IZ9AZDxC83yiQnjbK2rWtqF0+OMNDiNzYU8LKkFFzG5zQ7NC/oowN59PX
x1TuwqxNBzjTVxnVoEpC0jLZvBS2BYDnFFSjR3rMHo4NtWTEdqjbSANu+mL7Vjq4bJK31zCon8jj
4M3pe0iM3dyX4G211Vk90RJ9mPnAmYlQlDb8Ly+ifL7v+kRp6XK6zjybLqpoFNenXL6k0bgEpjMG
lXgSJ1RLYbJDy6QtQZnDwz0qbkaWtKEQ7uHrXyw/BQvXU/QitySzDEA2byLvAAAHJqMWBAAnhJve
02DCFrPTqYZfhqovFz/iAJRsES37qDvltxwt9gNllgjq/05TGtfeXgL2nh3iReLkvDesAxlqeVn0
s1l7ilQtUKDDhknARRRe+VbeZ9itniPQCfGZl0CvoUvh+x+ze9biYYeL1fSGMtDwhXaSqczKYpeQ
HH8qapRdHPJueWHVfFD5rQI6BsXvjUbCCsndokDxzLK7ZT6WwHNVoDIB+d+g3F05hexqxTvVYnEt
fQLphmdGSLFkG3YRwK6u9ymAETyhPKutkp0CxilxV+mNIGW/E3CFYvYRxCRpfUfIfjGZqrNXgEEH
+bOjZbmL/GqZmg+g2U6im7jewMwxl0ZejalqAe/E+E1A7ogkmypc+38gGXkKi3uxf3sN0ZtahRZJ
HbGPHJGZXufu7hfR2pt8l16e3vDrkgDw0f7eqUYRuIOIKvJ8afcpnynC+grZ2nSbmViJvuA3VCz2
ifyt1bxElwezjwq7OsywNuFdwDQMtDmxGN8ckcsDJpeuN836VuyHfjqyRhto3bj7cgLYeUPRJBVI
dWIH72hrdoPrY+FTcrRtFGBQlPbFGIK2oS50A5NUF4PknkdbXCf5bN3Nuej1L28iPg71H5ctpRBX
XX5ReGWeYF+NRogKtPvt15y6YRqHoZXwxN3u1dABYNdvhNLfeLd+9iRVdnRu7EL+HHnGdDtw0nmu
p3pm1ev+iPAIHihK2iPW6Qc+lBkXSp12u8hwdzKhbPmbLG25V6cStqjgJyBxTTfrF7WOc6AgOEJu
hVZEiqJ60r4Y+J69LzyBIOJ589ZBsuQo4v3i5GUK8m3yXi5WkZyrl9JmxqmqXlDVNzlHtdPKdwxS
btaGyqxBmFuM4jTgCE6SmiRrUhDrkPdIxM8yDlZ9z8vNICnnHfLt7LeaqJjwfUhTZI6FQ2vypZ/V
TaCDDD7J0ZWBWN3DKVJuQxdLYZmNKG7sKx9n9xl6I3lbQJkuE1MKZfxuTH9c6Pl+4zNZlGPfyl+u
EL3MiB6MqQGYKm5bydlnqJlSoW5OnqFj5X/BenRlkTaeeKLlRIceoGciisF6qMTV6BQikqVwrxZ3
2hIOD90L0q6SEmFKSowtbPMuoNOLkmGDlZ1qsqBg+Nq7K9hNWjxXuRGs+D9FAG9NXeOg0QrS2lA6
TaHgIJ3AbL3yOoR4/KQgDvN91I7o+j27oIhVTuznbIiF7q495tG8HbCQ3w55UuF55vTRbMe4Jh4t
Ls/PwTaKtZyoLQ6ceXxQNQDkZITjPs6WyGOOdONUgkRCst0D3j59jZODn4qozunY8AuWh4/S8Bay
/gPvz5LT8NVfPUdYYlnFEt/FewruUDLCNV9cjjlxiMnukFLbt8ZcXBjzVc0xKg7zf3SEsoKkf1u5
VIpJGVviWH9+e5Uni1D3FipIHSqnuNUzeoBiiEah3UiEoVF522aBxJGQJP076iHcnXXbeLdKbuNq
MElQ17JEcWpwjKVFVXTFPMB0eMlIeuQ2fcf3qDKRhbMuc2AteumucyUO6J0wXCOl97RmdbFcDBaX
gHCNuOWENFz0TOod7xe9WxUOm+rcpgK8WZEpZdyQ8CUR0cJ/mClf9ss6id5k4UAsDILSUDblqZtC
FdWKhH/bzYSnpoZYEfo0yRD46gcU+Pq3x4LAePNRZGYVdHwqTGSXman34hMGNBP4RJNCBs7XkK3r
kK1iFmlH71bPFGM+XVjRGP69m6N8J10ATE3NQBumU2aum64gozly+PiPmqnn5ysyWjKlkZKIa20A
VPszvKUoUKAbe7bbYP3ooseHI1VKfHZzmdVXjIhi2rY/fIOirwxVGHRZzHNREm37IMXtVawpFl29
mEvnLzCyzQ6SMHz2yzsCXHjPZjN133/MeIm4V79P5jX824TXKowBjw/dgD5PG8ADyc5uXtLN31YJ
DH51xy7JQTwljI1Uvmq3E4F4URlSmqFeBFpTyfCbR2jobrNqv+UbB/V6sIHp/bRstSfUyzpgMKjW
iqewqJQrmuvWGWL31Ed1+l0agVC8j1mR6OqKHPBaBsNz28MR12ZCLJz29G0QmHFnnSbN9lnGlaWQ
l+PpaQ2HrmTUXlRs4Oi9hWffYb+30Q279oZKX32VTdEdRwHYpIl9NpkD3Z8CUxroivGLwm3G2f6b
9vtutR3FwnBtxzzI7ATWEKfozH0nTiG0giPwWzXdKi0KJNn1jqd5wiSSWQMT+g3ZNVuXBiTP2ucK
3UXsRLodK8knzwv6Cx6yd+QQUEFgWPgCCktN5mBNMI4WT4SbqOtEcuniBeGbbE4ZxYVGBf7xnSqN
xWyTni4D4A4Uekmx0mTpr6PkxpIt4tH5W9gtcL6fwYQPghM2AgY17jYwRFulFFrFvUn+OT8su2qh
lyusg57xQNPnivwEFjd4PH4PxKdivaM/LjixdFpAF9frvtuCa4cefoU0GhgakaGgPrlH7Oml6yJv
u3qGKpr61M3tEqXV8+GDAvYkpgyLqVUySKsMMiYwotlHRT9MjwemgCEdiaRzAEbrFx8sZX4HuszJ
G2QSn8N9F18f75ts3Ha8wTeI93D3u2uQNuvx/fK66JYtlY0hyHa+6M2YPVRR2Bvxgxg/E1/K6+xC
lQnsXMPHqJSRlPKz01BCDei1RQt1NLW1xL9uwCMwzUfjx3Gjln9GrdxLzQouYiL4bdGoTfnvf2dU
iEPxGRsHhxvtIRif/yqlIlSsvtc4TuzFFtYejq7Ks6dbJk5QgWd5gWZSP7tLGshTS8QzUKJczCbX
e+/Z/JO/BujFpxiXRvDGdU60ra+TKUGpou1pY7TM9SKA3WqPS6Llv+FlxFzQopQwvSglgjVP/sZv
OFCLS+6+5GyGyt27MkDAZ/QU0HT452VT3RXfdoQimu7LRBOl07EvnrB2MsArvnMxPLOq8PO5Aml0
B6qB3LaldKI0u7jcwbX34KfSM2oP6tNOc1oX0wyiDzmrbvKK/OV4Vs4dcG2mLlh6SAKeMOrTRL7w
ha+GZnjVGRtQxnow7f3ZnViLephv148jbKJ7wuk8msWbp6hXcStV0bu4LxKqmHTCg6v0vUdsrmQD
dYsjYZeNjrcwaoZqhWNF7BCZBQEiDUhfQNFdnmJt2RQ6rFkc5IyjkYUt0qihBvRN7tuclo7ZtMjC
MONb111lfAn/KntPcFmqTC6r0WLpHQ//MHBk5ZcUNxJP3Mhxzbvu55N49vhM/t5jpMgAD3mlN3CP
DZsEBkGor2vyFbPDg7JEJV8vTaG4iPfJA8Z4lK6eXqyZTpKs9IHp0VKql85t2q7oOKE8KfbrGHRN
j9GNslqHoT4RZxtkA5VJUGGeOsLOuCY9cgeviT94YBx1ubWm1tZOeLjw3KP50erKKToOKdIJNwLZ
81NDek0eGfpTpjYFGtlJMU9OiQz7Iz1TloibF0Z/FzfmQoXXTHxOkVCvEgoryx/axUlmi7ISeBRb
30TH2PWdeKrQIGJtU5wZd2Xdbc/axQ2vukrHWNgKu8UrsITfgoo0UYMA4945qoEvTs78cIkm9ILO
STw7C9l4J3BSl3BGv9a6RgbJ0qKn5OKmstzsh0oIA1lz24rGv5snBuvfO13rVcv0Q+lycKRDocXZ
Nxe8TPlyY1Y+DGPZXJtOnnO7H+XSM6tDj76hwx0QCxuuj88kKlvN9rf3twV/GngGstj44peXEwEj
i/5EErjISVmCN+ocQTEDuI3dHt03uJ+9vVxz6D1BfAdKnRRgEEtAOUoDaz4uLA89SMEZ9iuIJ+yW
GtyzQC3kNl0PYRg1H6LoDy2TnSueZTxL+6SlPZKF4Myb40q0PI90y+JpZcAftPedDbHbQVW/eodT
hvS1kwh+GhQhXj9N7hte+KD99dSyeLC6W4ENDOb7vL1BefeWDtEtTLaKaRy9fhbBFGZLXPa1uohQ
Tem27Tkt4fOX+fwCJ512+xY7d8M15qBUyG22aaGMRNFFaHXEikJgcPAiDjfGl06D49/Rt/huJBDw
hhdOb/4vDd97mpjRAcbv4RYrW79r00GJAAomqvNs74AZTl9BUlkGFCd1DN5sHSP/Qv1MF2zF6+d7
n/lAaHvss37yD0LF8mRh5HUKP6Z11N/5hgOm6UAAu0CBqQhMWEeTgU/HS79a5N6kgFt5ocrw4HCT
dkxaPbGjhcSbFkQzvVkU+ipUHmBwRlOY9IBwAxsLdcYphHT9XVsgHO9IZUavqn1FDuTc1+nohS0l
FCNSXOOLcf1DjpyimD0KSYO99zgxtf0rcCwsqg1QHcusTTgs9+G21aU3rD8kk1fclLCJj9barYM8
rPsaX1LGHnW9AeBYsOz+vU6fYPz4m8YhYskNjwzjvh+d7Ix9yAXgpvJU6NlSRIjfFcpOHMWjvsVk
jbKsnOSvj03F3d++OfAWUzj6DqiwEMzdAK6MRjkgtNWTK1bvPnKAjXaB+YJxAjHloTlQpLWGcuqF
C7xAvgcoaUM8gbDNmoIMPhEuMeIHhX31Q8jNSCtncfM+isjUzcQqGj7PRA1P3Y/KP4yBmtDmU6sz
Uxz2mUcxsRwiSgUiV3yua+skAbaKD9jTSjZxaFwdjUQiQcKSucM4/z5QlQDJw1bKts0jxJaovbPh
9wPCpACe3wgbe7qZN5MqE/IZoZHsxG7Sj7mOCqSwRJaW7qnT0O3HdoZJ+elPrhBvSJyYm0IGNv+9
dpDoD8PdyfRaQl4dpmrLS7hav7h+yt6zSeJITZtAqSOGQECI0fZk9PbxiUqkScWapkF70Dyvx2xs
l98GwS16QS/N9QFyYZr5GqUm01dBLeTFp5NEEEtOcxxIr56Tilfesdkd35qEJYacd3+6yVLGn3Ha
seJCiGyRR2ODLJdXiknootfrlMZvYvKsavTEyYpkdm8rhEWXHy1Y6KyOiOUgzTE/xtNa53Ne1dy8
aAgSVMe0OFdcf4/I2N8s9UC8JySoF7zlbb+IOMpjPauRbXPlkdkMbmL0IkaMX2qw4ohb1tGPKwuV
n3ZJILA73L0XfqxQbxtT3zyNKOojUKNsEHlvpmuAjB6+D9wYBV3XRG/pLcZ+zoSKwUMHK10Vx7vu
lfS1fGRimOQl7HAqP8km0Y5Z2zzulVCVA9UchSwMcR+RDqs00LmO9pKgtovBVr0KnLSsZxI70MlP
La6fuvbDBJtIeEJ60MMQnCxfdUE2F4RSr4Oy/Mkq/WiKOByaM913Kehf0lTpuPwCoMS8aVV/uZrg
YClamaea75PrSw0CDMpn7PmqiLuXOt4DAjGAtjfKk+JeiFr8mct0Adnn/QfymAbYqtADO1C2BqFz
FQNnaK9OXd+BkDDtisT62Ks16mjqj2eCEvizhfKmix2+D7DiTNBHXt4bNAEpqEwgKajBGaUNJCSJ
i9lfBCRNVk7wqC8f87HxS1zYwnaiGIaDbEbI1pMVB8Eg3w+O/bQN03xvWxjH6OPd+DPSdwkERRUz
dAvyCXq9Xpz1uVfSSnvFsPKXXU13xKpelz76tjjHPAebMkz2fOYzWn7GMKCXlD3osm5cxwIpowyK
a81OS5HCj3HyGOGzrmAbsbff/jfH7GUz/xmyfJr2UK3oLg6CH69zcVd57rK3z3MqfBmLMvX035EH
eICFcnPGGCI2ERnyy25ynBYp4/ee7eG2ye2po/vEZ6wlu4Orid5W6+7PUKv6Hpf8yA08p+OdoJI4
Ejc7XsOsKgDQTG/uqMT4NBMroejmrRRgRu4Jb7wwf6MgC7pU+9yoPwr2NzcXLhSZZjjxLYq8fMQn
dhH+S5KS16cEy+QgoDxrQvSD3nuTo0MkViIQgQ3umQjDm+IvnH2QIiYYHJjZAvyWx5bSAIAQiiVv
p7Kr42JmZi2hF9XWVnmFYQ/mNQiifiW2a8JjPLsLm47qv05+HLmq9gRBl0GPrt381sEc87yuiLO3
7ProdZ98/7cG8UXTWDY4H07JwaTkf+VvlTyDnevRVWbsLL10KbVi9VbqmnQvrO3Ih6ncWkSnvZB9
VqzvMcwBSS1r12nSy3II8LD8p3W1/lLWuYOAZ/AQzCPzPKSM6HDb9iYowUhltAqmZgEjFyNOGcYt
GvStBBc4ULxYbXRfPL6r5qDtBly3dFdhl0kLKeH3xXvC8Aj//kDsKzBK3Gpe6qP7FUsYiKz9olPW
mIdX8GG2M7Ipo9sh0gg5qF6CMm7yu1nwVnWhImC8EGRsuXeQDfyPhyO0qV+tK75tkqiL0jc9FtSD
YCdE7aDpBdQwRvM+b5eZ1LDJiSViG0SLC26bUsgWWfnWzuPLuXiftph7AEZ2Yt6Uqzcayj8QEhCF
7HByP1WbudM6DmH/yRXgJpGVz3VU4bpzJErK87FJMi24YH0GDY4ru0DUmvCKMCLIdl8oh3fFDnEh
0vHQDereVhUzo9K/lqLdCkXE5O2tOprpIldS2WGDbfphpouQZisHbLFc0zo0ZA6j5lavhozDTbGT
9/Cyi1rzij4g4fivxubIc+wDgW7vjQMQ9W4zJL/mhFqSuHpMU64mNzUV0g3o7MTj8BObXvp4knVs
S9+9lZpKe+0bx7huIveM+c/1BruDvn1Z0cXQcv40zpBtaWUN3NLKRISvAif/4RY8brDVCBdvQj9s
h8IB28Cf7770AazP7qJ/u0KQ4wtovL0SKy0OT3eY8qRgVS6l8+h0l9aWWW0qAPQjDQ6w3YzkiLC6
RtM49w28kY6vJfU2P5YhdF1NQINqTyATKSFmIay1+KEOiVf8aVrmLb7WENlta2ZYLxNocZfeqFfY
1y4HQ6r0xVyfjJu5zR2Eq0T/+E5vKCORHQWgxAV3qVps5+2W7YjhKaizMD4FGiVK3j6LZtuSNQ0R
3T6OKXfEuWj67WE6+E8FDSEbdvGVElYToEu4DguQKEJQGmdXAfmy8qUbfX/POP1R2fr3N5wNbjyA
c8I77YTljWRXVzNmLR4Tkj2W3zB2NpyvXNP+dLVINReLiAbohV0nzGCy9JSSkW1VZ4pf+DKOhXve
0jkcK5uGApPxUjrC0aBxAAkCI4swviSf2c05TUkaZCbxTe3IsgmD74jCloYdjmj3D2MFvCudo8FS
WLzbGn+McFos5u3jusI1+YyzPQmDwVZsJiKJ0fD44cLTJ40L8L57wW5YIxxJ6eywFICcD5pkjsId
mMreLAHzya/hvZEa7kV2NoOOUsbC25DiMMd33gRAp8JVdYTIF4MdQeUswoOa2FWZtP0LUh7Qld6s
TFOmOjUmD4Mn17WJdo2Wug0DAWtsJPAQWKs8Deo8TYQXINIX12v2iIWMgtwqiuCEN89iupENl2xC
0250LAdu0b+zAV2T9c62GNvGpQe+XQuqQyzzcvinp/+RxpifL6juuDDXy+y11xrFrCeckoaDzzuL
YsNQZSvdyYDNMWIaebIPLmmCyeKzknpe5WqllUbwkX9yqrjTduRMok+n+6KtNdukwruN3Y4IMtWP
VacjdBcKgJLWDCqE82wmQNOeSRkg6fvg8m5bS9rkdPkyFpDi8w+Qx8cFAMKxMXCMtSfAL9iWtTtz
7LfKke6bRAIy2uzNiUt/QtQG+PUeVA6UjwlN+9RVZmklP8+FmHkSuOLk7YeWQpQ2lwoH2YQ6J8rL
YnEeb5m9/wVOIMjThPwjlhk4YnjK5SKmB8YzqRjHp9v4nIbsnvG1INOTKDvKdojpPy25u6ACH+/t
RrecW7nDd+7bHFJw0+x4CVNnBw3O33K7AG6lDUoo2lPL9nspa8ViAwXTg1haWNpTLf5y3zuLHNwM
4IBWgDW6v/elm3yFFWbcrqTtatkPo4Tu0NsU/mf3aJX9wWJ382Ew7dn0xHxE7d/s/24MFuPFc8lp
VdNP5qsj9kdJEv7LgI1JQjst5F+ppWDDkcF/Ol3kcxym8QtxPeVtvNxM/SzqVmneCRaMa70Bypjt
HglWnLmnxtyD5PedGeMM66FNKrmORRvmRvlo/q10R5XQy2Gwn4z5bj87dDjicPRXLAcaNemwSVTz
PQ48AsD49dLvuZnNAUITMngvgndom8vBn4HWBWeN42ojvhXxNLIv0pr1shH56hMiwPu2WWFoX8FJ
07RvNoylgn73DpX0tllcRxDErVj7luzb8wkAh/vMpTvLuy4Rzf87ylUwPc3ugaenFnlsaOjUb82V
yRnekkgFL03+sarGiqN/GkRTyfBmUHGQNsbyYivOdN8nYHnoAelveZXEF0mI7czYZcaSXAFBwgZq
3leGJfDD2GO2OxMFAfpth9IT+lW8q2BGXeRGEsBttjjpBOVEYhGc1uEjwApv1hR03GOkG+UIaR52
53duSQoxBiJh8J+ZkzlVy8oQPoWY6MU5lXb6wKEVh5b+m5kOLylQduPa3BpPV89abmgJl+gD4yi+
IkTj5OI66Yyx/FdJkapeYPl+fDJc0oiTiYCIfwqTOaVURxgWPy2LFurARRpODrpBjGC3YkhJj2SI
yrJ+tDCexvW5ow4ws3+FD4/4pN0eR/jT5eTlCNvd2uKcqwmlJ4WNRg+7Rb+Q969ot/9GD3oEqmMu
zhfjRUGC3RhdQvQDl8uIhaed5AbzTJr5xOyeJPVmxRqeZmKZ5gUshfp9h8TWG9WdxwgfiN1JYgbW
XzRm/z4B5MuEUwRuUR34bhVENcA3I7IOgu9bKaf8YGSa4OcFKpmeNklcleQK33MtjLT50f3Ap9/e
8W1W/yJz8NNPABLhIoMqJT5gOEvYF1IL2uuRNd5GR7ioFUv86FF3GmSSzpqWtSARA/5z7QPxRqnm
P90nHXAhFr+sq2xRRDqFqg+jporWYlsmfULljAratzjl8TMKW0nGkiqHU0ghWsk6etB5O2pQN5wH
s4hoF6WkIkEK9eaCHx6ZB17820zvKFPNVrySSN1qh1t8+9sb44efF7eVWshfnYNZZLk1ltHb9ahr
fNCYh9mJvGmELk3ih9KR6CcxEnADEBvXHCaJoRCq1vRI5X6rJ/+5ALBnjom/pERzdiemwUjlIu/A
GCz4W+GhQTa0v/wTLCJ/AflthoDhYQvs+IrKAS/ytKDUAVvrnUIMoBghlP3ri4C0jTxO/+P8DfD4
jEouALSmeskzqa7WJ/gcMhuixKaskWpVY1bAHxDYVgqMd7VKltBduB3pjMlhSxO5kGsdJSBBDGBm
nHlusH7tadeMUX04KAHJffIG8OTrqGh+EgPxtFViDgIIJqsLtwOaRcwFNaxJva4A8esFcwVTrHe2
u3On9QuvOA62tK09ZkAX9EyejJZx8FFfT8nYehXHWOEujeObDBMPfXKzJcMzj/mFAMhnY8RLMmuU
MrOSmSIVQOsn3Xjx/t8WKu2cZnLoA647DZVDKepEnHjW8oYpL6Wo3cdUg4T4kW/O8oDRx+87qY27
MQiNojR4cELYEX7KS6bXgmJQgUNsDguFimovjMi99Llo/SfWIwXpdoMFRlCK1LdW4S7wMkYucBva
z0N9E0FAuB7+J93H5UihtzMdOLsFMZFEM/2OfBg8izYuKJVjc+hqHIcJzi7G4hhX8hqMEAGx9dmg
TgCsRedYcXgKlQgu9QZCRKe1BQ2cvnInqT/Lg5KSubkaQ4hYTbMl0pXF/5UX+vryodGoZbolg3ij
UPxFeLgcyplpnvZkx6fdYF8kT6xw9X8UiI5sBP7J3froJXucsKww4/s0gwNQuaoD/bpwNHuJyken
Ppy0YI0ocNwNnoANK5C4Kfj6ZPv2Xi4zoeaI5Z+qdw+Blo0O8OINpykHPyKaAMZdQYxyWyemzXar
7so6Rh+CISJ+Xv3NZ39ET9PDwiNKarQ1hfVGcAgluzpOTySss0Z8nLUIMlSYPFcdg554pXJOSNty
RMTZSceNGabtpTcKRr40UwrzUef57EStcLz1unGtT/fTa5YU490Gg9kZLgSOkqFw99B3quLcarUm
U8dskxtR0KOQzKKbHSjI2KMuFeLWc1rt1VjRs00BONrvEi+m6XbLXHgmC9mXwjOkEIhN9vZjAM7g
ccYqHA7ZSNRql/S/i/vXuDElGWnRn47+fBkchHQMz6Sj3611N8JOyVL7FwB5NBcQHuBBVsGSoiut
gvdMf2PnfNLFswSB/3LY7pcFagKFmrdMuGwdRG5gSBy9HkCAaVPsnWS/F85sd31j6vZFs2j45sqx
mrCUUTj8ahoXTYqwqKk0dJ0+j29Cm3erI1pXbunCnc6/NvKK35cptwCrUWWCcgTk4/rARAisKE4i
Rh+bKGB/KCHyO2y/guncvTgjiA0jSYR2TaAA0Yz+2kk4XGhQrlOzExhsYPm8VfBkTfnu42Z8nHYi
Hb+4jGnxeLvorTk2gqJqZ+lFqfVSojHQ21bIZ1qyIowd7QvF0jJ8fVoyu0RJGStQ+JiZU9ZWea6t
wqS4ZUB6JhN2WzUWuOSucIJk/1qU4HLfLLVglBy/ObGb9i0JerE+F8+8iNZCzexd8no6nSaB4BdT
TSg69/34cnylxqEbsqMZAaOf816KJd/FPlK/569SIOOZBP2mgxWtMbuVGMDXTM9bgm5/pKI4ynWm
RRx2T5BcwvIG2d4SFYDTmyy0+KK2dlEv18YQk4UesdPZASeXqvSo20QEJUNXFdcBgnda8f7PLUfd
s7mIXpbLdjLD0Td1sGJTXlWM5zsU9XVDjgzCUvD4nqsBBqFecVAWwAmkA7Eau/Nj7R90+Eqsym7H
1UMStW4cQZyQTo0tEa7lewvTawTiZ9YlpG60TRvgePup44D5hyc6SxXsyRSWmOwbMNv95+19lvH0
VT2vlYe3Di/yxriDnVpo/GO+Pe4GHjoe84hdgFWKdYmaFYnAPQFtvc3FKVoadFxWQm+Iwr6In/u/
pDjKdXelYgoxHiSxU7tAT3ID6X2H9yjtt+dv7s9pcFKlDyWx4P8gbMQCKi2knWr3UmuIQm4p8QHs
IDgNBVE31B5xUENfMXhQ+tePYPgw1+wE6iCQ8+dHTBGZX6yLys+vBXkfVGi4AiSCXhVHMh/xo8YF
Xcx+LiUVgNfEs37ZGzyCrGCEkvS1EpzQGYk+lUsZXTQsC5KyPlxQDxAYdDZ5zU85T60bAZRU8gZt
fp23z4EUJvehXGsqG15AcIVWxCIUh8XLr9h4wjdD1XsuF+ddMUzSKb1Aw8lsQcnUiNZkGvqHfUYu
6LZ9wAbj13rPkcE41uO49bRXJ4X6FfPHybBsQO3lTMfWjnbGsJXqn/3oagXeWtXs4WI6whZkgz7F
GVBWaGweplN5jrIXjHehwRNikvMt1A7K574t0zR6BE4KsDQ6xHR1aWdzZRP9wlYsHf/72odnoUOE
GvuOSToRUySp6832G3zallfzlEkTpdFzh10oeY7QFrrC132fb4AzMUoWhfzaoqVToKqJ/TGA5QKJ
Q0KVH0Zcv69W1396oFkyMaYUhf1h8N0Y3CRPgVLHizK1V1N0CeMzwXCtSAxakuhUnip8cqDNZKnL
HKAv84CAtE8xC+tGT3um14bI0QJRNJxxpA9+Cuj2+8pK/DF04gNSHphyUlXm4/Ie2Q1sIF8z3NYF
v2iKkbVIZY1iulYpH1Ete5yR7hUAJjkhlBe4dd3o0eyDhCXgWBIFbnDRFjxXQhACZZCzO9STxgft
29iUUPIDywUj9C3+aFWw39OR51M/3rSjF668aZT+gOkBxvWZ6e7HwBKdbLnq6Mxeb/kiub+8K9Oe
bgaO5O1dONLBM9eLz2BeiHawdQpQJxK56FaObZp7RvfObwzGmfnq3DSUObuWS8lTdvFiNB5zoQCa
RS45WCxxxqzTlQIH96/GBYShiVKyHRCIHSmPDaRC2BN7+SqXpgDgdEHEYro/4fjXJahgosw9qaI+
ZN4uM/dHc1OgdlepeF579AtXPi5tW1VaZ070MK6wK8M+mkelrRhZTuTm2wMEDkO9nV/WDR8ACPWF
7XE2hn74C/iFZ4SqwV+RbgPxF5fKn4jjx5P2c0h6F/+HoHJxCJqCEaHZHPeXL5gzfe5giNKvEgHe
sp9CP9NEvembPyQmi+nHqS3AvPIMvdJYp7GIHeY8ETfiAFBJoLGR4XB4zQ75wtbxYEYv4XcpZpe6
q5+KBA33IX+FOooRMMQo2PCeULafMoyBt3UBun1FPIltu+Cq/IJpljkgq+OqtKXvBeSVWBSLGQjP
IST+psUqkoeuwZpK4BdsF9BMsSb+vY8Kg0EyEnxjhUEkYUhCEC8x34qj6y6YzXuXL1kCsBcPC7jZ
qvxlvBFWb5Ys8zE+9f0dmf2jY+P477FUFT1ctaW66+ejCqV/1iAt0et/I5N6xctppzEi1vchU1Zv
iFq9q9WktfxkckPjdgyGhJylivpwxCmY0XxbHoolfByp9ir6rZpHlgtoecn1iVClfBTcHqEHb8AQ
/853SkLYNFUbwHUSLbR975oH75B8zfnKWDqdfxE1IhCqTFOZQG8pABSn+CWp3vUGqSiTTzAsrggl
vJKYalb80IK8Rl9Z6l8H2qITPbS624fLmeYujMgyWiX/UETV593eSth3nK2MLhViNuV4aRTmF9Qz
BvP95afYZ8wIE7s5+Zw0XOG9fhJ7lxazyM+uxuuLYdRzOsepgA+41ymr2yyL66maQ6bf4o0kDi98
v2IskePJ4gj+/vLwbiKQo4fhx7JpF3V8OdChD2RdhTLtqFE9lNCZXyAQUcPIBkAP5QHDLjkErFbu
jZsdx5tHSHboi4S92rGHn3m/iG30ZgkdQ8E4Ycha7BgU6fQ8SjLZynBRE0Xgg9dXUcBsCOBc5vof
9OupVw9y839VEutOvtGcVsgkJzq1skZFdza6mznz58owZd+zT+PTI0ZfRAqBVqDxatNXXtRPkFGC
+Y5xCufn8mhZ5+DxEaattp1cs0ZTVqoa4DPqRtqQps8pPgaJMurLn0nc91uRnqti2ODgVlwuzhp/
lLUkNzZeRqeZo6uy1JaWmH2OwxFLt8Tw1SuzT+XbTWSI9Oa98RfuJLCnCI1x0+/KUoW6D5+gSmQ0
oom75Fk6CRggpIBxTHupQqB+IK5uB5Cfu9BcNlfQb9cEbJdm1rKZKFNW+m2azr3H4Yd88x0gV5MS
KgOkgJ0+xfLa99CFTajg7h3r+eoPsuB/n4aHhOxVVfQ6/s3/oyFb9MfSDtKxMtM+qdqyqfgMUib6
tiNpAynrZ8yvVVv/XdMMuQLqGMGGGmoyCWsD6CtodjmCwerTpL2HwasIOO1H/yRZYHpV212oyrqD
Es+5g0zrr+J7OmUAlW9YqM3Z3d0obpYXZC5f4FAzrPyLFMdwdQpDcRceVbiCgQYIaFUXada0LPYT
F3u6K9vJQRz2lQi5v/r1nA+x7HjBiQYBeiYdfa24d6tfSUM09f9eMXmsZHkIFuSB63S4jSzCgtnM
tfFJnbcIHNKm9aYtmYoCAaTnU7NttT+tpYOXwUxF0v8THJUKNw1mynesZ5bmOFO+ifIpLO/nhzax
eXn6/59xBjQxj6CTmir+KyNJ2RiB2IZ9fYUsLtQTSP2AS/G4C7u+usgENExX1t71wINevcaK0DWp
uiCD3na7OWg51hE65pNGhB+JTB6aEvi72WT+Pyo7D8eNJT6aqQ3+y+lzoZhcz128fimnCsrswLYE
Pedrt9DQpZtRFihd3tjfFNbU3Nb6IGCuD78ExCaWgtvNfRV83NPLICEgZ+JTWF4rcr09y/Rk7X4i
A/tH2DxZo6MpokPYUTqJLKxXuwmPI7TtDV1/3N5mno5e8tPFuOw5aBRVKnG5qS9P76TVAJT/H9Dr
D17kN+NsBqFGmPLifK4n9P+M9/8IXW1opHUFD1J3qgLZAPMtlg8uxE6GjM05Hrj0TjI5FSD3AyK9
l8zzpNUplH+YCv7v1Rjmyybp6LOeVoKabE2ulpyDg/4FI1+hhATF55VsIxQ6YTtUpORPWNN3Egml
yyxHd35KfkKjU11qbUuuaJVCdzATWASHxFgD/B5Wno4303U0uBU69Gb+HaWyJMoDjEn03gV1OoSv
UULOMybCPgzWp0RQ6zlRmfm39sK9fdQsxUTqH5C/3yORLGhnLsLR72APj+eu9Lqs4X4a1w1+0PKC
M60x9+d00rxKqBJ/8W3LrW39G39fSlSrJEs+sTjDKjfbjv3CyqepNfAjFZIffeIo0cWg8uy1vQFz
xpMpyPesPS5EyEUV2QNIVjhgtProprSwHpSyExqsKnjWaOlGInHqd0tVCzL6H0LyEH4KkbCbDrGZ
m2JyGQSjeCZFjM6rY27+3se8KDbTGlimRzuVL4b7mJ7JSAifc3ocpR+hrn8p7UnlkrHZmnAE2acz
Gr/NRzhWTiZLMJvnsM6fYrvVKIG1eWStQOCRwc3Hb/SmkHx7sn2QU8f0VgcJAkEQJ5a+rd+aVZ4f
WPoCODyBw2b8E2KbjbKf6yPRkglzG/9229xMquGDOKEu8uqLvZxpucia0sNvnkc+uMa4z0goIm3z
yroJjOWntYSpB3l0Ze+ZtFUvWeC2ZiLiklDVJL0anS8/aqQLnQ3200VybRLuKPRH18qP0ffI8OPG
ZudYAOebc/zKB5fQI57ch9tQrGihN8UfcQIOz2PLJ8zbXIsV7OFIDyjpJWVFZuIxClz611d+Ye76
6vjuLwKOlpNLv1CNrqrKSWJMJJ/LHwtJ46ITBsXc7ahAj+VX0ILRrVC3bgwsrrCSVwlNYkJWaH01
4y8oLBFvksSGlu2DKFmToLV/gd6StT24ItEm0gNbPgpGIS8Qw8+1zbWpPCoagFGlwHQNatLUfJQH
KSzhDeJhJV93dS6rNrXnjsm/2tMgMgc+tsrJEgXLYEn2lHU1x41rsJjc0roH/VYjig8nkjDRoEYX
CjsCKhj9Rvj4nZKT2p267xNVSVZw99mQp2Et10aiU4MEyJrUP5EDv4apHELy72yk0edOEu/RqDTg
MM/nXRrvzXnLsZJUlBmQCZ9MD+/Nqa0xi7UpEsUYq/yeGD4Mj2bbw4W8wOjY6wf0DvHmC9VqOUHG
1sVkii2YltpFhpDk5OQk+SlnpbSSlbBvUBUIeyi+8TM0by3Lf7rY5YD1iaRP1A8O15kSHPbYe3h4
2uKtx+SB3e3ygEXhoScqZLube7bnGVQ3xEMdfwE/zVYaTeSynd9VMnLzy8dngdGVXHgJMnGY8qmL
dAnZ+r0A5mrQTH6EZCN61g5fGXLg1qxBhzTeDUjL3XxhagqfXNK6Xb0CQhA4EQNWMwPhEdrMByaS
XL5KRu57fZ0kF6axeAVYaS9xOsUyTiqDFlIJTJC5J83vGKu+myPf/jSggZ3oDwzLlZLBE+buNIme
dzysekwRRG2r7V7mwiBXbybDZN98JAjo+oV1XnjIqobO82hf3jyzXSxsfVhF3gLoNGsDeipqo+4S
yeQMT7ghFu0SGUl+ZtQLy5OIP+sHAlYBFeF7IuyOBMC3iuvmUHjzBQoK9WmO53lvofJiMXPPz4+G
O4bPnYyC25ODWTJdG7ctQYXLlYunPmuzEmXG70k93qmfdEW9Dhw0WZg8KHsvjfxwp+eiKWgFtf9q
ntTTsVcR9uGqWgLpq1oSJ/bppERpNDPORFM0OC/HDtSS8xcIepoXYzEiYsrJ9JdPs5XQVjfjqb7t
I5N0Hi3uLmGoCi3ffpnGfSjfDmMBKwfvJaBiZHAJM+QEc7gx4/GgNZD0ijMi7Rbmz6htcdEUmz3M
ol5f/VsqCkliZjRSEPOPcTvDtndJT5Sr+eYcQmavAk1mxBZdF9cxCUoRyDum6Qc06YpzidnKLXVJ
RoeLXNqxAPazfTpqDxk/7QUoeAoE+PsOPlW1QusQQuDmwf/CpkSc14oIn62ZtM9CiDPNxR1uayob
2Lwm2A+8aA1vJj4Dc0Ejf4ySGGCSRBa3kkCby1iK218tGgitj5bSVDKVB/Lvs4Ov3ybgA6JwX3Ar
CEMbPaHUSV+oAnPiJHKM8CVpXiV+Xe0dd5+wWKEk9MeLUte7JhzW/epovBApeF1D0hQTxo7tweEo
BtslyFmIigd+lnWynw38t6AxbpMAJSostdAFpUfoP/cs0QJcrsXIqXnzCobROMZIDpPo6G5wXj82
BMdKMrJn+rXAsVNbna8Y6B3iahBr0dHdJ4GAi3L1ilXhEDTLz6kx5DmcoWyB6V3ir2ndoKpEovhQ
S7Yh48nYhrCN8W911YSzavPHBBx4dpuGY1Y3Jw6xrZRweqot2v2+TCYwR8xisIK/8WoaI9db71+a
8PlUGXh5D7A8RpFrqsXu9+fpxrDmtZyX1l+ByeVJgi7GJcGbrtUoxcza5BBRI/6GPS3fJrI9Wody
q2MCj3iEdSispVz608Z4lrS6Jv0kzWVB0wlXWgzOK8SoIlSJbiV0DBUR8y+48kQwsbeMl0WTjt3q
fMdS10/PIP5HGMwp1BQ/fxhDgUkAbN2Xc5YcHE7xshNloxdSTfYVP7ownP64xzu0+V/dYiCcsK5Q
Pw7VFYMuIwg36usqQvgQ4C/6tsHjI5cvyNqgHbS9OCx1TXfi9h60Zek8VaeyHp3CRDLbl4s58mV0
pSpyxm+l2naFK8wh/r+iaBuZKltQ5LdFl/O5IrUQvaz7UbXQFz8vGyNiFrnCBODmLfrkVLXH754r
EmOVwGLOCwVt9UWh4H8riZnV7x099wSy2dQshGDFUgA6H6mgVuD3mMCmeK4RWewpPvuQFiaHkTGf
cbdjQTHhVrb3KUN20GubNPGKkt6sW7FUd/eM0yOUIX4FXhETom8tn6ajMkhAqJKtY5qz97eVTph7
0pRZHb6bhGyKDIq37g/qnl3iZw9N+sD6t0fHhJnEkLNR1rb7Z7fWhCOa2tXc6jW6PJKepacItJNO
ywATtKNZGF3xx2hrBymssUQs0zlvqPATD7wNdCZrkn9lvei89ELkEJ1D88QBuHGXD2DereeDz6M6
zw9cIX1UybUJ4FRIzBbLH3mHn20qJqVnEn/ElzyjjE9KNWFcYqv9VMKJE0yczmmN3LRpfpETC4f/
5Ps1Ql8K8W07Z+cZATrSQYPVouUjFdowRuw0SK2MCV6CJZen0hIbXdB+jvPkC3WdBDlyX1N/XdMi
iaHYCiL7+/eQiO7ZA8XqviaZX2Q3SmVlm+zVX/i1HNpOeewnhB+NvyvDaftPEKk2E1+/HtkDsm6K
lG7AhundeNzcMqkxMqFG/5rAk+a2YPHtnT98cKYXWE1WUNsuZwlQxEwb2gwI+QJXBOH/w6spEf75
sJErm23P/0WPbmA/PI0xrBB8aIvgJrA8RjMTDA++TvgHjzlR+0B2D8qoPND4G9SJRrAKYqZuHDVa
aQ2iNuDIvympPdBPtjx1+uBL3/ehTcbmdmF11810mSYRmvAiSvv8Ea8Y+wXEGxaxubzAInxMuyzg
DRijHForPbDICEXP+QPcsAOCv5NkkZQmgUYHBng3qh65EHxcBQm/ciJbsOAEIEhjNGth/VKSwTaQ
PVi84xhBYqhnzz5ELJxFUVvlJqGdEU9yz5BZJxAbn73yvV4ZE7cXg2yNK7a3N2oOop0uaPhhelAS
NbnxThmn3yR4Id6Wj931D1WCOBBB4mQPNQQUIFEZcaGVuuMJdNcOYHUsdllJ405yDpuqnxCZWJeG
tZe8CPk2NFDBjGBdX34E1jsIzoTLHMcHPCkyTBF7hJkCxi6NzYmAdFnfYTI5V7xoueZ3fEnQPjXr
kgZ8rPB3jheIlvBybze1jS/hENjBhl/tO1jBI8wjRRLN1Ez1EzqTrOq1K6RckepcOkASPyOaazLt
yQ66mV164eeHxCnTDGiYEpnW110CH2BgdiMWgbGX840pevhGYEaK/Dh/+FvyGKtPXeeVjxsuD/2F
WUwQpwuYnSqReUF8/uBGmkjkr5hvqiOANXd8fD+Zvn29IAPltUeEXFkac7J1DHc1eLc2J81arBnz
HajdYEwxTqsDoye6pIM+aIDmNGZWkNVGlJxujMjO/aeE2vLlBey5Doy2hp/mJUlbHNWnpIipXMu4
oLD85zEgwlpftPsePfPDjNpGbZ2jvJvKShcMB2zQCaoSlkhBbiTC0paDIIVqHFZCduYK+q4dBls9
/cewVl8+FYq9XE4E3p8WWuaL2oDvmMpe1tmx1aSUhAYDtJXXBqgxJS4z1kV0GBjfQYmq0M3ZwRU9
Zh+po5oVBcCWm4Ropda8Kz/Egw0SjrK841aJIWebTPNGYwEMzYOcPZSMCV6Jemi26nOxxfCbeUbS
wVAhsLKVyKU210cDax/k6ZGmfqeLzy784CXRpruOdKy6tz1llmdUoORh/E4C1LiEQO6U3ZlNTWUk
PAbZzyduIYe22SoCVByUJw+GPhXgPEa0G//od5jysklAQ/L0qsOGiPP/MRmDVlDfFO7von067tgT
okwIs0mYsz6mtJ7dExPWxI/TbcdB85Xx/9D4jNXqltA/l4s4tcv0GxbdzDB8Q1Re/5if/xe7gK3B
zA7M6aUJ56Riqsm4S/65A3dLKBhnS2F8g3WemBPchPKGvdz+f2LqN0ouEa1MGd9sabBgdUJm3lZK
K9cz/IMy1xe7rMQPX3dZogr1nmra8ti7ZiZOpoaPTdDomW0XeaGRNoj0Cd4t5qx8VJMeYJB3cc6h
FcCvVfZL8wz3cmaRm0YQ/N/t/ehD9Jv16QTQDPXvxpyU/YzXpaJrJ0+VRY0dB+XsDjN1JlPUr519
mcGCR7aVJY4BuGwhNUme77POV83VQcus8nmSS0uIxj9QysKSQMaaeuSVrYDY3SeS/lUaq0LmM2Y3
uLrswAmkpaO7OOtEeIH9Mlu+EPRMN3BjOCasy5KXU0Iuk5vmYlBveKHJT11VfX7/sYsLMgnCcHXK
nW9iSIx0YajifWCK3qmwV3Oh/nrf7bcmFdgzhTitcPvFVCXK2gOJtpKq6u0sx54jMQg9MAilLW+0
4C5ZkuYBsR/t2mjV9k1/W5ytjZVXNJ93+wdCuNdc30kVR56Auz5F0zZmmXmNqKOfoKSUxZGIygcd
kWP5fdsrsweKS8Xpq8kfaIQAakJd7fcTAc8jWhGis76bpcyFL/XOZ+dtvuKQvQFDCumvO9GlmWtc
B8vsXDtLwipSxvyYU8YqBMt1tVTa2LdPdQ0QyaXg7CiFYVPV82mDKRKCkH4NALXRzWcd4PgUF2rW
3QjRyu6qvji9VseLJbGWXlM+dyvnjYNnY6NI2EylB+yLLR/ws12CxSchBUQRHXFCJYMF8v/PoYSo
2YfwjhwSAM4UTMk3o+/T7Q7/cKz8DJweNgxPMxjO1Hd9HrVGOu9vIedBRtYCz47KueSEsFlDX1w+
2iCQjbZZE5bCTv/gBn1vAk9lg/AeklyXHMqDCcNY5kvuheve63TThEgdkiulkR74oKFvIYlraILA
z7UR3YBlcLuzBIojSnH8/xOz734oGAPI20jRTyRX7TeE2Bp7XIn747AgAbgMpVnTmmPaIM+pzSd6
39tePuHhq6oeFaR0b9JLWUeh+LdsVs5hPjqjASCj9b0iJoj4wDFcGncbmzQxky/XChix3zKM4Y9P
AEogiNiFRpKL4MjRK99PzQVPf930YDju4FwOVuIN2IQ70cRm3169nndyByi+ZBxWk3PxndNWbb9Z
VWj8gYo3x21lDwoKmCGQf/DqKyQMAyf73e11Q8YUo34vA89/iHVqP3kKLvGaA9LzIv/OCG+Zz66M
Qd/5gD1QaRIMgJlOKzLyacTi9tPXhPYci+ILtBi135H+VAkFUjOgHPJs3JFbCXKG5cm0b89szIm3
QtU1dXDNnRAKvRCxuItYpbMIWQJN3VHw1dvU92krvUc/2fwvjHIZ337S1ukaQXqJxFAtoaLdiGT1
CV5z73cS8DgKcu8PslKfz2A7yMF5paY9TmiLeo/v1i4/RQQ315giJX0MspstiX8wymUb/zsJ9GWR
NmoEU0Htf73zUDXtnBTnUG/PgUGmKiA8aF42tnB+2YEck2nANP7UHvIq74BjLEicDOEbWF28/Xrq
oJ/+SzHFcr/Zspq0Wrh0OSQtI4/kxLcchuVPQzoGjLiyVfXi6lb2+NgSFdNzNzMr/r9JH6HPdQ3h
45cEBfVBZu3vDo34VU3b0FIuPUx6GWdn+ySw4BMAAxzeQjT1s2F2A2S05ymEJ/mB3SuvQ/LjMRIU
DNaCC5raCZpq5p85lyNQsMwUJR8CswOTDXIamf7ohdErYx54iP7jbZuS6uIpg3v/OPgkP9BPI7vc
s4fNw4fxY/LkGQyk8Hh6/5UmhcyvRjgFxsWHo15g3+5ZfSzzsxnWXO7coUapcdgguVUDp6rBIGMG
9CAaUjC8GE/J9eeAnyV+jFnimdCGs1SEwFIRGsA72EKwKk5KFimI7Ho+fjVSzPEWNmRNaTyGiNEA
qYHI0pAW/EpnABhRwIB7AVXMzSzJEdsJUe4Q9jSsS4ETq1+kCH3Na096sPADVe9lg0KiuriPGkSY
yI5y7hcLCT3XBH0B5oyk3nGxXYRuiOBgHO/Zg4etGBFJy6SbpppgCYEktYb45AwELijLWl1TlDrL
GzoNsM0vSNy3GL4crIq65fHy8e14kHui+llsfKcjfuZdoOwo/b2TDw2K6Dac7Uapxyp1zFefWfjG
2cjYydDQcG8QrV4ylkKjpZhucFRhY3fHEmr4HNhtF1GK+nHwQ3nxNUvNkL2yl2K4kIniya0TUnKj
Iwd3QnnK2cHaMpPoSSsN4V3lhJ/2vfFHgTDWWJEH5yFov/GIujSU5T1CGUm4HurLRAEQoGdRew2t
EWR3GfmUnZoAnwkQ9rue8Ay0WN3h3h+itbQUNH/lGOlcxYVlpDW1fTVsKocRZhE7/jnlRQlyz9lb
wxUYZSm7H3CpkmKsPqGRd7nK1cbfL/1CIj+XR1KTneLf6SwB2azHqCvk+CgkddZAhhP9utC8Zb+Q
n0Y91CnWtSD/KT3Pjp5Ezk01TwJHTt5G6v4p41CVq1JUtREtnGrFzMLVBVjINpKYrHWiL83rVZ01
h0REfcYyzkqlHKMI4UzlwJeJrxhkSgFkyU62d5km0ytSbbOUOkDvTQGpioCKU6fscHwyP7o8RVVu
OUn4XcjhrS0vCUUALVYU0vsLRogvQsl9RYiT1AGRkFMaJSD5v5Ym4NFQ/lr1MSp5KPRc/adEG2D5
6y2EI7WoqzTiffk/aSN6kFdP4qs9IqNibfk+AVJzaSxknNKwf4SCoLHXcwern/zwyoZ3SSzxChQ+
pCVqY3itLIJ6CByzE1guEYpO2fvTn7MsbU9HfxQWxzgt2Nfye8FDFdlaVLek7Z6K7zjjUPhQDTJ8
fbn3UcjX2dwZmKCPSNi9Lg2xAzNBwFSEK3hNEtmBA5UKIWhaly2t1vQqrtQw0r5nmpNHV1UQw0uu
1ECfg7g0qhHN7rRu5fQkOaeYuV8He5p8nXwzE4g/frHspvUzvQUDxneBIWHb1LpdAby2T5d1peSb
Pv1iPK60R3ObsiAD1Lzdwfk3QhXJl5uGebaTLLJ+cPZIPKXUNugk3nOXnjXR1WKYVfPO+mK4vH2s
NanC9jtBCojUOnyUj+TLJkAMBWhOTfNMn1/51L2kQuYmABUKtmarobRTtEqlxQaxtR8ArBy+YXdr
dQhDInXS2ib+qbK/45cr576wE5bOhuxHNjU/ZtzdlYfCE6i1dRakzXFuz99qhec9+Nisds+TSLQb
M5Sr94c/r6onJZqKhAHr/r9UPAP3RIhmPwC/Q7O3cwl0MTt69zcwmHhZRI7dolYdTAhYghDXC59H
maRIEYavIdtD7mMpHkIvy5/X3T6oWju8BRUUqkIUGQ8Y5otHv3376MAUNQa0Z+AUo39KvyTbuenm
703uS+B2u0vpRNmsOFVMKcQVBPzDFH2AZXJiU60hRwnuCkaHcwkQTi57+1F0L3o4xdNlzyz34qKj
zTC7GmpIUeMpHO63xq0SwJKdszY+ZOWkNhW8LrwHNUzup+jt/Zi2xEVQnB1s/JHMQf9AtdCDWi3W
NjYDaZsrEcFe394QCJHkjLZ9e5bS2NaelKmhU1CRt9sEyqHzCxe30PIF1oS3YQ0q6/8ccx9XvXiO
DSRxZW/NCpibj6eAy7/bnfDVxXh93FlBTW9G/6gQ17YxyESv7vsG8odkzsNa2VgOiEeGXGnEl7yZ
arvpfqrPRrCRzZDFk9NoVNwUr6JN3zxFux+BIR2RVMW+kKDVk4+9+uOyzWGn6EXX3BD8yirvQsFb
2flNWF9wQgKFFSjzkVwZXiey+rPBpoZwSm9RuYZK1YK0bXoayB96WQHEvh/7kMB31lzqR2zlc9QQ
G1ya01zirO0FGHZszF7mqqu16Wjpv8EGaHzqYAko+CwYKi354spY2Yf0W9jzXVVvgXH8YCij78ch
3oryWoJIH63yq8WkuCwKMUlQjtUZ+PFbd/GwK3KNRK63ZVoODWLt3/+/UJZ1gH4waU1ee1tTrKkX
CWqBiOtH66V1kXTNMjU/1UAwWrMS8X+glPRKi1jnppHnKXZA9+iQm4UUKyEw8icOWyMk4ou8mNRw
kds93+mT14evVOUpmFN+a54rX+KPrZNqbiU5V2XiWC48SqwOPZXfl1e1FYYQ63P/rCr3F5vEZ/iV
irxxTv8t6aTIHYw9e8nWXTa0Kyje43SwstD13DPf9jQGKEEI3vhEPWCEvN5q6pn22S5igdAX5l3u
lelhPBqyZClTsry6moRoooqpPUWCmh20jyJDEhIYZReDrYkWxrETRhf+FmIk+LkDLoO5wSBIGv4g
iJ0nKkcbQhoJFD3f208lcSCZCFlhueilcWfjpCKHImy/qkC24mGxTjVO12NRsFImcfV5vF63mz6T
4HEZrZgepCfFgQaz+9PkL92vrGGqraVb/5fd4+q3vyCqwW2oZtChRy1X9eNPyRf0PUidI3kP1VDz
eoQet8ij7AVuboGiOvNvKr/hGOi10f7TewZKYR9crqhga82qRuTLxFq3PGD2zyf6C792QREQ6D4z
Men4+dkK1vAYblQ8aanUY/LDuyWySuvDTJM1cGSZPQ9DxXjwBbV3Gw6K9sjnI+KUGh4G1siAiZOi
CiYPSCMOfM70bSVV1AED3iw28V7Rv/1rmt3zKC6LlUQhUPRYvvbDnD3LjaL6FBruHkFytQ5ZB/1Y
ilRquSF48AdFqZC51BGotaOesctvg8V72gBY9mn+IVDJXZaTtzTINTpM+Ydr2g6Tx2bzk/fRpx5f
TTpugAP6v6dH1N14oZlj86nLNb60ECalEhuW8iwT+necxXisDuySQlBdJfXApkjW0aelZYC5EkNi
5XWwdyRC9HuYrNqNlU6gzulunfW3czrGTobD8MhAGBTI2t7hySS1o3LR8dcAy17D2sfW6He0zRXU
MwpiWd0BsJklPtWg/FwBmWbPDBIHGjlPMCxbnIgv5+Z7TTRcmJnDoCpJjq5/GgH+Fc032pzFxR8H
4Jk0OvBxL4sc24Hzc0Ev12lLoiPQgFiYn09WLC5kUmHqgVFAbjmEQKKiB0q/EYhVEA9guunJLyBZ
Xt3ZhTWOIKHiwZsmsDRX8XaOyeXj74OduxT9vMYPJ2LRKODBdN3Gf35aFf2OTKA9FvJDcAKsIdMv
5eynJfd7yWnJfMiiTKavH9GBVYVnFDpxO9g5rMsCHBEc2hgLR4+9wXG+kJZ/z/dAA9f0n0B22xKp
RweqL+LmO0OJT9DL6+swpUjduh9OYkcJ8XOxB8tNHhRUlmPOXeC6kTFJ1Rq03Te7T4leHMDGq+Z4
EgsfVhriYPhWiaAUN0w92isLTkeSYfvbK575WD/zoHKeswIINLnvXzyF0EbsMXwQIRZ7EUaAU7XB
EINfPc0R78eC3H0VN98PRJtGkeaIeWplvPPaNnyA4OQctHI12UFLdeCEP61CtkcEA/niqmnScgaw
xl+gly2NEhrLk/xQxQo2M+IQUPN4XafbZGTprquKwap4bGLQswPVlQSb1HT71ZPlkFcrEJiQjVi3
gRFrgIsLKHX4HHKoyTavTceJXE+I+8Ka8pSOOcIc10hBCcKXtVClGkespZnEi2BLeMZbIaHLF7Ck
wTY0a0oTOHtVC99JQoaRp77crevPBjzcfakB56PscttHVDhiJEMD49kEbGvwkXvgEVf+b74k1+tK
lBdoVMPvHvJygHKTp8C7Tok6pSAfsPoiRQ6yeC8qRdzkHrGhpYn22/ZwIJO4LCDIMehn7hOwXBVc
6I3rc2fROVALcF38TuPkNZto/uYoh7o6XAjlbgPG2TwvQ+YtRnCwQIhcskYgLnN6CeUUoAfwN5Ve
sCI8POhDXuYyUvSSe7a5UM9eMzPFCaZbm0mZ9Rh5bLGmP5Wvhq39MzXDTgCkNKfdLbQ21ce0fW3v
8i/aK2fiukgCVyA5ile4k0lRQbVz33jQfZo8uYFUKcaeOeaXWtm0NBuH0AhfGU0fN8VqQ0v3INy9
5ROX1lZ1Qjjlzfb9L8hnaKdgv2bLjAjoAeOf2GiWj+zDad8BWk0HHYR9BfBoYxBLaYkjq8VtfTTx
nwAE9CsP4UU3JIjFVcpfOUeQqY2AGKWtWKpVT53If5KUCnU+2zmSqKx3Iy0lS35MPwJBxQLjqsX9
uncIwc6cmumcIlIj8KyQL/htMgspz2B07ueeI56iqex589nP03rUZLRbvzH+yJLfC9CAlwf07Pss
c5eJf6CjXahStATd1IzTsAEzKFdOE5n5KHTwnwyA32pZf4g3U2pzREo+Zw1mnGwYO735k2bxCJNn
Tz7A2TdqEZxtjuyMOnUR9JKn8a9Mt+2/n6i21lOp6i5xL0EXycUwYByRXSkCfYpmLbjmG9zPkjDH
fYH768j23AEN+1hj5YW0NlebdKmCzB0mTy4YT8MAD7HiUltJwZHcbj64cViqmqDZIDkjYzqJysoI
R5bV3pjiZdq71m01+faOunyeS466HE3Cn27EiQrfiOjCuKPC/CuqG/SrnFAw2/zOx+Q1MdpiIbcA
N4o1h1DAULi9i0Rxuv9dplbLK1XZAFud1EAREeUD3fux+QzJhkp0knmN8UStFFxCfWpi+MzV+0Jk
uZinM6ieH0OMPyM4SgUxQEy3Xmsy2QA972MjeLOl4qw338g0mb0eHoVKuVIP57WLZN0gxjDZYReG
zFyfJV1a4pudylgxylvrBdH+jrRhirWVB/4vQKj2UoZqnfucsKp40iikmdFqU2fJ6R/kPqDudpNM
120EXomTBVFzWAJbpiSBd67bGDibv8Qi6koYKNefFJEunVraVbcqLRolkv2qJlpJLvJFrVWkVVA/
WgiNSJNXU43O272aZON6DtqGc0SuolXUpz9X5TRoScy0ZOr/HNiMgGQqsY1zVatgeS8JhYCWYaR8
rNl7rPNpHxi2zpu7h047M7zPliyFfCg0trFwlqbYhQAHu5EZyn7pZGDXRV0jAuLhzGsl+1YHs5iC
HtYxYUThyihmGRpKNnhnONxR7LEKR2ykfv028iJq5tykaDg53/Y5E5XfUgOq992EA9CsBRg8DXPd
//sgXqjYSEgpLexJM9bR8irEUBlHsbZZAH0k+zx/2xAw1twnaL/gaLhRyMufOHiP3Mjf4QA6Xuza
v9JH+oqS3BhRqNAlgmagAEhx5YFtG5qHTtlqkEsM2K2BHjCycjOlD2GnEKfeUEM9eUH6TuWTOLIB
BUnszcQLWYAwAP4Z60d90hXloRYmKgngwwiw7hUpBeID00o5vDwt56uA3gKlIt/2wL7uQQERCBDG
9kma77NZVuMpoJVuxuGIKhhZ2Cnu5aDlJACA09Mq9mJp/klPxe5O3tOc4m30nlmiXZ16Xdu+IxKZ
HWf3/3ukzE4P0wXGFp088os3A8G/vaCMJIkVd1PiqZygfU/Jx2dsQ+4yq1FWl1zetzcsF3g+XB1w
6iRUIU8JMr8cteBmsbppIc+t9bTBG29shZ8p9xq1Xr1QbdND5ag3fISYZMULEEJCIi1+2XCbyQxL
8XQAPT6g21Opv7UfBgTKQUo1jx5EmJDUJCfMrcZJgN3kzK9REUbzubo10b/PWQY43nZnoj+QSqu1
7gcQsJzM1fU83teRjRm4qlfdT5Ia1wayUahJuvTJ4PitAZ9oiXQ+HbNhv2n/Tt2y0ISkfxzJHF9W
OcqJe0bkwHqHu6XcHLArlNR68W3VFUk1cMt+hbW5cu9nTAhBkIQBGU8p08dNXGn5cI3n0JPcqwtI
RYs+RLs0DRpPlCiTL/rWfQfJ/JSAMg25T97gZ2eFjOfgS9rpZqDDstNTlN4r5QGT0evxDM60bTx+
GLDBP4PBY5qrn0F2OKGDYFOZwKbmjAb+G6ETH4K7/O27nP69HiwpkJobnYkhp36L1awCegO2psP+
2qvN8KioXz0RRv2cd9l7cZkFRW8vbcKDPBrmsveosjVYVy1zUgTKG/XGx4DAHdS52cHt0g7CfvAH
nqEWq32An465eQyC6FUcHSc75D3fzHvVHcWk+iP/KTgQghd8WIl3oyJ3+NpAL4Q6RTtyY4+BOR/w
t155a7uF85R+zpHyyHP7zostrNi4cbnSDWGtcM/IUPrwbtTP1RPyqnWBAD62pZqTIteHTR6UXJap
Wa6i5LGmwnABxliP3jK5a0Ri1BSZ3zrMyP8QZhA7JDK8UOFXvk5Ta0WaVSmI/tUZB7wkYe0XJhdh
1lrbSyDo/lOkMOJeUrOarxUnE6Ygk4Vuq+/0jtUHjLk94XQh83rvdGeRH1Re94uWz4pqXKW/38eo
tr4KeRv0yR2e5AUsY3rM0PmJtyOLU/gzdfXJ6tMBMpU4avNoWf8E/YynKRtZ/YRMa7b0jcpnsrBg
Md4/oo7HY7ec4yO7wX84TJvVFylcnT3gJ7oywnSNbba2/RwLj2l31LRRAl73nZF8JT0b1UU5xrxj
xPo7aA6tNBaFmw6lFMoIVMJlFJ+FLACiX53aEpGFjQ8OivIET99NmqIA8QWK27wH1NOpqNkdy2dZ
No48a3RIJCKqyNm7pc9HPLK98OsIqjD4KYLmAy2zC/6+xKWPgFcVpyDUDe8W3EzO0+sVRZlXoBkC
T7dvXaHZNba/K3M9UzHX6539G8eqyAwUi2Eenk5dzffzV7tYD+PXurdwWxRsnjupRJ4+bMIC8XSU
tKZNFLV8TcloOHl50CaHWtX2cbbYn7geRFmkRWsZBB0fdkEsD3oIbt+KqNrLTNzQJKuN8P/3a6Nh
ahi0PKS/Yj9yUSQstba5gAsKW4fYPXLEWWme/cV2nfqPdTvnu0cfw1lRwDtlhb7Z+tEg+SYKTwT6
BxSA6Uv9bdAEVldcWwsnDtuyzYT5vLeMOYNZVqFScKctNVL/iqxQC+s3M2SVoPWpW9siIfYGXVfM
py5R5A2UvDYkUyFcgqSI/55z54r/nloiPowlAR8AwND2UpiQ51zUIPzo3mIqPEy8GQliN0Rw2vFg
EALFDoIhpA2/g4NPWGRZ21LKUNC97wYjCwhFSutJDAwXHDWT3ALUpZCiEDpxeIUdYcbsxdZskCao
iEZTI/M1JnyLnifSj4Sh8nQ1BOXPbjQvgpCp9sfEotQPQ3KLBMS0XbEzafDKU4pY1vq3UzxCmeTX
b8TdBjdYKojdzWX1TvWl/myEE8wRqa0olctXDrjrDwMs3LYvQDrtUEBsAzv2rFZXyrcsD3BoV7lO
inSXIK+/MvQSpsktgRvRddGmOqGq9GFOTUPvAxcXaJOE2qEXCd+xlp8R7lmrFC/ibzYv9XsTD47n
mCBPd5FqRlHEdCwnpLEP5J57LMNU4ROI88GP4v9Cyh7BCzNcTnT17R0kFwFBDChrVdnygNVnmmOW
No1pGQXTN7KRfneRVo0zvJ/K0aLV5y2CG+bO7KTepkH5fep6qmml0t1Q7CVTmmHMFQz8JTEYTW6+
JtUekgoawuerVHICZgNhhxC+emiyOQVFjTjFInNzcgT6fHNq71qqpexSpzGSlaRjnxx/fhco1o/3
brmIplY3TrhU0X5jkVbLVXheok4sQSLmEXdCPIn5lvg/UrA1pJamsu10Tnj/WfgS6W8rHOBl2WkW
wEQYEq3cAzvuzCkKZ4/sNPZMk2CAO3jAUYGYLOWEpM10ZXxfvyx/vyZXZ5h1VJyuf90KGxmnPhdi
RedokqOXxrpaSiW1Lie75+Zy76YtpPodN3a4BYsXHqRKUN75PIzPwpvSvXQE6b36vqTDPP3qNoaq
SdRWBdeYHBwYG0qdNwQQuNJO093f0pyB2R0iy8WSEhiu6aDVCtvOoM9r1FkXkfbHiy/0kBVmnkMa
i5YRR4/1erO5YkKrE9/5z7iuMHABozjFlir2hgbxwiSEt/omXk6eRHtfD2fg+eY/zL8+f/DL3Nk2
JZErkNRH3Bvtjk9N4h/rJaqvYSmmt0BT7nUE07GQz30xdP2bI79Vsv1wMcfoCo2JszRSKGb/bI6p
pjKLgCM8cx3+y4NWAX4zrb+Eavd8J7q7aDpF9TW7Fp/3N0Q6iiSkdjjaBUfBT5lvzZkknStIG98J
rC5R/jShLLfiR/mvuWv/l/stVamSbXXG80fAnnyq9nyJXjngPTgT1sRi3kh/7kTbhJQe0PVx5tPE
wU/DqIR3tNpph0bgBWQmRlO7Bp96J9F+RjM2DYX+vItmdUbcKO/ICLT0T9c2yb0mkSHvTxrjEjuJ
/HP/aVKA3NqX/W42senwscCJgCLrjjwTyIBKlrjjwblYZ/1l3qFZ/2MWMRVrAk/ggD2aGAyv6I6B
2Cspeg9bsspm8H1pqBGKGYZodDqGADJoUbnlYlYlC1kaA/4lYVo3rYF2gmZj80oYOf7I6TKWpUyk
3DpQjjKxmYw5CqZXJrlKXyFpUIXymrOHJMPTV7fEXLgqIWyyKkSslX9x1sDLfgwUNYtRc5zvgC6B
l1RE2z7oP4seqEkg8FtmhpVEEwLLFTPlKgzapIHYuEyF3oYYi4SPx0hqQsrZhsTnJt+dJ+hTDvo/
RkHuzjVarcjNjsfeC2f74bqUlHKJ3F9YghHR+NtKkql6QwBJxnUNTocNjz0hh8GDwL0s3H7noYFm
Z7BHBduSRtxZBt0PdrIePRkMnLfKyPyla1WvmSiOLHZcnsHFyEZT+sap8EwNkLn4MH+XJ1oyfThB
IbI1HwgKU0gQ/zIurQ5XP6HcoLcHkINTlRIhsZkMsMKpc5AsKGovw9GFrcv8r8oxZD9yHehhFaY2
Cqd1a+oixbNrtQuKjfIe44W11yIk3FpcF1EpJ+x/W5XIN29sIjchEFEHTpA6UCOhLWMDTnfpcayy
sqMftbv68pjVJ8CGUvbwjT4x46tuot8dZJrcN9dP0AQ5ueTH1irlENbmIH5iFdrDyTID1rG1O/M+
L3Q+wTmKgKe+O9taevb06QIIU+CJb9PyDarH9r3VU27XSVa7MwVmGocDIFlqEEZkMX+n25HSxtUh
6LAVyb3q+9T9gPe6QW0kYu1CkN27BVMBskA+y6m1mKp9A5yLU8w0FzQdWXeCCJ7m7bHAuIFMgSlF
XMkpvVjwb9lei1CrTlH5SKw9SL8DzrVvYkjSU4OaRze2548DexEDdiWJ8fhLz150YnW+kbkk58en
SvoOJ9fzw3gzHjsJCsUimHH0RwJFmYjvoYHOjspUKE4oBpjDAw4ceZU9XQSgpOV72aNfPKBvd36W
cfBxLd29qI8OTkHJ4fjluIk+RLQsQzBVj6KohT17Xe0p4k7AnpKA8TMWE7XPOMJdnVkRdl0LGwbA
hAbz2bONaYVHVqumzNBwLhMld6ZNwmyGAkmsfM0Y5gUJqbcMo/xZK3W2pk0ewBymAJYcRhmtbR80
c/RAtwHJGMZSxqSSys2ONJ/FwQZQcnMjYNLsdyL1ggACjM24O93c12DsugnvzoY9aX/1aP2cRmv9
kYOSTXQlfzfkokYK9FqPRCDqXP5yEuJ1a9YmyuXhP+3ssSwiUzV/c8iv1gsRkT8CjLdWa7aah8QE
U7A1eI3dygyJlqRE9o8PyCiuTY04mlmo48ApAAR9Bc91hLXHpHBi2s/LroADj/eGKU4T3UFC9Rva
D2LBbR/0VkcxmBKoaRzS/BhoAhj2V1oVvPjzm+Z8Nnfjj2nVwUBU3uWA9f1IAg8F0iR41dMac+lF
TU40ORQRvlGZ501I/nLPvD1IOq59xx9PXoDkQyAN3aSMLQYPPDVEkLwJtfV9W6xT4U+SbAiCrwzh
S6BCC9b+4+dIYNTc99Pj4SSt+BMcIPVsee44GRJLuNkYGJqBNWzNF5Y+rz8MPTeUT3fxKpaNMiwP
WGUHasyLfiQCpy4D06dfED2VCANw4jpTgU0DRJzP2UyaA1NLU1uvH6cNS03P0yM8fALdpbjWt9xL
kd5tbAKTV28xeL4rTjsOv02nitUn1U5KocZSwWZm8zTgrdK/W3MQw4++3CuFPXIhmu4WTDHMqY9W
tLfMYTO9RcQm321KKu7SfqpJ5uUkgb8jenRZj0aR1/4h1F6bVr1spzM4EKKYXjwccA357YLANR+z
7J08PbuBzJW9xe8TJ1NoGamR/w0P3SjoKDTbTnoVywnycZfu9Ho1hiZN9nfWpX3wT6bfUP1uxCpD
sU4Y4GeJVlqeFwNUtDG7ywmwmEvqvIHXoRr/SR0wlz2BhuOiwflyw08tOujjqc/VSaIarKFH6G/C
wD1+fOHk7XmPbTF4pUNTap77RggwQpbvFrBmmy6lQD/i6TDMF9G3OSVQtDyDlPmIcEOQUvR0DaR0
2oCpX9oSjDRnLFj+3oziLRwKYWyBWK0K5pKYlmm62c4xBzAEQgA1KioOZBvC6lGXX2WE+qfrPKND
V2Z5KlaoBoUYETvBzzDDrNWlkYB1CQvaEvO/Fg/Qhh13yLwUN3ADJ0JhbLa/cZyaRNJbQxpHbqGZ
Wu4N3/Yx3wC6r/M8NWZoLE2+D9je8+uct2BbY+1LKiBaoN36ajJJ8QHxl0U1m/w9TTCUZ3Cv5CGD
jLnxjceMmsCUU8lp1E2wNWlV8xfA2a0aiIStnbN7IEi4KEowlnxSL11oXZRXrR4T8SK7+HgX8wey
iYwVNwIlOt7/l18DjIAfjLotSt6cfSgVq/vaqyl+yPprMJprdnp48qcKwZ/n1IHs6shGL3QUmlcb
s+8djEa/I5yGmgJNrHDw+5rX8vqYJL1NVUHQXQ8Utr9EVMpIFpsm8kwT5UZ4lYuEEUKqaPnACsuN
VyIk0V9dvxyBxQzDsMyZ9wy0O73KBeoqYQhVwo5dgLspCi/lSi0Ie1Y7pYxnuNN2Zx3hwNq2WfIG
+C/+ZZd9L+JovCANQiaXecvfCK9sE+GgWV0QB4xvfo9pDmMVKNuM5/DuzmOmXhDk5aVKb0J1vAyt
3BsEPHi1jezTDhr9joW7dKKA1DiggO1uaxoJS9RwvdNJNZOcQa18ZB6P9DtkoHv8XKL9WKdnxXm/
O8dIkrVSMJMthBTE3adjcOQ0bJ24HEpYZ/wCalj5E4q7gO9oUdWICYjb7axMxiN2wkqW+WxtDNja
B1BRb6kASRCis6N7ZDsJR8LGGf9s2o4XFiinljeKjtPFlhuY+eEOp6yXDUK5O6erJXzKivBSfk4L
8NdA64J9mPLKMffqUDiFlL8upGHE6G+ymrFkv+iA7fSGWkljlBs65GA4d3Fs0LaNGLIa5ltWWwe1
d5ITnlj5Is7zK/H1LpUR/t0m8XS0AsMrzkNgcxPVDNqWsCXsc+JE6ZcpBdOzm844YjHSUFKxLBob
5tZ0MXO09mV68czx26I/6jQlS+M1eUG6LYB6O0mHRwLHrclX88Dso9lzbrcQpkzbUQk4AjAuxuqJ
Ai8grQLHl2OhesMy0EzMViUIRweWi3UvxvAE2TuzVs4H5d/y9FyPXHt6O1g+V2NtGNREwj+0S/+i
D4Wg0qqyiCQN7qdTF27QM2iu5kTPlscHFe24B+roJKSKj/v8+nEdAACaEqE78VnigUeRNcR8qaGQ
Z+68/GHUigpiUVKTfrRhnzdOIujk+pWNvby0rUfqkj4q8CyS71ZQ0HXr9LJ2EubcvZj5wrdsetxh
zNCvHZsBnMOjZfLC6VcnlTEvH6CuolA4xET58gGQDAvyTChhg3QxmfHA16R0V5fXM5oEVvtDCkB7
N2KIb9zVjJaodi4QKzBNF29Gvvff8oTLvrd2Db2FAG/Jt0eRpr2cS/aUMmqqddvUrTS0FkhoTIUM
u4iFzZtLmP2jY/2fcodz535qkf+xRXoMdgmVt4gB5SOOn81IMQcIuFjrZyK9FfXCtDnWGuQiTuiW
CcBhrrEWMALFNdCJlbNVAqHytYLgZRK34MPEdWSXTqET/pzs++XgLgPA5pmWa8OXYjDyZTB8rc7G
meGhkXly81pxaEHTtyutDf+vaqIIc2NK7WwOf1nlSsm9PdcdXsFdY68lDmFFsQSzMV+pe3dHi9bt
+fEunxfS28+iPZU5lsPaEi1jTZzBW/eAUNeGfzp83r5tnuo8J9DyK/QZxDnDT3g3Y2I/8209nXia
pwERq1ephY1CYkv/R0aYCTfjtgWnCdMcy5Kg0jhMUGjaiQ/wPh7UYs1/DaTJh0CIIbQVGerR6ZpM
VOUsA80Cl9tEuJytNgBPyAeed1ncJNRm32laec3uMh2KT4dcj5p/M8ej8iCXfO2MgaJ+t3aLV+pW
efZ+t5gGKumdWGQc4yw5KkENLESaSiLLlnUaf4hCUAftjeCpQZ7y2aElNPFNU/m+5cFbYYsEMRY7
vf8VYXq8joPm6mhFUjPGZsDz3CCMLNlF5eLleukeAIOkAwu/RhM2mfW1/sShIdQY8m2Ft3OrYFtY
iuRwyAksXORjfqOAdVCcqyCWlfjTEOc/CCjA7ccEzdytc09O2F/Ii90PD7KV9l07WfaOdaRQ4oK1
Uy41bKM35w6ejXQGYDVZOTp/fKVklzdMRFUdaR8fRvHpGSFEupgx52HYUYuPoHK+PQ6it93/2KxP
7mXTpefUQuoWqusp8M9YJG+xn3BM3tCPHcOkmOdAxeYj5Oi9AHaGUvpdIUnvFDdhuoA9ozACqv38
z3U6EHcujbTxHZYnKl7pNIrjKSTwjf2mL0fnD8HHymVWM+4+A3m699+W8ppKqGzlBZPjpw2wOGAQ
AAeB8Gyc1KIpbyFS8wKPGZIglLqaVP5frns5UZwYCbvxQQB5eijxN6TvIL0xfnYmb0RvNRmOl9FP
QegCfFqHYGoUYWPaXaTqMbalLplVWaAapvefSpH2OSBXXyDuyWPZGdZG4HC3s/qE/KL2mZ49zzvw
De6XPJKElhUii0xFg4ucyF0vmsNhW2dhFScw6OS+LV2Sm5Rfq4Szz3MyHoXvh9OtUOU8s3YGG7Qc
5LQAvAzPqbpzOK8AtZjKuRfDmj+2JzI7lVlSV73G/P795u0G9lzHt1+aT0bgJT+28Z8wwr/r/Szu
n7fIArCZ5PrcUBev+4lEMxNghdk9aXoo9nEDO59Ha7x6mLKoGP0YnmFmJ2lps/T4QMkpubFLM3DB
DvJxF25T1pIaOrSawVMSim2PJ5+piY1LgXCMH3nkRtWaKiLogdBNk4C2jPgb0OKJP+/n/WwcVbDq
F0upwDM3BDTrUIET/RD7+NTOt60CnqyKnIUJQXiXuKQPFB2kJW8t5WdvjTeh+Qz4kphl4krAolyF
T3Bki8GlppePc3rrSY8HEJIbKRwHB249olanEQIK2B0ZAj/xuN23LqBCbssr5Atn+rViCvsOnoyd
j18PoiT0v5pviuMq5riaT9z7FQj5dTqhMmy8Nm2AfbZedGWrl5oRkLE3E+uKibgvafoO7gXjo80h
6SbuZg/tdDi00N80IWx4ztmt03HaO/FJ6rgNkntR3NDBqc8501y4hotj1sGV4EqSYY1FcAz4KeDp
DAbfGE/VLxzkEYfJkHF8QpE2gU2nl0Q/ndQFGPLBfBC66yAlOEHOc4G1s7l95p5jm37HmxpdV9Xa
SWI2BeiVYZXRPBZLMSZbHdopoRlhaVtFk3C2Y2Pmo0zTk3MtqSZHFZ90if1yQD0v7ZBAJIDF8154
3TFUyEjKBrEh/3rXarMCxcAV++bP+Ltin69g986J4z+U1RB3qV+WuqnYg37ISgsvyXn723eDmHbs
MaI6TGyE/nXiOn42/Xd76Q3/6o3pl9WlO97Fkjz3Hjw7uxuGgLQrq76XiMnowxOSEvHnz+Xs9Xfk
ZXcMLTSvesy3G59RPb39EU1OeqS1BZR/BJu+v6a7gdXhWVh9BnSOpB/J3lTfpipKKZLdHdn+w6cG
Dkr6HaVVV2KgqBa0zsVMXakWClzOp+luy9Oa8QUHXM9IikeBslZy0LIZSPutUuNizcTtKqxk6qNy
2Nydr3xlhjaxpKNOZmtWm3WXTtqnHI3SGXopxEe9PwsdYpEnbzY+qfaTk8ggA6XyAo0NSqD0BAi/
rbMKvgaWh6cNnMGGRoLogZ4NqvpWZo028SU8YVK3vK3ftKb8avmBWy+J7MATGajSjo2zfUhsz+3O
1X2BRHzpvsQJZFl8XiMS7CexFPXMQYtQmI/nCRLnr+lCaJ/4dwP/jhwR9YkopW7Lvsh5AvWZOR3l
t8dBQ1Bd0ZFELXEYXFxfG76Wd6kJ4+uWJqn9vRcZLbLB7sogK5YpLOfwUk2JYbSZ8f4w+9vohEI+
+IKDPjPpLcNh0WEw8l+68TUpDlB4sEfPtLG24v5NmGrsjyBXHZbHSh7IEfUgiGubhMWBkqQqO5qk
QB5fqYz6ihlUmQyU+caz3Pr72Hycsgi0sBuU4EHBp1Pmoxm/ttIQgGnKlvvCwIsouZl3VONm2fev
rCKY/cs77zWx6DYOSIJI4KuXa8AjPgcR+m29876V4bDmq/JkWybqXwuENxsLdAOu/P/DizzTRN1l
gA8SpBiCKr7fmR7FX7OfgTwFdTKEOSG+1z4cPB0FKZPXP3Wj14y7Dav1CekLWMKY9ylOA7djW5m3
9fllgTUVgT+gXEtJNhcDVLqdjaDv/6O2IyOjVaW2RgV9lfiyJAY0rzvboYvTj1Q2VEPPNZ5X8iLd
ZzRM+Xapx758tJFfw5Hpb83Zngk0WPsin6ua9MSSo3JSXC88ucUT95m9SZOIwsDHxDLgu+AD5BOy
de7abd2xSPPwzl1+YaSjpfU8mDQUMzEqfVm30XJ/5IHOD1mJljlXtJyjGaauvLnQnW/fMnrycuTv
tT9/Gu9Tbf+YQP3gD1C9mk+nmacSRXyQHJfp93iHTbg+z0CqWo0Wf1vsRX3URThMIULEfdHMoI4J
tLdy5jUxqFJ1JkKCr7CrO9Qy1Ei9DInU+mgwtJacb56A6d+e6sRkmR6ATzrhgfxfNg/5diC7KAru
PwLC/wciMSHueS1jlsOtkQOFj8VRrWYs70zKAJO653oRAxY3ldKoORkWW2MZs14Ee/v/tLxl2ZIl
uJ4h9q6ZL03Xd9CDOUHWSW/v1rcsCThITsJ05/ayxYhjMJdmbKSflimFBlCCWATtc5QqvWEJ2HnQ
XWGkfqtXDw01wVepki9C6Ohy6CnCd3/9FQ2nPJmYccOjr8NMOpPuvFkKQu/nPxcRtAoMw+nLNd7e
bfZoPSDvrzRAjcN9AUBXwgFF00Jl443UDKCb+EoccIW3eqT8qlCLTq2AmZSbCYiaLPp3HqwD5Kwi
+Bk8iUyiHFyoVLBm1sC3Zv6dPvkVpupRXLX+ib0z5DHoc5FzsigaUiKnO+u4fokolVPutBZFEpdf
yoEdjop6Mp57YzI0Q/ZVDps95spO7R2weuoTrax7RmihV2hbjSCWr3Q2Q0hRKMxu/w/S+DrATGha
JfbuEL0dpZsMNbZiXzFvoYUs7xZKvD+PqNZpa4QnFPirUcmg/WuxHlDz/KCBZLQoU5ADOL8vDFw4
3jlooTZlM3glLjCbZvtsVY5lwtAZyuwa/ukL8RQOzPezdsgLx5A15iOxRRQY4FI+TBjRCRx5e6KM
l4n6CJhBmTQ+6XYBiIbr0AjUGZUxW9Ecvx2Cwq6j+q/XTPeS4esUjiZR0N/3O65j7s70b0nImjfJ
OzrN/y04Nq/DPyh0m+MOlTPVpjSSflBtsavkywQWjqXOZ6QGy7loI0OHgKMhoE3Jx8SpQZzo449w
t6uk5i1BvlBTVr/pIQpU7ISiAzeRNmkkW/f9ZmJgh9/xepuSoyEuha/XFVWRwXtj33peO6Ca41xj
HYrpP+nylkXhpt0u2nN7nnrIrmRC5tMmMTdv2jgFzeXJz5W+to0oYiakfBm8JdjERuYd4rX/L02d
EhbDpKHp/YkU7YXtUXqGj+qej0XtgyqeW7YVTQG2ipHYmhRpS/j3FPiQPLXvWcPuTgr+Fp5IVyt5
bn9WLt8wyz0Sh/xRQhSgDSO9DGWUK7gF355+mTxww77SK3fKG1iB1RpTBC+MZkG/twxu1A7OuJjZ
ktcNCQstRj8mUbbgRoEZ09dXZLsgKDZDWkHSBSjn2vpsscNH8Wx/JCJiJdW4IPOaCHN/TilTeZG1
qTIsqvJKjIdsrRvIwJyma+4OKYrvV+7keDQ7kO0+Xxe7U6K8Z4MUrngtq6dKlSypW7ydTc7jsYMf
yx2iGFKZrvRxKsdkC8DvHam8kL8fyIakO4WCsat75oo1LqQJuqELWxi+4KQy14TuynGWhNe7feyh
/OIUmpf/JB3kxX5LMMhCoiqtdYLem8qNrLnQKfwr071gW70hC3k4TDJz86sZH/ZX6ssdsMPswLoi
FJbUHKiQX/NvIbgYb8EgnO6i8u7QsA0JrWEQs8LBYrD4uRsLkGZW4ixsPQQ3pj3NTwUSh2Gm7iYF
LV/UCfwv2TzUUS92Vig3OLbsWdlenXNQiaAmVfMoNZsHUNGcqZdVQQjLcsfnWFQFdvfziEBdqcis
UqpoQfQ6Epp0o8JGqzLkDOkA8+4ypU03S3B6HWSqM3R2M8z4OsID0r7HObpyAQ22nCxcMDO1uiPA
83quoC7oipBaVT/I/bj/xZ/zzJjchEdM5IZ0NSRwV1oKMZBc8dDMD3jGT+6cxXHi99fGPhzDR1xs
vm9cXhU6qizXmSgvKag3lfEQvzO+xT8DIFzx02CWrrh1zJSJMXxD13yjIt5JKjNscssizC2eVqk/
qrZ0ojAzxaILYFxKzQqJDISUF7IFxktp4/Eniz1W62tO+tNKGzgDNnLOi207Nwf6jAPLTtjg9HG3
Xr31MR5lX7y3gZd9LGNo5c3D9Kkzf0x48yo3xCI+Xu9vqGKng11Y79kIbNcn0MbIfpIhc/n5OFPC
djXeXgRdayN3AuKIxXcWRAC44ywi+55Ry1+M10jaarF6YLHXUQGeRmC9WJKOcQ1xJOSER8rcYwT2
x01MA3Ym7bY3u1y0/1T0FYCbuUscQhUNX+5fnVulIo3LwhwFWE3T1c/Cbu5EgyEllPX/sPmPpyK1
eyv4ymqgRHydi48/YI+7I6hV9zFCArRzpeyPSwTLBxHiaUvLJoyO4pyyqmDXm/Umpt+b0C20xBOq
QmtTPQkxwcE1bXvEMikuqA6zSYk3Ka4p98mzbmUMElqTxpx+KfT0wTbTg3K07mcu+IRq+PuS8Snn
Ze00XosmKHN0dxiah5eaZ2Y+aj/mDZfOzU2b/z42vLaWgdi42XLKh6enyWPnRLG4pgFhXEAGvjCd
95P1LO2KNgmmmSMbFCges3DgD0jnDIWZipmINcKxA6pdKynY0EQbED9VyoIiv8COU9Kuhmjp6894
GpSILH9otCNMHEO3vsHHrYa0vI9GZ2iFNw48UbzkhoMXdNbrQ81ro/AyYjsD566mgwWK/WwNxdVd
vByXIdaTRgZhvQ4VXbzFerG8uBfte/bpxBAALrU//ou320xep/5ODvIISYOG4dONcmIh+ttadpfz
z1Qd3v+J2SkTewQ7soFBi/+wko1KFW4ADOds84+XQCo38tpQBExi1BX4COXk4CKEVNPzbsUR1B7z
fLtTkw9pmiPmXC49zPIEOAClfxkXH5auoOLBsISdKDHJJo3jUrj7vDf+a43bel1T5biLhuzXfGl8
3L5XVWebNlcx/8DYSZYalt8PlYfiQP6rnOVyOWsyRRvwxsUFkGJcj7MKQBHiPMMNg1Uc7Yx27iLT
JNbdThKZlLu0PPNS3XX4qdDKqSVpazXjKFuu60esBG+W5Wtwa7JfgRjDJfnukAZ9JsBZsWjOqUS2
ia7Q5xzds3ElIpsjOc31Wj/UCxhGG544wqNkQzwOZ3miHivB+1DMkQMOlUfhMcyNFjhqby8ObPop
lyVrhz87oDDQOIwu9ZAYPBg0/LalLXaIC2NkSChjL4KnmEcnIOv78kleZ0TVR+eu3HFVlK/pq0iq
EBkHGQG3e8CxEBa4lN76KoEoJviCIklsoIC8R6sFBHrJQtO9FVsg5svjn0adNQCmxxYq+3n6/mG7
I8lsWGCCL8PqND77WmQHznWIDn77XcVyGgz0oh75ZdyWk5gBur32/15TvneYdRMg0/4WnD95JLMX
oCNxli5y+YVGI2OdwmDiTSWPDp6FZOAu22iAuN+WAixLdRsoY3EJ4W1j2HsnLy002GD6bU0JswFS
mXa2HXSwx/GS9JtcgeOuSNlaeH0Jp+p97VOCpzn2N/zSNe5Htolmx1lafZiP0oZVOQRqcmzPpYmT
zochW7uCgfbTRyJMyr68p8t+fpoC93YaPiH/CzKJy+AvjvSboGuUO4ytB3a8QH1ADb4zVzxRxS3T
+OUv+UzOxRq3pcsSatL5tDIM/SUjeZdc6syNAAB8Uo5Bhr4m9+miTx5iyxI3k3y0zCZdD9BsYmap
WPIhMd9a49+NdrJWeBktbiGJZTFApJX/17NRYRrkQ53OGVL8PLoJCqfHgRqE+OT+pdr41NqqB700
tZVnBjo6Mn+UvuQnY3PImXihBE9XoUTfrExFxdPWmjmOXd6sKSDix58KQU3hnYsUuxHLQCXy4zf3
4rz9wlh69sqgtoRYcOfmFEKyljRaTZa1nc7Y2XNVI1dvpvqcub12L2pa4OyAm9KydwDYmkzQlq6t
3KfEVHy956rgkINtLuYpk88BuGFWf+qUgJRQLfu6I6gTpKrB0QmorRi/Bx/TRPcSHSrd8zdNVzh+
4sZTgmweOxFz3+sDig1Zn74W+qv0lUfd0zXFo/vPOTjvnCULa6CD2VwcJzOla0RwPvfjkIB/dEBB
K4/EksNPsJpGiNo4bGo8RhAV9g4t0V2/4pst9OhSl1D1aaD5FR2cJiH86zoLBAh9UBsr0fsYRzfx
Qi4GIRj1aQTOz2L6HNoCapTY5tWypU9j6C1IONa0x/1su/7q4aYGV/q6gacWl11niVVysy+mcUOy
JHqwavsB14KifmnIV5+6Ox+gXw7+qYJhxCBfjcKQzpGWU/tHtb3Hv13pdCWniyepE9veYRnaOV9+
+GfIsm0VutO446hFrpx/5bv272gkJKHULxj2CAujPbCPuYcfk0Ol2St60ckCYRtmBdQTjD2qr7cb
84lpDQkEhsphKtD3OEiUi99oU/6q2crpJBwHUDJjHoPQJ4SMS5hJm8qCQ/7vlVf4/G/EJShXrATS
QtudGPf86HQSzCXOF7zxkEG61U1EonK6QAjZYumBOPp7+j2vgZIZMzokeE52ZXaYlRiDhhXEgL+Y
Ksw83HDjHXB34FZIDO4zdSc7Esg7ySHuRnl4+Yj5o+NjPPWh1ULKYLwMOk6048LJUwbpsKBOjU2+
iNgzw8nONw+Fj5ZEFLETxmJmstNwMlrLgFnTRpgdANg3u98VXpvgy6OqjZSe5kBmI5Qiir1RawD9
bfokBzIPQjBfhmc0fHbygWj3Uyp3RX7x8SAxo9WoFusx3A1UP5hUYxjsFHAJakz8klDimsPiVq4O
CgNo2BpmB6VDppyw/0jUBdaAMIWeFSKucBTc1HW3c9XNvRbWvLBZ0m655lzhuzm9dmx/zgtOJMMO
Bii8WyX0W5V8r5P8fNPx47O/k+qt0juv/svohpHvmbh+Ql8cprMNw3iv3RRZW5mJW8xQm2BRnSmr
OVtqQIch85jbkGgNzel0A6Cvgi6rpLaFGCW+YYBoi49vwe1Rn23H3y043bG7uQV4PmGd9LlBqivM
I3Fzs+XM6D3dLJrOvKUBoRWM76O1eRQkY8/G8YnnpoOkf9tWSXRZRTng1WdG6LJIOpz9IrcXwp/p
S6tHaVQlvK46zNQhQC7eJ8V46Ss6HAmCo19tG960qelBu9XZageyI8np94RB1m9LvxyxBlcA/P+u
3QrIgVHofsWixIQdGdv2K4tLNcFDzOpmdaIthmhwzjx0VzCsTWX0kYnakfq9YOO38kNkGxXQeZsT
hzmH28fOnAwJHhyR9r+hFkocsZtDO4B3zGHQjxta1A5PgiL988nqprXwQipPPs1m3Rs9A/tGpCCu
hRaz1nTQ4pcoKpCItppufYPWs5N0s4ZAM1bofi2peuJIDImlieIAlxfZpMfva7RRF/C7tBvKGiV6
H1vDVABTXH5cL4HJU7UAle64AqrAPMs/h7OsjkdR/+rP+/4LKpZtqzfRs0NvL1DsschkI7Z0X/LO
3EBkMsjpo2V3grspyqgfZcSVuTTvZ+OVijxclhaKI1KhEZUELZHTEbBfemVkhHyXBXh0s65HfqZQ
W28T7upG2Yl4IxRxwApXIerS2OzGO8mRoz8iO83VyZfXEBQ3CMo3hAFV0OMz8ZfyCLIe3oZ1aua8
Tp/lNStN77XZDl+zq8gdJ3dYDm+m6ZLF/bjCOLf95ucEB4XN/WScSl1bZa39iicPkFzTsCNClRAU
2MrmxmoBQmLx+rXZIOIt44yKwHswIc2ktFRJJwz1ciWSfcrqarGjHDdXEv/060dSybQaLl6Ly/Dq
zsoK9PiyXMvFhQjl670/VYbyAZ6s43FlygsuujC5816cGWmfbmxjq6mAs3Dqj2EZ0d1MPHO1MADN
QvCK3LHWjBduyYova/6+cvmLatRH2ddNojr7sxlGVh4404INxreD1AzAfDuco0ixcwmwkyElhZEN
Q4byBAiE6q0Ou7LIMrZJYh10ZsnmEtaJydE0jL/xBnbL9o8qqZzkRpTI4Ji95DvyrbmUqVAQy3TT
12lHpjDws+1ks/fkRiscg7/RpPsiC822gvlNEwf2q+ZCV2McgJTuqDpYo0V2IiCklUiaBniuqIxV
UZt3b6iGhqsuBNw8grE0n+pJ9wg9L2ylYvt3tN66HkZXYHatZEmWB3Cy/VuqdM9Hs5vQ/u2ggME0
zhJgYQwmiJkhV8iMrDS2xXV4RDSt4tbXqI5NMtVlPdG/SaN0hy2FoIG13cxENlcV1Dt7riPu28HP
GvroliV4B+X2aoWAR2Sg9D7pZKDLMy9R30P2ExoKmTPXS7vyejGqRmLhlcxbTHtzFXSnM5ILlC09
xC14Hq3m/1Jd75bd9Goh7z/MvMc1CK1TcNgKR23XoBOq0GBIwFcAr+j+rVjT2d3Dps2v8gw3ys5X
6Hy0fEB1sU4qY98yjqtnCJy3CxQkM/FA6xNJwe0vXwtow/ZI3671FcWo6taiW0B/y/JKUPJxaVa0
wbtIh+hjLjMXypIkDh7qm7MqfUYKnY/yawWEdAic4v2Cd2EYuPkrAe3AnJlvV5vlQUntAqIfhiLO
IKCy+b+Nue2fPoQnjDJqirdNuC6Q+A6wHr+5+FEY+sTZgQlK9ZQjjG0XlEacy2koXxWPztCnuG4z
BOaO5GI4ZigLUPs1xa3uvZQ0Kfqjkme1tnMtmj9oE03QPoOdXooAFoJdpRGBWt2Skrh13mDK/7uF
D4wjE/E4BblqAwZ92IatIE+NCiaMgLVC/oR7HwjKycTt6RDBqaB77+y/8RvpK/ervsqZxYP3LoHX
amcmQ/ejqGKvdAk6GD6rYuQ0LOLZzTZwcLfuiC+huPZhE7efHmVE/c3yDfrxe9mP1ZPi69Y5w6/a
U1AZOHk9xI2SnsvdEpmFtwGl0ePW6k1tQie8u6xLapbNWj+Xgfmg2Br05zJisrUfj0xEmWm7Fzln
8GTlvpBS5Y6DHwCj83X10HglIlqUFZv30CrXJV/KkfsbFzzDSwY+E+C78+GN98eBrewLfKOsMHKt
wXPomPn5Jy08jq7GASDckWHURjJVoTHj/edNgcTuOxAAqISY8demaKdUFiNLzgHebUm87HGTEM8L
gBACrzbzsPyt72HvAt6zqaPhdfo3j7A2xLpV52tv2EupP/eJIVi/BgXLp/8jm4sS9EAPph/XtlBp
4g1LIPbkWAUJpbdEj9Yq8E/nNolB92QVn2ZdOuUPlmK8ralH668k7+z7VCqYLmDCRPiTPsUpMh0C
qP8Y00nEmbMC5BFO860w+v9AGnxu7u+zqCHuxVrIvcDpe5CzHgru5ms0MGO2dQSsgkxK+usqqxGa
sfKYjXbmlkgdY5TEFlFRwOd9+HSk8hk9XtN3mLExlTPCoH4rc2xGZ83ddC43gN6KaiWnFjdlFXsb
0MuF1jBuZEbU+KO+siEjDdWwd9VhM2X7t8xg5RDwAMGSghexxnpGpBkadAc3T68E2whBJpEBBOUt
hcvOIHZ5iHeZBQ0fsYI7ToCZbSv7LfTyYHzhg2O8OHtFfLmPTocSyZkm48FpA7D/l2P9MOWj8DoP
IcK5+8f3hg5p6ejZ3Q55rNv5Ni68QIp7Y32CS8FBezEkH+/lKwGLUyALBkvP1FDd0Qe9n6CaSrB2
i/sbZdD4AtuWJEwqaaAZUoL2myJ5pq1dk6m7gMEzrXlXfsY2SayESyE68iO5lOzDNAqiVnQespW+
bV/cIdMG7N1cVQlhef8nB9i0Lf07AMtU/uet+NeUOqPiduMRwcuZ5SMsxgbxQQeCREW7LYqElRBw
W2UsWji3Mxs2oRIQoDhUO27Tv7eVS3bhvj0OLHdaDsoZrG9SuYduC0iQU9ZIBIoxf8Tp2++NcppO
sCRmcwKw2M5cPCZOb2MkWyc996yhRe7wlk7mIg5AFrkFcWBSsLKNFbhXr8ttl7X7/VZMhHnH1OYS
ip5OYCz5h/1axB9+17Mc/O5o+gRX7TLAI3wyjPkH4rS/nNZA1/s8YBWadjXW+tZqU3QN567itpHf
oHJOs5B3e2M8/uqyPKe4dJFrIqYc9gfh9ko4Ty/RmEVoePnhGNK3cC8OIOkmGuRfD+OJ+aOaCdsS
W2V8bVg4LE/1+SqcgBHOZV52B0RWtSyBeMVDtptibYez4ONzFa84OmlM1CHxVogl9v3/DOOM97lZ
AfBxVJADlBzktprI6yTVRyCbHgIRx8Y8MhMEHUpQufI2GzKyj1XPAxW3Se2/n/4mIWny04nfDkmb
lbotX9gOy5y/HikTF9oIrdhOafDGdfQMXMgC5Yzw+iSguI+lCXXBMbg6mfm3wxLbdy071ZueNNhG
E0gZV0BT7y6q/rk5uTfcQ0gm07z2Wxtm8kU5lK+iGILSQF90/+KRHIYtGUGq4c2rUvc13CTEvNCP
BH1DNpUcwS4oOl/gBRr0JjABClEVFtgidc/Gz7HLXYJtlrZEZYA5pTRRAJt7oEFmGykEuPnTvngW
2K57mpS8j5X9kI9UDjw39QftQlfHqw79fkIGstnfwv2uiYwNdG/5LLInzkZ94j4YDqMrXgt4yOrA
qkwp228i7ASBxRRtznQ09qjUjB1i9ql7Cnnz928wZyuWTpYeCpLD99BdqE8SjYCxUe7h3UwSO7qP
4bWFkLq9kbOFGv+JCt/4AO011ANZ5Q+R9yi2MaH5uwfkybbOW48yUrN5NMS9sohZrEOXmoUqAzeW
Je1KxpuYuvWCO/3X7CZ6vqf6FHC3faJzaJ0Wufn+XC6EDWPqH6bUsnB8UE0S+Plwh7SFjnhh7ph5
w1Rl3P8PpYuLd5J+s+fOk/P8YXLdRrv27AAmO1nEC7cu3PZTc74gqSc6z5lY6X4qBaf7QOYbjM6X
wbdTeIMp1q4cEkgmrjmhC1S7/jlmFSxpdvizVa1wylZZEp67qp4O5LKaVHWj+y7V93OeI57VT6xC
TifiAvbfKuR904Wse3uyTqoUBFXBIuSEPG3vr5YilnseAsulmDIboLkJW+d/nhjB6WV8abt/ULDf
q6aXHRfv7tRyBw5b/MmbP2CFhruM0YOIxXBoJmRLCNQsMeV6rFjvZzhHqo99Gu/Jbk2NHQCC8Znp
3O9DXUIwBL5LJOW3r7BQFDitbDVoiEDvEpoMNLhzhJ6bsJDP53siEix/1Rabn67sw1ggBcf2foPi
ygAES4Cuq4gLOQMy/TRoHSlk88PvRbG1cBLOb32K66SkcZjh9TSq/HtiQ8P4vSU7apGRSIsT60y3
+khojYK6Ie87o7jAQSOYsveqoFnKPDsnOde5XbThuhmoCDD39BuWvEGEnRaprwojE7jSlt6RQiKi
vhJ9w3PwVF5mNIB3yLGRswlAKuD+HndKAdY4Xl/pfk+THwDPyKkEsekuBZRw3JcJDttD2TaL6+21
gBlHAZjOSmYuv/526mvD/k2KkcPpTatV+WMupafP6u7CP20bSZiejpnOPNf4KAKWdZvUGvLuvxeO
eKA+dcmEm6DCDc/IEPP6L0bH7IPeq1MJyukunB8EuuBlnYijiJffZrVKq5LT17cNxH8krS+2FHZv
xf4my6HVABm8/dxUNV7FHQwgdbdiWWhqWls+b8UBXUiH5WEqXRl9bnrYeqttYT53vK3z+2/qY/7G
HXYGban0m1tqwymjtj0l9nlEf3t9rCt4CevzkXIVnMgzh4B0x3TFIIY2uMGRCHS9i1IoKRIPXQKz
A5i/WwDlzSuevCxMvV5yStOP7ILVHkhFIPuMeaxf4RIfRBqSL6E2JhYXQL1HSLbFULeSQJM/6FrC
VPEZhx5f2ci7bx2nsfiOKyD63U8LlmDc2GYvKuXk+8YZI7jxSWGG0MvyROWsF+Weav8YnlqX+AsC
/upd4L1+eUVg8Kxfr55VOk2N/VzCKphToHiTsrfESuhS88vKd8OieOSt6Cj6nJVslXIC9XMY7D4d
wRFL+Xb6/ob3gq+FpwcPfyFkpVLGVp3CVJjdbNaB1BIaG3YqUfeSZwas/+/8GrM7whmPqIdQyf3f
zvgGR5Fu233Jo4hysvfjBn+Bn09ta6ipGaIxs4EEL2ROLTsHDewbSs5XQqS+4PPmcIPYKELmyxfM
mOauJmkx7sfmRcV6XKQdKm1ZW60DA8jCcz6Y03y51HPTMYDXZe/QdLD+lQigptuuj9irS5eeNu9y
+Ld6CDCO98TGr2aqAiZuH+OUBHVeTqxUf4D4H9FIr4p/rSWaTovtPoAcKWAk7Po/KKRdtvtxZk1n
thhkKDQ+VFTP6hJm3aKvSCE6Bv5n4vBXaX7YICu8lTiufuQpdb8O+/1XZIodwo/cPFYCouGEhPhm
sr7mUF/p2dvuB7ctsvDs8CzxTjRjg/chLooJ/IBmUWPzCudkYrQFJu4uid+nEirbpbZP2Nrrik8z
JxmtXP9Y/b1yd1ol1X0fk/TzA8U8I1IGdi5gTbFqZj6lSgTp0ID6ghgFKyTPhHnuiIulCyacdPrN
cpIU1S8TcpUBlO1/Afo82aokaOsCpheqNXtV/LeWAANsSx20CehJgd6NGLTNZRNiQO1lbP8pAQjC
GdHdBQeuN+7YtO3dqKLQPLlODII18efyLRFWmsoAGX8SY/vHXA0fUhkMA9cmtulS+lgoPJpLfG50
B5IUODAiBpPZYYQ2q3Dro9lBKq/qK4thfvcwDfjFoXB5T12G3hInNT7wMK/ngqFaOczFGKCqiAqM
sxdnpcaW52MXdC7dFx/2ICCtx8kw3NSurRmFXnuRL+Hx1R0GT+xRZs6hASVUe4mJVI6KAvmhdL8x
bXiXMC2YCvWEH1v8vyyjRIEQ+3LippqUhzU5DS67o5Yj6lrOehPxEpu5lZgehSIXivKbbUFHsrMN
LBOGMOgLQ7u4vuOq7InE3MpWVcD5by+6ln1w1MwpjTQM8+Rhk2IWbqTzpx+vZGnTSkxhe/jTZBDx
Hem2m4Vg2bzF0VLqtOpGE3yQY9fVGTbjlCeerkH+/4wyWq6OehFe9P7jUwqozfM8QTSUjFVpxpZi
347EqItBXKRJlkYs7GkPQ2/EGuLvHl+Lwkd+Lq+KwdUNf9Qkotq2tinqhUo8NRuBUHyHCH7FV4T7
oZpIlEnFpdFXCVXar4nZ2a9dIykdZ6SewEYUm6WmzxmpsxoqgYGIQpU2JoH2FE9Swv3Tryl1wIeD
1ZifiExFy1W4BemBAKa7zPO35d73tJnOOeIaRhRq/qpALpJWYU9zZwrDHlQtDymX/or1FW/NrQQw
G8hEnC+OCQbaG0RnkfwRLGcttb24/tVkPRLaSWE/tQkw+zqnzrOant7XtxsgjGrvPpqgu+UEPn2U
LgrBX9HGYhVmnaXgOUTV+OYCCcqlAa2P89Vn+mSLS7NXdJ/CQFIGD9GHXU/jzLHUg16Ikkc6SBbU
O8Enom5kmyj3qYCmJLtmkMJSLhICXAybvL/HChY2XDT07E4XnXUimXvhPlbKe0lOd8NNq+sH7l0Z
FiEFu0oZq/nyDxm+7fdUC7TVwqj0oCX+rWylpARPypXfDao50opM256o5f5O93fRxHZTK1xni4Sx
mVLWDbR3Z3P1Q5I1bDMJn+zzkYT5NxuDZa4rEkyhC8Jk65xKdfKRrCzPTA6JjToo14RVKSL4LcQ4
ZMnJpprGRqp+ssxVBYz4Z9uSwnW4G+JwPYjdzvHAqs28wwZ083ToJMY24A+cdlqVvJIWpAwlp3NR
yNdk2329zjKOtBH9+f0Q8rEUGh5f5bc26tDyaQngMUE574D55G1WXUreZSwvT9WslZ5qEPsD4n7P
VJiluJrGtrX1Xmv8xGvrTyjim6rOVII9ED1BemcogLRZvg8dJTQf8fLvch8zEnFqP+nWov/KpCNJ
cnxvte5JgcIsL8JXEThZkXmoiDJLik0djgzElsa6Jr6F/4c1SuXlJEw3sQNkSF2xPCnkUhRdgRzb
9su1SkqIo+4f+fdfYBkZAh4Vywk8C4FNsh5nK+05djEwIP6LxuSU+JYwJy2XSy7/64wElvYNxwDD
r1pdyAifY4XLc2Bf+//XC4BTZdV7Vr+XKpn3vK5pMpL1WOi9qLFizcsTbV44RtMHmZUU8DPfUsvO
AaFiOm9wT3MOXR+kjYtTz8T0qnNYny+s3Jx+O8Q8/ZA9dhUR6nCXIPLWeSjB8pr0+HIatTCBZuIR
eqC+zcLJ4/o+CSRZZhzizZwi3BikZhfeVTcwVDby62XsTZ2rvj3UCPdXHfbUjKdYSKXQX064Y9jP
m2/0KUJCsjC4CIfuEOQSr2UwCsY2lEPf4d9hruCbBTIJaIbOok31lEcK9r2ufEHy17SEvyTZEQRD
2j5HkOaxq4vbp4AJQXefgxf0axQFDudQgN5lSuO8iSWEscYjwRS7WdytqMHE1D2bWbVYAFgT5uI3
0X7IP8QEb67B/Yy6HI1UqTFz5cMrCukmnGRe8OL91gRPbLlfHV1OtM6C56u9rLLDw8lpoQihRQLV
uRUY6VhbxKyz/gk3LvU73NMTgN02km0cUvfH9qONFfMSvAOfD1hpyUap2VpDDYYEu0y7IWrAHMJG
sT5KtHo4uK6qZwzjD4BakOPS7h+gbMfNnf1jzpiT4IqyThibWwQX3UxQ8+So8vwI9Wu1bJXJldxF
1jfDxKDUcK6Lt5InH7KI/GcjEfxgbWOPvb5XwCYyk9UuWdcgKo22IkL0A6ti9u0Bdb7CC9NT3iYK
keEdDb47PCVavgXv678TZvpL0QfUyjSaQEVZpHH+CNQD3jxK8PkyueIGwsjzFZnv64mu5hKKYwzS
aoQcJUtIL2Uzk97TDtXkc5gCo8hpqNPa1EhK45qdShiHJi99Kcdd2rW8u8ERwZwg3UfbdHQIAVOJ
yRsxbOfENYfd3nmETWrp2kCyO6DovIsO/95iGsWVy+huRAg8KiEo4OY5K67n05qhgPiWY5sbG3hs
2G2cih5KZsR+3+DkUmMhKxqBKScOl2qr/E71EFZKXpu4FZ8SQB34mQ86Lm/3O7L6/sZTG72i+eKT
mls1OopZOwEhvPYiwe7eCMH/g1O5ZHtGEr3w3k9CLipteyE/LDi6RJUIX6bDuUMhttsZe3CLBL5D
vg21LuEY4E4m7ybziiW36ByeeHwWcrFf68sVxJ6OSD39cXSfIk9rMGmL1URg4Mj65f96MfURPjae
gekwGJyOGpfZpaWbftx1UeLgRNnzLo5bEVswH/ke36P66QWQVsbxdqd3Xx56JUQrXfPzpAYFWrqL
MrefmYsHgTF6FQeNlFMpLjnI8DnKZzO8MGvUdJcc2D4N8rwJWhTUG69giHt1d2zRoxsHdgfwd0/A
8Zo85S/WnmyqI1uWYwHFnI6+pbp1N58zKu6uBGLRzGxFow/Mp5uYN9sz7OKl0m+LqhvDuBxBK2Bp
F1mSJZM5r/nUTx3xeYVjcPaV8fBSXK/iTvn3drQnb6tX4lG7YfdbqDe6hKYRzKvX9ZoCTkbA4mSh
HzBU6vJAcO4J48AtHYZKW3BaAwernlpmM1cJ9oK85ryzEhwu8LJzZ4gpbfe+j1D2D+N7iRkNOgYx
5JRajBrpuzDvJxztqg8lFAoOpOf2MD+WMBiEJha6G94qU2ehPwyG28booi/w7PMp+vkXO61c/Dj+
iunkKRlUGGPIevIh8CqgCU/7pqfQcLUIX0D7BP55Q+ozZSy7yasyBx8uWGsKvYiuywu5GINT9dWB
e8aw1GYFWKtw6y/40HlcxyD3cxQ4g8opY36u0+pdDSBvhGTEuWVelw/gSNcr2AQbiPIX9CQLEWIq
trWrXB8tDh0tdocXdU1AkUMyHdvBqXGlt+AV4pIjbHKEgV54usveSkOJAwOyFvs8dlTdAbRsWisE
Sbo/npAZreCA6Jjnb8tkWqzd2OuG/2hXR5P1eAu7n9e+Eo6C+AsPKad7LOVPYXyA6Qkf4cQuVIdE
SEhUX42O4Ug8HVHCjPAIierCmycOuj8MThXcECMuRxUvvwc4ZzOg6uxTt+erkY9/THHP87kg8wBH
Uhhp6LIUueo3S0892Y8V40EQKvFixjcfLT63hLEM/0MVot9U/g+d8WDhyXh95BRrWl+SwmtQpAkZ
R7KTaDwTh4gEqLlfFqbUQcAosXkVW8uuHutrrwXRn6BZZFRcA/y2HDfw6pxOXndZz7VvVcBOpsXI
iBfg6dyy5XfOpgCpEZuoppaXgtbc0q8aplB1Wg7tantvD8CdSA0rGe6xzINZWca1z+4ZtwAe/J64
jQn+HQlVrhdUiPg3UODJkAki1/1RxrynMGfdOZIvsbJsUrmM8IVQWhQmORo6A5vf70C8L2qullP7
Ck/v5wvwnOkno34ptVq4OVDumNfUp+yof9DNdoLqQ+RTkjSdVLyPSc8BhF/dhOUkjucn1dr9odd4
yxvEnPP4gVZpQsO4+GkpWMBR/XkYctdf6KjLwnGUtsDBl9anu2ou+aITWxjtHqKCpiGrLIz6TRY7
x6KiwjBAzUEguMG0iOQfsy1WjpaypnQsTMv+l1qtgILOIPGTguRa4u9nz0wkXL5gyPOLoUxQoDs+
ZXzf5wnn/WWakgRbk2pwpkpURMtSzw8wPUQZ+2eHH1jcgefsYVh0qzMk2HXM1zqjeGZkLYyZARko
+hNI4EDLxARTYOLZ6SZyDP83//BcgBcfFpap6lDBg11vUTmksQLiEO8It/hDXanuWRFKjO2SUG6G
5plypMjNV7gkd66s/8Z5/SQyXeBpx1Nxuby/P24ktNZdf1NmDk+CCFIvt8u/dwpLfKg1kOr9GBId
auRSzcH26Z1yyCaLWR0NR3tyK+CwiP3FlxwVAiHd2K0RP67hAWXpL09kxQqSAym/OWgp4iUXDFtD
RGGHAJ71B6UkfOWBxBskD/XwdC7UdxvEa8Sea1rqqcHPLYvkDbYTWTRAMsR5VxhUUKtkHzIYPMZe
h/wJczq0psLA+mZakUqh4R++yRUpVSFR3Dtg6bbJlVQ9yNJM51+f4J2YDWKqDe7yHS4tOwCKzZkR
6jymHkjYIbdUjZB6EjAZDSC3HqAaqieNYB6yAHtf1T7iJsDuI5qW0PXjnLorT4AD9LcgqjapCOXF
MuNKpDScgWgppmMYewcTn9YmgiMqHvC1rbRz7IzCVfElfc5wtscEDcUTyxhizAbIKpA+R4dVyE8i
2uJmjrX8WFeNTFQ/KuP4eNXA5TA9QBDIyqtqyR4NqO+ODpbfLO2BTS/sBmr9v6b7zFvepsLnltsH
sz1d1cvUqxUB2oNPC3chk23wAWPxEe6eo8jggbCdNbV/cKaAEHswPziQvS17kWLuwfcVSYS3rLjL
0sMpA7OQmnZ9B9Vd1kjyDJS1V0o+/Fa2hv4rI2fsFjsFtcMqlfvA9njbQpUFa53d+noPAqHd7k+s
GSVJvs6TRjP3NIJdn2nh5S3c+E/rvr03YFSDQZzcscpc38KXUfycKCkCBNfBwoFqCCbZUO7HIVI2
EYbU4eaFzPCu/uHujac2JSHIDEPVt2k4xrrxEy88vfLOHNQv1QQIeWrtChNBxskHi03R2HJkT05+
4IaUz8EN0MqNmEzEIeOFUhFWjpdcdjMdhD6pSkDYmglwMsPM1LPACUTLaXyLxRL2OnYyld7o7oK9
3p43BXOBGYdL9guOc1elDsJFe0mZqsPM9BCmXeRDyjLxQqeTtCL8vrg1ku/7ryo7MxlKP2tagdDm
rdG345MwECs56RklVVBs3nDGJF8Y9QtwfIpIETtneCUhZYM//5Z3L5TgaxmxYP4wKjSZ/ztjGS1g
8yE06S2hI9VQgD3H2VDgm1+HJPX4fzye2wMsP4Ms13tZWyEd+esfywQNje3p0FLnOSYWMrTeJxJV
GE6oGS1NOIaXg+hegxkMsYQp6eJ8s0BQm0zKhUcIxVY0r4VrDvUPpk5kMJPlmbY65UW2IZW40MEA
V3Fj+WdckLSe+Ty6wYFgjntjDBrvokObXchoIzBn7HpLxqMw5I7e3Xksl2l8ZxLVz+puIok5TsQO
ULSlTzH3dPIIC1A7aFGEYYzPUzURc0oIOdLV7hUAaoSRVKZOW5lYjyjKBA0T/1XB/zd30gnW3kg9
YSZrgNv4L+7Uui1DvyWKfar47jaarM8qJjnMhJSEGvXisK7CE7BBW0dyOZx63j/N48bYYbhzv92N
ptbYYdPGIEBcz9k/cO5uwq1D09Or4yHSl4I75CcSax9LsjkxnD28e2Huain4xara3HTEndbhGFtB
roS/OioSVK7hdufwa6UvTIUsZ0fuxZMqbvpMqiSlpFFzGugepqIawFxSqXLuZQX2QjdrKa+XGB0e
d7FsMySgUhM4rZhrVFP129iUdYv5MAt1Ta5+uwqiWZf24XwQNUjqjcosEDfgXe/MpCjwKIKqFQkQ
Y5avrxoDIm/nt7XQQjZ8Ve5/ZKh33kWRlg4KuC8m9/DtLtvLKeBp68G8Q9nt+EqJeVFirHP4gH6/
Mp3m3Zj0pEwET31zSVUgpvGOuIkikrb88IODDsmAoW0K05GQC9P8jKQJFQ24upfJoNZMT5tACvPA
u8RJgJKA5OXsw22/UprnsowOAxFQiPO4KTyrfk6lxT3gN7qTBg5HbgaxP8YZiDFS2hyONepxzlHt
o73YVpbBqg351A4z00CA36ZfJ15TZmFjr7FRVwNkhnnLuB23Bafus0gpAs1JlMmXYkEsklICyqcr
bh4nGX/dpIEYIHMfmpClln8TUzTGIiXZHbRooB6r7H+lRWMf1cR6MXxLYxWqj5SUQp31eHaCw4mE
++7liM3rSaviQRIBjGsdN+lN/rM/anm4iOJtAX3C9ZWB8PWy+ophzePFB8jGq9LKliQETRfUcIsp
sO7TrQQ4tdxeaZmHre6m93XGbL5lO0IgkfHdB4c7HE383QV9DbqV+GsWo3VHzLolUvp1eurynPKn
N/QMp2Dryyzsh2688ziZE0K/H1rvUb/6sXtaXxOvppSje8skcSVWKuaBQAmarh27tLKxNf+314w2
Y5XVhteQzm4qiJl9OHGk7Y6BNtaLdtamuycm6pOKMN/bqH0izlh+qeexjGpiGgydVPoNE+nuYotR
KL9Zt4ECLnI1Dg5wm0rq4y6X0USjiVqxyit+fXTQK/Z28vaieoxKEzZaGzWXUJoF7deCzE6y5t8d
4xC2lnGLwtgqgW9JDLKyefAoxuME8eTUReuc63i0K44+z7Huyvej8EiGOhCeTA9/dys2Y2LEthna
ha5ZslwkwV6EjhWC46paa/gHqr3kqhK8jDc2vJC1JXfEa2FIv5P2fguY265UhlLaf7pbabfP0xX3
PxOoVZf0D/uGppOfOQBGcJ642BMXiefFzkWQqklPpppLHwE62bWwjKmR2xshkFK5weGkTJ4gjXFz
Lkh4MbWZH25zW6Y+/Pd3gZ7/RJ1enU2by/RpMZk5Jstffa/kuaNxwzz+DnSQE0h21bWShEVQesMN
P0eUoO9N+bjQ0mCwcW0m02ysKzDIg+f40QXPO0oqsagWNxnd6bv4/hJFgZ6Jos7AAB1AP8hEPv1r
ou0ZRlDEpbTLv7A8wjZKmhzQ1Rpk+EASfdl119ZH/a1GScQNT74i89zINcKdyGKQg6gPBQJTB/hc
TvPr7uAMg7wsDJO7lwGOwFPR6I1sqT+k5qlKdatMRoY71zpRX3V01Lfe4cee0w6n70pZ1fJlALZ2
RQeADIE8IM70hQloyHGa+HSqksf7d2eZmXinF/r9/JAg4pysYRwypIFuf60QOuw4ClX6uLi9/klF
TIP2fApU7x4lY3lcUUt5n2+gp9FE3zHd6kOay18kAQ4absPnjYVr7VUD18JnziQMuyYVQFezVsIb
ywSJ5TvsHrY5tE0j5crRVRtl44H9edNzMaCUwNdBH7hBxXWnBBuBujT2E1KWSHWN0AJrxNqAp58Q
OHZoEbNqH90OekJNflBlJkNcSAyAztVdmUQJmE/hRixUzQV0iuKWMd8VrYznsS668WnfwAawVXt9
p18EGpXqwGCLJg37GDbV/Hg3NtUAlczJ8N70Xg9YEZtGRKmayuvcdfxP6vq3/iYgMs3Mo+h4WY8J
P/queZ6PKd8yT/ZWlJERZ7MaTLtVkRPoyI6Es4pdpcrcPTDoe5HcC6y8Z9XubTqBUc1SRPAF+GNs
0GfPNYzdCbBNgIj8HxKtDoCXCjtkI+ztAvS+vvqo0UFRhMIrzX1SEIPq5ez7ZfscRkHNIQLVLbD1
5l8uUQ1SPB+CgCrvftgsgVsqLzhU2rbrci64OLoKha3YxEd/LjGw0D42CAXEscl+5aAY+0j+INo8
YqZPkV1Lrx1d0erqF3ICvHjY5HBW+sStxE/Pu3p6sQVzxlZq+ydFrtT1Cm/q43j5SMxjMYewjkyK
2PXyj1n5Xn4CGJJgBKSEBR2teFWjWoxEmvqoe3dH+wUgKfZEzvnfmqERIMfzdCteH8A90ffWFFFn
9jjcfmnHgEBHw0vIVtWYmeuxZpGNpv38Ij3fIb/kbzK5w0HlRaWudVScT5WrgYOGEJ12TBfbos/h
j1vYrc7L1u+sPPJBTBlg0wj68Egd1Tay2jqADKGzq5VyqMu2xy2a8x6b/AIE8WgLltjyBtA/Oihb
qo0mOwgj1XS3tBB2Qz78iOIG83qQtYmu+o9RnU+0DvBroOuCq1IRFtVZZfUmNt/JBg7QVCXSwYDo
IkvG1+zCzUi9IBx7k6qL8yNtO6/6wpZwq5seWaLkZnZaovjxPZoIHtGUP1K0dfiMUgh+DLYCCxY8
M5MDQn5zJyfZW2cvL37XYpkKoMv24E6K4kb5eAnpSw1Iv8tqj4Br390w0Krjc91YlPxpuBI/CQIp
58AU6qk1G3B101YIN7zFZd8kxHtYvUtNYt478v72nbZpqyA0JcRLAgUjsCIzKYsbmHJvimK6nyZQ
Jd3+87Su/86GbmE2BFmAX34Kouf0LIHw9EAd0yDJ0ueRRiQrCAd6aoYrpTnm+NFtkVce9KSFQ/nZ
/+9eWieAuqyto7wlYNpFllb5si9xrX5zT+JHiTU5Uqs1FXfbNPAtbr71386vyg+dlvAdMvJatcwg
vTAHJlmJ7a6lpcxyoyMsxTQn827sgi3fhU1DENlFbS/WnmZpcBgjEcWTPPXR5KlHt02errOeQjWP
9ZmloBLlYBrXSLhA1Y6p7u7CEi5kYLb5iReSNWlGYMSAH4LxLCv+pbhIlWkN/cBcbitQ0Se+dJ9x
9V8oQOKaTFEfariR36pkqd1Jtr0YGzR1/7kOw5mJ2PWuYEWaGVe1IiEM1wshK6Qotn748VI5+J3h
mKtz0rwg3K+8iJ+nDjkrIRB214FNHcFmjPG6uvSmMtaMh76whU2HkZDYM6E4FbMmnCy60IwrpoMw
4WwtF2iAtTk/q+YK2pSOVn5Y4RSB5sLJaLvcOmy38KP36lU38CyzWF9RKowP6aKbu6fpTSpye4zF
qFmMGRBMjxkOwhwEHUpr9Yblgd9W+CcX31RePuXUKtCo9biHPw2bIHBIHOcbxCeO/Dg49XTaVALi
/Xu62LeNi+cTKGWsQLRFeZEUa0WaP5szPINvgjcv56W00qXZPHDHwCUnGaJole9s/9LSBEVoVBFp
OOkPtlWMEGhxILt5aexEYlUSIC12RL840Qv5Mfnrmvw5k1R7Ovso06Wh1d8gNx+yrakC50VF/KSR
2iK2ED0VyFi4K5NYQaBU/JEhEJTGKdh+Qnc37+qRvWBWzjKZesQ9Q5SgCO/hPjySnU4bPWn/9UXo
YIcv85dxd7ki9eZna0zEE4EuzP9mFhspv3iB542e44A/LK03w5kI6eiQvjr445w3EZ13b62sN0PO
SIzSYukWeeNZV+yk0TYXOQtefV4zXB3ob+2cEbavbxaOfLYcMVmZeV7usuMHW8JtlJaQCEcTik5v
FHThHTnAvQSh2KrfCGfLi6gRTpwmdCtHon8ocAAJyHj5QF7EVn11sTgZIxClh3ky1Ril/cXHz5IN
LtnuJyuJ4wvaNX2/TRgkyhNIgnGsgb7Gj/lP6KrCfEI/Ll2skE6y6e+MHjEaAvfjtaYC2/fFceOG
znwnSJJ26W65sfHBz7UTCu79maBqjKiDQUtX4yJiA46TvPPeNvFbkeCmaIAFgBXrg2cmpgrHVPfE
XOC9KTm5TrqWo2Ch6W9BJrUZoSCJauOLuNIz6vyV9UNm5t5of/ty0vqIgT/4uZ3rlqmSOk0ZZ6Qd
bwiFpNEJWTi7tOogipJPgubKtIDo5M3iJUOoBtHWhf6/PdikuUAOHnWnAuYzQG1zS/cNt312e1KL
6vF2ZhsPIHmC1Hy8MRp1ajvKNpAVuzU4EfRq0TJkq5z4Y2if31zbwzOWgaFzNzbTbPbT3RJgCXAN
Rx5hODEDzPL/fv4pdj3Ej/I2q6au7cpnFaOQk8fdL6qwzWTo5H8U7BVU+abU3D2MRE97JmF8WBMD
7h4Q6qkY9kd3OSrFsqlh/fyPIWtX2F3fPm+Zxg6M+YbcuyQ41AKKCx1e5zGdAcD0bd+myAGB5WY4
xRrYk6mHkKRVUEvXOxVVPoEDL+44naAZMhm48Pmc0FQBxxQbWeG1gyajTV0hoiKlXVDSC1nAonqB
SGw/Riwe346eoZcb4l7MSbMNinEjRxc6GJzTyiOkcHc9y8/G0HYZJCb8PW0HWnJ05L9IJbmmDD2a
x3WOVtrmTxR9g1aKfx3ukadL6qr5ZiBp5zZk0Y6ZcsSfccDWKobDT/aKP4hwMmXYwhAvvWk+5bmC
BWliFA+4NMAgbfMthJ0xBjO1dt/7JFtYUfuDvdA147oXEiDBXCN7Ouh/pozcPa+6lGxXOWlIblcr
IyNp2lz+jdbZaHvPHmCYhuyz0MR3uVj0Wa2+RlrnX5CkbjoIJeq86XKkryWd6nQHyOq1UauS85+N
PZHvSki/OHtJdhUKnMxGlw+8nwyJFG32G1QRi2DD65MjZRV5MUdF+jbto/ALicbSKZqKSHY4T3fs
fpNIKriCQ1KQ4vSR4EhX3J3C5HztpcJlD4sUuaMl5YZNAmbZZMcGmQ/1qCCh5M9b9o/joAK7OjID
c6FyzB2mq1FDjf/JEioWfuQv6mPLkya8O5BmKeF+nMTIPz2gFw+IjPFYJx1OsD6OfJHKEBayRU+z
HE1FxvyidrgY2fYR0ztjyv5rDL9p7SdHfwp1pmiwz8X7Vh20SfFzEqpskQaAOpbB/lSOws2KT7gn
uLsYo93wm9g9sNPzECHxBTA7hfOjKkVJJ8RnW4ULCRU7lt67EiW1XB01ljzh2x5uS7vfe09aZEhH
TqU/8+kfEHcghDY9kqNry2knKeB79tf+aQdq9r3Lt/5aHrPMk75DKvIxuc2aoK3VxvT2W2gtX02+
ubmKl6b+vu4k5XNZduRxdzY/bNODZJYIIZ+W2yVmVs1M8k9TdRAfCOaXcxGrPCODNHt8vH1xV+bI
u41HyCyF8PHKRB99MQ0dXhqrWYkOe/F6XU0ugIPIur0jM5mGG/r4mRbVoP0yaSVW+WVkDRcEZoRi
ynhM7xdn0z/aZkjgFWTqgyxEfVRNEvgwxdS1up+As1vP4afwDVzdMldlUprREOiw/ImV5F2/gqAY
Km0kr8yTAddiNNUxCgeWLG6mVpXcf7rnBe9xL83ZQSKxoo896j7Hi9x+KgPJxnni/G+J8kK3GlwY
/pQTQvourw6ohnKhJ1X7ozsbTSXdGqZaLkpdGVsKGB6T378OVU6p96grC81woOjwqB3IMSyrWDoL
+QIZWJMrxJYG+CWcRHerPcBRhk0fzdwb5jSpDHWVrQf5txh4thySrnYqBKWrY1GBmRzj1ANzICHr
cVLEb+sI4KedKZL75c9+OuPeH0S+B3iklzLoj0KntzLKNsYsjTBKDqEjru9uHzcEKioJygsZwJ3F
a0pKoxcifgywNOfgqAogK0f0sHAe4zVof9E0jbGFCV/sA/C8dJxg3OYL2XWPEj1pmjI9MQO2SdbD
vfX8Zo3monlRpHrXIjZUiSpZybF52SGEiUEhP3X0QxwNRkIo+JBYktfgifBnwoUxr4/jT47vm4ka
VzKJBR5lmjBclyDWd/ZbmEwenEekDQgdCI33XCav5pOp1U1qihdsVI9eobu6vt9TWw1d8c4g6qc2
6a3FoNT9J6I+U57uaSqjvcIl0TMkOV9xS3tcYmiUcmd1BuHjw9PpHqV7OJ/sVJLJMfjfXlBTy2Oi
jxsXk1EFlxrChM53Es4CP2hcVmiXuAAGZMfm8VxGIurc5cJ9Pt3gw0ZbQ+LYIfuOijN+3UeIj0Gj
CIO2VtvZsn2tt0unPBDImFGbt1lZSmthzhSPrAEC4fnW/DfvPXU3sIqWGaSAAdZyUDqKZz86lcuS
6u4SCWcUsJkGL6DRqQmkWu62Nx896ovGPEtifWxnerNsTylus+Uf3e2w7qGoPlc6JABRYPypHF7F
zn+w2m3LTYYpmoOT6qmgLmOuzqocoKVHWe2mSDjoMKZIlhMnTOcmmUvL/sy+gps0mEvVyVEyDWVt
9MMUb9slEauRf9a/Zx9kqDkxtnvR/NH4457FYylIn+vTMsd+v0bm/QeC8/Tfvgl25wykoLdJCc8C
wV5I+cebAsz3aVjqsq7yF6OPLfbBLRI2/kTvsAg2IxFQJEhtCAZr0We38rF7F9gjQCd0dw4uCgEZ
Eeqk7NAF7HeksuxpHDqrNI62vkp3P/A6RqbiC2UD1iCTVZIYNgrt5E5NAg5jQXRLhaOHt/MMmDrQ
VHu5Y4ayGy5A0jNLCFp6b9zv8CcapbpSP4pBp2pekVz5EAqT1fD0bS9lmfAJylxOtumdCZnTdnaJ
fgc5F7rjyJVkj+pHGClIGX6213Vu1auW9GB9UD1CzU2dsl8AGJNaPyrkoFQ2beEZiHKJmBIPafKH
wo7ytcMLkc5ygL+IAk+XAR+Ql3OKUCqzbqETq0n/NtGklCc9MJYDx9XSRkJDnx/ipvh3L+1TXq88
bagoItfL88obA2JGiDufJ+MtgAQMxSNMq+S54oL3VkanieG+EwYfuhJGpRhaOdoEnMAAM1mtRtGX
og+P8ic27GoJyyMTcxxyCgbB+MRrgrHLxuI9HXav30PjmBlg1ZOVL7gLTau7RGHt4Hp1MoxqfFzQ
w/DyuNCA59656W3brshredzik3MYjUmTRMx0TOmSxrUzfLGSGC1gclmyGlA2Gx+jxC1+VSBl6WnV
I1UjOWc1D7cHU3+XSpncfp2wJU3AKXTbyQ+bnjQBVYvWIXoMMjdfxjXhJ7pt/YqvfeNDeXYhnCEF
O7YMBy8Toke9swVMnSIZT3FTeJk6v3jQCTSb6BL+RaDd6MbrG9jf0tYV2ku+5HL40Vgalg9Z3AvQ
l6OVS0SS0YMaFTatSgqJmQH/GHLFtYyl1e7dIqXsjYxtTW/kaqkO9zAvnNyaoOgOjidOIUcvktys
itdjkkTZ3+aQ5Fpd0cWHSe2U92fcNQJL9wGaU9FQG2RutBdQyXcjBxX53DqM1P2G2+e4Qec343p8
lSkjBN8WBE3kI2aTnRrVn/Q3pzMm42xAltL/AnCvGiujed9ibg0Ue57QsZvy+9ChKohumFnjrZlX
eJK92/WQ0hK5fFquYIiuusHdxp8fzbE50CmGW//6RpJtHnC2kvTP59wI8iVAKVDc3SAWL+LyNOfV
oB1Ji0i0PxboXx1nYJ8E2NbMTZrxW2w0t9IKuOsJ3G2R2iO7jwQL94iTQvK56yIpPCTGOjyuvAeU
BR35HvB8mfd1y49OE+HxmYFoRuiR+M6+afd/Ifa7mS/KctWhEkowipZEg9fPvs+kRFkkbVlrAc1t
F/h2HVG+YIuQ9MIP7rnnfszzNDQa5aSkhkHjHOJgZmD/Zfhb3FrEhJKV9jqUJQXkhE0LAj8jYz3/
XPairOJ5XM6iy7CrqzpV1ocEf7Vbr7ay/Humm5mtTfcbA8Zd1Gv+QG+v1a2NnlEvs0OH3wNWgMes
IaI50u9WMCSZ4lgZFOZ4Nxz5woOTh6GqJMMKqNAMYYWYJCCFtYPNWrGu0J7h0YTxeAvIH2p3qXik
GHCajtH5B2F9XzrjHOvkbR0P+lapmwDQALxkYOfmsAUHpKlgo4VXAsctATSb3KclGu3fxaxzLnCu
mqrCwio+kavbhEoU+ZZHUsXP4cWbhnaRQkcq2yZrzsbFSf2wfw92r02EY3fWZGPmPJv+uQ3hRj8U
99Zib+E3JpT55+R3iv0tgaYMPn9hjr7J8ZN45O7c+Z2Pj7I0uca5LBZR6Y2vLtEK2R0xqTua8aCE
2ad3/4yt8Mb5Nnk+04UMv4Jto7ZaeB0UWtP5r/2O4pg67BTSmG32F5cg28U/+8qITEvH4iTX9Oeg
zT/ts+9xXCAEY26dJKUwlIbE6pljibZsN2+DJUztAm/ZYnaBmbPOcTvECNL5PIfAD+hy+JLDxjqo
THHyxYUtwDT0dxE5taPVhCgYbqSBYql9xEhzeBQqdgaGNxceRHGSkPBJU4wovIUuM6Bgl+LlUDUj
wXVIOqiLLHjMW5UKZfqYbzY6F6mboyORa2SSra815HtwIwjDIxswkC8fWa2VtRuffYm1W+2LS0Tx
S81Y2sWwcuOnzEws7dTA7K5aVNUyFG6oXCbkKBTDTkoDdWJFzQ/SJlwtPUmzr2KlEvROr5j/A+0z
0HRCEuo9ceNdhjlN450rxjdvYHaOxtn9JjyeJH12pN9JvcNwAaV/iB4O+j/U3DJ818nYfl2GZM1N
RHl5cu5IcygQH//zFrBh8Wk6mlAt3EAxyMRhP7LH/rebOAegDHgu901wPpmRWNNHjIjJw7/Rb0DD
9x9RH2+xFH/A6VxV8ItSs7aJN0veyeVRkGYmSQyoiPrmqPCHHkljClx+aZ92zZjS1uQeFmh7v8ip
oNUeqhncNpk+P11to1bEiwm4VNEXBa5tqwe0X3+K8/hADcVckZxet/nw4CQA0hggJm3GvqtTXzbP
jKlnuU90niXNC8mxrkiO47IOCMXtqTgB4SaxJDYlQZicg4y4NAMSFgggWEJ8XrH+BW4sgh6HcIMq
MZRcWJp16/9wMrIyMj9lJfrcChxpMlFomJnj5pr1n14jaWtgR5rtiIvQBij2SEm5FBzvpsjHV0bY
AUiLZl3m3SfIQlqhheSqPmYuBGRdmj1KReN2VjU50czO9igiL0a08UmVeeZ9j9TxDck/t4jqiGG2
lzjLgS5f04SJtXxs1DFr2q9eOfJZVHWSLypJ07rOR7l2A7cnxh3tGyQXwA8xnqhbaw6pX9Xmz3TY
Gf9RFJP7hUfPSixZdoKdWUj4jwRLjqIYTBppbkgm0N1+kIDjY938/6O6tN2ntv9a7TaOL4qi2t1D
EFiUxrKt71sTr+Pmy1U1jxpk4JYPzvTmvAIwOvDGljvHDe7u1+wZ5L3TXTpoK2FlzZe3aIJb8WUp
n3nmQta5gheyjGJho4msJcjmhS+2kLNWLMGSTmQ5CiKbkP0V6PI3c4Zj/0AAQ/9lq8+ch6RyQ02F
mFmoNQ0hFzuLZMfdkr/s6p3UKxCxbbgAfUdcmDlMjsAkK/Cn8VyWAVBWQ5holOmHwz/p244gAmFp
iPawEuS1TU0Bkr0wLUhYh09SCpSqUnKetL1sz1IaUuhTtmtiWXGZK7gTWVDCBdwD67Lqc4wbh78j
6dZ1qZnEOu/RqmN1szJmzNy7GHphUC2yNKbM9fcAEKox2r0+tD+Usxvq4MUzpF/dEWlypjbeaqdf
zoTqmw8nn8TIuiW+76+89TluW5w1chEGC4A2EnX/WUtgtjA7FbMeimWRO1EOiLipuWYTQRJZz9ZE
JuqzxgiWwGHAKeUvtyFPAKs2YRMwJerorLF3znBq86a5Zx/vpbYPW20n2utvQP2osteDTIdTJb9I
4DA+Cursm9Z+Pf8wCD1vHRgjdg5DwYTWEy5Tu+/1dxvF1V+A0CZnKDj6gSV1Qb+hAZ6WEkscjviw
eDwtLvKgrsNRXz0lcXEFC1soMPvlvZz5fxf81b6aP9dLJXDhC2NqrRiVuhFC4jv3CpAsiQQsNEML
z+Z20879XDGeDWgEUZu3Ufc/jpyoW98V/npKQKKt3VYq1mGEkXIWdEGwK+Toeub/CzpQQw0Yc6ad
Lvtljabd3+TE52DM3frC++UHKgfbzV6QgasFksM3ktYxeIgTWKCfBjE2whQBQaQIKLYelkwUFRDK
PdBwhaCaraRjU0uxzmonMvXcAOxUW/xHfVju+exHABYDhh8Q24QVtO/6JIgpl+biJiaTVB+TCVQs
8QHwFcyC/TksEobBhO5BvYUQg6W/ONrDSztae1izXd2cjW+Rk7vO9i1Rxlp8TVBX1fJQ8YUKcbyS
y+VqiIHII+BlZ1IgTnu6HzPy7iA19O6k02rUlq+7+ai0IYOaF6SCxintPBv7Gjt4RqO9GWSFJ+0i
AAxhIZdhjaFLuK9g0rUTknfGkXAk0+68HGYS6sGm1+A4S6sM6KSQRkfXkuSPNUnhipvu7MvJ2yr5
xdxl5pYE4iGYqiXSgxrCxzPVRy8eW3eUwETClpxX0p+5UNrlYEK49HcX/FnLewTYjnmZo35s7U3Q
Jk/QeVrlxltCPFUFw6a2lZf1MHjGTRw8IFnbOcTDkO4ln7WeEROUjpZb4Ylv8Lu+xRnQOZhnvSFK
yuLCY40s6u+DA8U+pmdGIqpzSDkAuQBJTD4kPG5f28gQEwNJs91zZFEK1sPyCXnUO2hwtGM8uDlp
dJfHd5YjdOXf1Gs6ZKmtWlSk7w4IOhsFyTmx+P0iUmOSDV2AbkT1S1ZJYwYZYaZUT4YjRWVUhBOs
r7bHegIlpE8vLDfWm7FnLLsnR7stsnOOpuKYe+s44WTRBkJpWOtFhUld50/h1iFPf1ndOR7oqVyi
IcQQ412aAoYIgB4O7IYwMGccR+UxN1CgqttMBuvWYgUkGyVCsNTLP3huEUoCzE3/M3635mRIMHUY
x5BSEpqBcR6thGFJoebE6QkegM/DZckPzQgQ/OLEURIOJzZKYQ6TFiP5KaS0Iqvd2D9nElf/DdfO
yPB+HmNXP4y/mHJYh3Emr+uoQM0sYdGbrNBKEGQtoWIbv25198uocXN9w5oO+5A+iJQlFB/gXv6M
YLpTVNR9AtY8vkJQWRBz0F0sFF6feM3BVOuja2eqI9czWCp1ijPODujUEfcJagncrG4lBRNGve3m
6gB0yqDk2BJ4ghGQ0WQP1Nz4LMEyCFHxg0nwO9r5o6+M2sU7MjXvjYuTjM5z4S4sWHnfaU46E78l
STgtU5mBhm7fT2Ycat3M0hjNdHJFQb1O72So+UxDoaH2u0H2LjaLX8NvOvgBTNQSS8sJhAMMpUxO
90pGmEY0I7+7AwCLRfYCkOsPvBZvZmOvfkxZhaREug5dWwoCu0ZdMykeKim93BWomawwqyMjcYYG
RSS/cXflZWmSzdLs1u4u//q50nJeSYcmQFMKRGz3AKWk7cDGlhjbt4IwHEwkyphzJkIoM5vQwkqb
lUfbFRp4QGb/vPbNvl4BDshcuV8uRIUfIiafK7vZ9wCZsSW8ZBuIoLSwawY1gEjq0ws8PR9lf+2w
LnGNxgX7T0grKT5Ggyyqbl7btw3fyeMPqWGXiiwzE3/kIOltkIfdo11hL/fpAJE0zq7e27g9PeC/
7c7ECxMg89vwH06rpPTLQkj+AcqPyBuI8GvY1NnVnFkiFwHO6o5DRxDSLnSWlkzq+i2TuiNOVPf6
3Xuz5kcjl1R/z5Iw6jFfaqt0FgBo1mMvrG3Mc/EvBM32nvdDOLR89FLhGX9UhwX24rHkp1G6WCNY
kLQLiK7XbI6L5YZC4LzPWaYF+l72hflDORvNU+BKiDHf1tqEK/JuEIX1WrgGWWlfPNhjeLuLjgcL
v5Zf1lRr4ix4uFmMrPD9iCnnPejsZbdFd2ggXv07SR7shAFvXfjPFL5CunwY3FOhTtsYFIVX3kZn
4lVSXMG66Bm1iSIu77EYB7NpvcHqAQ5yFk1Bj8m3o4rJH9K9/Fdwtx4fm8dxUyB3cjXBwfc/vWm0
THzb3e0Lb5MHwBys9k5YC+m97AxlUw0uIBRI35tRcR3BKGEQIvwPsJKZv8zUJXJQW1uZwjOdT/ri
XvIJeHCpKLzA/nHNcV5xuG63dJiFehWfPrvvVEKWMSIUeK3t/a2FK10su08t2qtenTLRgH9uivtM
35Z1lFddHGMpc6IRiQEEmeyb15gtJyIbX6g3BofQXgp+7iuhaTw/9Dr0BD6ksq+nkUw6zvRoi02J
tUCJOuPIYFlQCvu+pIB/tx1G5+fC4Sdk/d1aXqLh98XL8WNQPFbEBmhu9op+x2KGKd3sp58eU7F4
wKz4vVF4Nu+bpD7q4rQn1qD5tkQ4i5O1eZL3f/MsaKyNVsAJH/autIVMwDUCB5nP70CZkVZB7nzh
n3PMvseMJEXIEPEgv40bPeq/4HUqMtvTp+Kb+I0iH2/Z91V5dzZmPQn4FfGTi8s4IlQnrxKj26eU
JehD6Q16NHXEf3masfYX30RBeDJ7hGVJIymoOsCKBGcyuCAC9Q59EbxYhbczsgDWFS0ZeQ3eeMhm
CAB2gKkS4GwCRBGYo3KzPZrbBZEOGu6MNDXEqXBWw632SqDz5qZWT1a1+P8VwNz7bCNPQvm0c6Kc
x/kqGvmNSd/Wan11YQrbnIo3gZWhwPuzWmKWO1HeiVuBKJONflL953STMiUc4NtQ93gPiIBiMTaZ
SuOSN2tLWjnvDM+VNMDI/HKp/hF4+zuvy6zrzCQvXEybeR10lzf9eYbQm5yl/9NvGCLWjv/c6k6D
S6+p8HRsLfXnPR5LTplhBc7UbaS8Zzsooj5RyMXCOeK1aWOW6q0M4ER3JdGBb9eYUzDlcGUrhlx5
/hId4idVVkePx5Iu9eI72FyCI76v4ODOyAJTcILuSisZFrDzZtfdmIxFr6/d7EfuaTc70oQb2G/S
WCA95Nz2UUaoJmkflrOVoN5T2bLZ2OJLylO7LCqj9Wq0HZMOKrJN+QRoLderYj8JC22WWMOuO16F
2ulRDN5ewbzmkZZxZOL89sKhb41MugSUAyn59+BQbQAF5hUAF+c/CYLpBQDSCu0TtysUPtKcXrgO
NpRzQf5G+0l+CdKN9ISiMeW/ihhapqwvDvzF8YVLEyol/eatn6RDRaztWthHHB4HWxH+PUN2/+ae
4pw056D/n2FiX/pGcrIzIf/OUKbeR8/LA7bFh/zdhTvIgZfFHA5wvYd+H/1rZS6l3u+cu0IkLaa/
Ppi55fNK466GPXBZiuBzw+r23zcCry1XeYzpAYNtvwDwyjEqfJVRaWJ5RbpZ4/dptN2Wh+Rz9gDC
rCmVd4CA5P+/9B/PrmkYWEbkIQTn2zJKILNeJlAF8t2YablNI5TX5Nr0907FEKi0tsyxZdME5iIm
/LUWt9JMq+2h/In3IlPbd6EGzlyR2pIvfpv2AY6ToJYu1stoaE3bbSQPZyTM9Cz55+DQv1qvRz+4
wTAQ4rVf+p/WIlEOaKlpH15nBuY8Hpeyqc8uZUxYikX2ZHdfbnS31T0crdN9kjK8QIDF5jyKdVBo
5MnPYBx2UTAN9+ItrlM/9slpZUHGj1gyvhvkwDJ00hsL4oltrNJHofgL1x0ze7gtpfCK/B6/SX+E
nyBfDoRkpgOCkvz7IYMhuftwUhCmRgE3d+fyt9gokanCgV5H7PBWb7ho/UsUZkCEHqEzuwrodGAe
gxAtcDhmNUsHUlsaUIdzpt5XUstjwMsqtMvHS6ggU4jpbKBBN8BX3/CRv/HEa9czHf4Z20r57DWa
SxJnoEunROvL8jLG3gfFgccS+ElgfYSlgj34qOYz7VogKbU+tb9De+5ug+imLZlDMBXExJuji3/y
w6JIikCLsth4414xAK9af0coHTNOt98hXpeI9jCMCDMqMqW4M5JtC6ufA6se65cG9VbG//JfQfdZ
7gG14bXz1AcnrtfTTXWbByA3vsKbJWiM/rqV2yTu8u/kXbNtV6cWYvdLdTqrpdF+RMlC27x8lK5I
uQCdVKFAS0wNIq4BADMBfZnLmsalDRPIgracUfql7RHmTjzhWfw2xlQR/Ez+oBElRSS2KpOnuul7
8n2yz9JsG9n5fanHiiHgJPbtuCKJ6drNu2+Hl0S+TgK+LRY6GF3eole/f3H30/gNeW2BL+qLs7cc
2fiybISQmf4XSj4/k21NUgNACXhNJiz4oxFs0wbuiP9O7q+zgMing9miBKJ/0wXDl9FSGUBlbiVr
doEWNSa5uKQwWVgZHYJxITmKktaVsIjvNOnjr5qdtXHYTADB4GxXkNVgvDZi14UZ5vXjp4wKEz6d
X4fyLgcBNSOLe1vY8yegF3cchg0HJAGbl7b9gNjPYL37OiWClaCIrH8KioRcSM8Bga3O2vdYdUhh
LDfMOq5TBgcf4gasNx1yKCAx2D1xA7UQ1FrOzwT+B8G78A1h1kp7ttIJedRqdprZn+N9n7BDPzrp
4Z4PdDEpjNgBHZ3wD/mJLy2+VUP6HiDszOwJNbjApIG7e3tluKlxof4HuVSFHL06zdykgfMPIYFc
mUFKCkueVeZNXv35DcBj4j2RLUtyoo/bPPnKQNi66hnfJAv3c/Ag1/TR7v0e9FwMe/OebrxET1oM
pFktZPjPv/A8z2cmOolPG2jr2IFeQYnJ6eG+rbKl8/A4qbOHX3WPCB04MdvOyd91zLNeO5mtKMzJ
AzdlkBx2D0dnApz7tMWNoaEuSsWnTu1bIShztnelSUZygQmjDLHkq14NDbLz8hdW/QuBQ0Q4THAa
Vkso7cnGzQSF0+f26gqQZymp2bv7CyipKVIKeDrw7DviWvFW8lyB3OZ5zIQfyjqI3OCPu20qVBUo
it1vhf1WEfzqf7LZRGfrAhV4yKSxQEsIUdIN4JKycL57SSsf8oa3ICtaSLdXl1jUZQ11tI2YzIaa
eN3lXkRvF2UIk445EjWINVYv7SzjEOitNv5qWB/YhoetCapCjKwXdjqQNtdazEpnvWGD3f07ZMTM
zIZkSbY7E7TXEHz66M//k10CGIL+4sP0HT8K4dEmpaRx0M3pVs124BrZAxr57yS5wcruas0B2Z2Y
b9BBIk5ma+ZpeSV83qNoZpGfteEh07C9lzBH0UykVlgPT9IqgD2VJTXqENh9nVPCUsyg4bhRPuip
oBV7QvcMBlYnqkvVTdoHKtz5p1OGU9qhsHysnOYKxzY6/yv+VdvRPiZZs5RPQRERSk0rEnxUDBKg
7r/1KJQGhseusiz9vCBuKz45l0QYW3ww72Nt4HDUTNpVVvyKtEKc5ywn9d474FdtaxSSBPGiySvh
a4bAlX77SmUo6phySn3Xm1k7pseg03jFkNOA3ZBk/8XId2PHNk6Gi67+JQDdXuTvkQNDTO4a1CfH
pAWSrkhW6TR6dpLkoGTJRg2TAkEw/EzDjp5fr7sGfm5rTFrVp7uFj2RDTIyWNn60wcA/oxhfnl6a
5V25sgv/3aBi+X9sEj3M0X8ZC1L9PPUmw362HOn3MLgaLCBLUFvIpQs4GPM/UhezeDx7vOXyMvC+
h0ce/70V5SB3ASM8otUIapYlJuA9ZtkHJpMh7VTzdq3OosK2QlM5jkYyrRHKP64W+f9Ut+NdyTrl
P035yvNhLqnJtZB0fcU+4fwvHfDirWJ/L71NcSDTnx/pdRThPK/PSI2P/P9dAohldIwxPx6zA+FS
R5ZmoU0E6Mr1l8FnlZDXNUyjBPbhdfiiBnxI1190f/edfItIIhM7Sg/Nlcd0q+KxaVAHZkm0kl5p
cNnM0ZSrzqmTT6kgWBHegh5JUDy6W4lbNmVaXCbQ28pLmPAdrv0SJ6tmkVIcyhOwWLw2pnLivt2a
JOiwnxoWvU0SgnEO4yVOxbhlyMmcnMYXEu5lsvYbqAz0vbckNMcLhz42p4tH+TOk5ULrgOB9Anvd
9rcYbO+UBWb8t07TvT1ladVQjSHhfIaqXxvZSb/dI6lguIExkw3fwutcvQ3wVJrkcvZCefVTZA5r
iormcPBzscodpRazX5Popy/XWSRMRFA0wAXpgu8Jmu7twuHHjbuEBlUP35+8J8fue3pNfc/Q1jpZ
4YguHAD3c8DfK/9TYu0CZgO4S9AKDmNg57EwA/rYJfNSp5cB4oObPJ5jmgrTcQngsi7U7P2WJ66K
MKehj2eTINlfkgDOOzLXllaJIyrlDk4KulZgqo32myT7bPxd2FM3oeapmpAK81ox9AOOIjrY3o6I
Fy+0IOOJUZkI9ZoTh90s6zvRKhetlhfXKv3fCuGxQf4Hikxzev132SpcmC2yid+MtzS/KryepSU1
4WLksXrTnimhOzwVWFUqEmPshcij4Q5X+V5210xq2mniXuMrGU9lLjWoT0eI/H2JHKlP3Gjw4UWf
IsMJzdNmsAqfuHYYVxQakohRPpch19o8GqXkB+Tcm1KmvvsvjfVNs0ej+P24uBPPXbS/HTq2PJvR
1dXRxUTdoEhsl3PSxI/sexaFryR1a6NWlGCqa78Fl4JY4KFxa/XRv/sZIxVFlcD+niy6A0xjp0Is
di0WV7p1h7cKUwawZyionCZzSMVjy7ut3kTYZPboBYufzz3aN94+rvzP+J3kBq4tO0EohSyW/rBc
Jue1L2Sv56mVqyipO3Eyet9TQ10zSOB8T2oJXNWKzgAdWkfEdN3U0KJ+1sWygSyk3naY4e/xKl98
4wnNcPhDmTgACIK10x+yOjMXPCQdfA57BrGzOYF/nMBomPHn3d6O16Qa4Tv2YfSR4zzl66AoFXy0
Ev2cLpy6cbMLzAHjA9w1VvyBwDe6/3mazVHTaCebduyRVsc6d9Ext2wx2GVICEAkj+O6I3wHeF7g
moTdlYxblxm1LeATKFVBCIa+2avYrACqSkU1foQNY3WjPROozxD3vRQkQXZvHwW3XiM+B4Abj9fO
FDE8qRTsz+mdKP/DduZreee/jSkkQK/IeHVfsHVmi9Az/Sli2n5Eju9wMIvPd+v6wMT5qshbN3Lc
sIvblaslFM5DGcMuCovASGD91Rhz9Rm/GyLRKBxTny13wd5i6I8iUAuoNiHKdJctA3TZU3JmS0Iy
j3KyFK8Iee6ZgaFiiXX+hQT60t1nV2482Nny50NEk0Zt5ldDugC0Vc8qr/fSHhZyU3cjyWNBjb3+
Gxu02ZuC6SUAukq6QfqxvwgW0nDFVepylSk9nwbBKrE+eUbfnrhyJpS/sSsvEgLSU1QXUKxiXQRW
tYbiWi0YkMGHiQvDYcQDFxhmzzFjEsMUaFgcXxBvScfr6TXG17ExW9ikNBFAO6Ji/w5yvRAkrOEu
kqXGiq+3em4802ToGWe1mbDiCCud7noGQLDGixvoPMQr314RkgtDFDx5emyW8eyOa3eauHmaZ65V
eNP1bcdMwwzcgt1qRDkl7MdcATj+T82HFKq9rHyR4DS5+o0iHBtXzVosqURlwNlnnOSw178ml88r
6QR3ELASKUhGkJQfXsmP/aPk/D1A+eR8TMDHvQR+E5vkuoqUgLXs5YkWVlQdD7BrffgSa3ZBlaYw
4JgcJze3SdMjXrlGIjaAatrt+jcp60/+ipBgGaYF21YtxDe7IMo2AeXyYehy4awibcm1V6Q316Lj
DqEVx/mtqHrfBVFgxOzkPxk2I1LYnj4shsoSt9fatU+qcjX7kox25i2Xqey9NR5XSd0ze35IUn30
w1DRr//9hTe805/QxKrLP4WXLuK0GO3t3uewBLAODu5zkWhgOAHWGBTb69k0IPsya77vl/YOVZAf
ZYHBnYnsTS4zlfEZZTVVA8cEzKnZM1MKr6Z6Xt8wEPNZ1BBFV9r9fsiBdFc1Nh/wFZutAj+K8E8z
++eSnR2pk1O2dzgOAQplZEA6C/qG9uDwd0a/6qaBG6DewGdhaQUa+8J6GW7dy2m3VDXXfABKQPIJ
J8IcBOj0ltCkzrgEYqY3bqAFwo+wt8K09RN01fLeJZOZZVWP2ipUUg8da0RYIqyfSS6nD/gaEMPv
CjtGl8+KyllCcxrqdZCRP3Ie5BJUldXJyJMVnz7lpJL5ou9ouDEpXsZiaQLp+HeD1T76ejLVMcrX
ZjpTVpIt73QT4IHvSYj9FpLfXos3Rd52QtPt1iWjpnCT73pAMncEw4TmKRkCna3WfG99V7HlHPF/
uky4hKRNoduFh4KL8vpc6JqF3ZwAIbLyLSJTbVD2y8O9S8kCrRleM176I5weO5GeNbS/lYBLtesz
yKQS6ljyqSbzY3QL2MN7xXvpYa1HaoJV9lOkJcaRQziu3hSUf+mQ1NFd1ejh8lM674WwPZEXntqS
IWqyqnbnVTtlI+QaUV4nbQVjANQF0qbgNizaeWEn643mzXV46gS3c9AsRxeIfbuuMyp6XN3ciRhm
K+uuD5rYJv6G4yPwARpZal8m4vgUj6X7oS+wSwdbOoF3oxmMYZ1hpwL6w5CNWeEZgDGt7M8mwtcg
lotHlRIdbnb1wRI1VPVbhysQa7Rly8R70VtbarX0+Eg+kEoaSOVb4+f0r5BLqQNSJJq3btLMTEmP
+J+9IM3vlrGE/d7uTVJbXJL5Y/mbIzcDh3R+nGSrUC8WrJu3cK9swF+EKzLr4tfyQJ4jEpmOz5Dg
bxkXo1pEZHb7CpelxLBGaoecbTyPBlZ6zfEvK12vnjcmxfvGtEO3vcW8TpK4MvZn9FObHrAyvfpU
k0BMpBBTqoVtWLg7IkGa5WPWapOhuKpHIz3mLKhbjzLLh3f3YqdWhlMLBbNUu+2OxapXCcAeIJbE
gJqKMlKqBeCRpBxtDzY4S064w6mRKsRrX1DV0GEpYZLX2/Qv7u7ojop1hAPyBOVEywsy1NyYpk3e
xK/GSf8cPx4Q02Y1G0bV0Akc2aFIabxKeBCH2XLYMz7F7KmXLrw2ihlFMjw/HpmQtqDxTy99V0hN
7AvbR/tIdYZZ2KLiid5vhUYr+VXH8Sv28Lpj631PDuF7a2Zyz8GWQ4v0vu3IU2FNDFCumyCCBpeg
JDI9P2jqo45LlYm5LgOtyNz46vM0hDJr22E67qO/tuAM0rgIxuKTUtBJwUHdHG7GisLU62pQEFGR
3hTat4qV/e2+4vWvdkNH2v/RN+ZwYh/vHzztWCvP3/O3jaPWjaDbuX2l4ZFzIHoQ6WSbjYdW+8Lz
MYGVYSFfK0WOInWitCo5j5Ibji81jJnFkSGRLv77B4kWyLsbtHZ9Oc+YHVBCbOj+CKQFJMr9tCPt
XCaH3XHBlOMPSJnz1BynoIJHiwLEDwuuLLbtiufC+ng7f/PhJuAgpb85kS5DTFjZyDSPtTCxSicK
2nLQv7DFXpxXgvfsROvLpxM2G5toRWSsXueHiE6W5r4NqiUvXFIDTkJ754u2kEEj6joNFOzZrIUl
Q/Cic4H2oKVrTzEFAlwb011CI5TdBTXaC8niYMOip60Yca0/5K5tYCYmLkjRRqfj8I74ufLqUsAq
uQSxg44zsCP/30g3n60WfnC/6LLUXl7bua+3gIiCSowli6fH1QO3soG1v0U0h+YfNlRlNDPu5yeI
27nGkKyVCqA7iB+JHYD9Yu8Ii/2k2+xHDmnaJ4rQ1tkwZkRLACOUIZ9rSk36rWVclinezU8wHuBI
ycEA3QjV03uVy2zVCgoriSf+qViIC3ZQgcV6ofjopZyJxx8dCfZZmxhkEKDiUtdNChSF1Rv5siRx
x4DDXXWx0AStuRTJFDCapMv7bwx/8w2YC1GAbl/cj7yXrPUj92Ri7VzzufjGzaWAZdeNI4SIXA5Q
nrf0jSlLIdK5hLCVN6E569BuvJ58Fke6SgxuG5XBA/foNO0bF/8CpkIPht6hycZhZ5DnQIO5C0Gl
KZcd88mz7BfKnu16RYm5zA72PQmMSaoI5MaIiB2PKhEM3jztIjs//Qps6bVaGwYpjyieWYYzac0o
TygjtFyyBCfWXikymdwqQiO3Wj2rDTe1N6HVLYkV8ySTGHmvcQ8G4L7cWmWCDj/HXo2cZWF8Kknt
R7vBVLgi8WJ91tdQWY0Cg6K5SlVG3Bzx/FK1lrYncDc1HAZg3EwNd+pqhaupFWVVBXW86fCYW2/7
DogT3Exq+7AMzKh8oTxw7T6oqFAivRz3S1Qz3n4hy7tBXX9sS47jGSAoxHzlY/hik1cxC2hhcMmK
B9OjCyvyvpunXpRxD9oAuaxis7Xy/TxmEmPNxXIO7iKWWvhfcmzXf2ReThh8AydUgdaBGA1ZS3ov
X9AbAptIKv25hMRA47qgFp2Weor+cjMxxObUq6a35Frrsq/XAqP4FKKhzIxNUaHhN8BmHRwlDiGL
B4PhOS2qkxipEBp/pnKaRFXGvILQv2GC5oga1hAAUX6MrR5zgjJMjEwptL4x+b4HcFdHoN7G/BU9
OEXRhYARxHX1mwYZR8y5t1JkFc1ElyD5UKA3soWoU90DPFId5RYES/xrjlEPff512gnUYbGp81ly
wS6W2RDujB3vx4quJ8xSoBDHrI0rUrkEXyC3w/A7pTfYELaC1LN7XeLlTAE95rl6odZp0+Ubv5Ij
gx3ZrCCbAkol8KI+qFrwMT6OVhI7BchE+lARQxebfmVth260KxkaIC1bfY2pjIJhhb4fVjEh9B3y
BrAqoy62OQ9F54NLy8tgX7TCnKrlQMVdztj/pZiQVwQhRDxFWNpovCEAlsqMvMQaF8RU2RUQHNW/
heaqH/wQKvb3+dMmRwmkNksK15OJScwZ14qKReVN8QWgU6oOdLmc4Togi+omfpV/yQMKwka/tfpN
7Yhs6/kbRUk+Xg3XWpfyQ+HeOIbefF6XEzJBNYI/T+4HLtFk3ORH8TFeFDGAkrtwMZ54txRzXSru
vswuQETjBDlfU7lZqI/Qnrm5o9616aWrOw9mVFdZ3o3dWNu3FgYbbCF0KPjzBrmLaE2ScDodPibF
F0J7LynWp0diUbgDHig3kxmmXrMVDYL+79foL/VnylMT16E3tLcmoame/t3y2v3Qyho+Upi8jNJR
hqCIroO0bNoq1LHsaOe2YtN23UvPTiT4n4IqQ7nv8waa0IK1DL2cRWZuQNPGkyHkpILTzbINqLT7
mabBeWPXRsaFSYPgchpF4ZNfIu+RQhPvq8GtKfqAvZ4vQvBpb1ZdDTk6WD4sm7INDgiUWHqWllDj
uCZCZGYytWPk/yg3yeRF+ishT5tXMEqjBIZtsqB8tC616VGa02TorVBWUruOE/APtSEMZPM5nhef
L96XbmyJbY7XFFTl/cvXAgDjVWUVVR21p+GkM3KF/RgGpdDJ16gVTyK/u0dSHO+Qc2FfAFrb8OYx
sSKuZR9Gn2e1nprkMohOA52hchlxmmOm6QJ1Pl6qcDZaJYAa1YyfZT8lzUe+tSPG6vxBFXO9nAm4
gaYg7+ZBMH7O6/TMqboD2If8NWHYEhWJpL5jfWpmYenC0Iq9FoMkjas0TUOooLAgWLsxUbRpEPta
W8oCs/3pq+f5dO9/I4zCKKFvp9yWc2yMg0TCY1yiqsGq8mCbuYW8Lk2qOBarssJ9q/hoT//ON7UI
z8Znfa/lZ975ISqY2yttnIbc/zBfhHhZfyB9l005K11tLWuZhzL9lz2YVZ3pJ70v3Xx8gevnuD2z
vPBy53Y4lrnijCNA+UO2oLwbTPPf9eRADq0EYqLuhvon8S4ePX2pLIQ1zfRfkYht8x9MpeVKqpnA
XSnP6xNYTHPeawvZ1EdbnZkHAdLwS84EPmW9Fpa3ICVPdSMFwvRdL3qVxA5/pzYYcD/AolTTVe9f
eAByyJJkrgic8m/hGdbWoQ6eE3ROsfKOxhoJjfB11HRIJRwHDRCJwe4ki+psx+THmYrJlJcOn0lB
nioBCK17jjc3oo6nVssFqufQAP6JL9zhGATwkQKnQakGCwZzGCjsdOTUnlmtqNvmFlfKPG4pMCmF
bhT+eNmeywgxoZTYVp3HJmIMSuLIR328ZyWI6X7SRf8pOiHrhsmkzq9l9+ficpStuMhln7IJCl7q
+89tHg35Q8w4qBu+kd0SawO3eEYhkttSG7lZTxD9hFBWI2cf7k5sGihUb8skrqUPsDE+iS0fG9QH
6mFQxEuOgGmG5LpUcOoWlOs8pmTx2M9INMhigs6fqEIA2nYZwWlzrzYLRfxAcysj9n4eq6+XOhfL
hhmhZxQ67f2CeH50WZhCv1WRU3l2wM/aY6pI+206xArdp4MlHXtfvlyhnyj2fmS8iYN8fBFxohkY
dND/sRP6eLd2QpBMsRwB8gws/glNTkf47OpV5+DZunV6KpoFm4UCvtzJHKGYzRg+rLyzT2N779i6
y+Ensk6EfSqiiMD1eRMGfc/KZujzvWk639Q396AayhwAi9orzhsfmP1LQsnE4P07VknSR0H72a3m
VwDW+bLHg+lFVt2s2ZSFraIPseqJ5WPoKrqFG2ayKqx2h0rqXxPKabcYq/+9OdswIjJgaFLHgV0r
z6Kwv2lg/JKSg3Oe/VVBl6PTZIueUyJINKZypHwOIahsdanm8cxP3kcEb0spe+GtUp5JyO+W3rva
xN6HfXNaWyEmM/B8vBN2U2tWOGw1VVHfFMWe/E6pky5Uq/woaWylz7BctgczZh3MSGatSgf6Q0ON
ARtxiXIu1kFYV9pa4qWLM3sSi2JLr6bs3w+duVsmDODGQqCmTIx52jnHg7CcvoK5HFbD0j7XxDv7
lP7JmKRGgng4mCha5oNB7NMSCHwjs+sAYBX78yh7e6qMMVrB+huaWgRCdWPriFac6zkZwIQ3kfGK
2jSS4iOC3ltgcpXHq0rdgcnV9QbEqnXctS+OqjW5xR9xl/hScQA44ADU8UvZR6/It3imXsuWRI5w
WIxhD2GSB66/1TGcEZkZ/Rz/lLa7mOyojWNSAbQV+qNsFR4hggcMEgxZX/eXppOe/lMKWKyMdzfu
3lG84lUzpxc/fO0dxMAgJV9HLGSVldGb/RQyWSaVK367ZvvlmB361E2f2KqAmG/u4+fJ8Ej94IHW
co0DgQcWJ6ON+9pRaMqftVmhCKPi0IvTcaikHA7YZQMUtw0cUpOF6TrtrUvaYoD7S4Hk05TmIVld
693GLAee2z1fJ1WYhFqP2raOvidCDPQqswyyDKlDIESygpADTKFAjWBgfjEPz673b+UqOKnGJVfa
kdBbumpHyHWYaO7tSnZvWoXBdhax9Xj0oHqprt3N74YARjKgkQppTZsesHNCY3s6R6vZMTNaLn4W
k3J9vvbh4KrhHLEWVzdL4hcSC/dBMZ0DfIKa663AWMgLaQ9NMBl0zE+U4d+2I9masLdzKKKm5OK8
LG78T1eC4Ey8loSjo94T467EzKCH+ydjGzQa/uOSpnDWoJKsFTUxE1aT5LNrxuL9s9lQHu0p+yni
yW1UJax1+mSxvak4LvigJYaLPF97RUrdXRQ1QENbJZ0H6I3aGGAd79iM5AyuRj54MHWIIQh9XviM
eYdevuIJFOrfIZVwKiusFbHOOpeZzA0eoxhf0kNu/d9hqRc+MWASzoEVdZwnYVb6DBbLMnCq8wtB
uIRywdToXDBj31g+ckyWtagaKCL79xXML2l0IVKJVyoDiViPUutuoJQobDNO6+6gjezk2/pj573w
xnEPw0QJ/iNTIGgFQXuFDaLopWSs8FkvIx+EkOUXHBPajfEFe0szwayX5K39eSteLa+zZ3BWeM+v
z36LDQ7DoWucRb5BM/0T+Yi7wCo3713pzZZ5OyxWA6WUoRLGdbyJZmvkOb1R5MOgxyQkBbDxmFhI
IFk5rM22SdnfWjXauJR+2a5uWIXt2xbEouBkr35T009kSELri3dnMT3r8UCx2eJju6t5wQRSUoHX
oQqYP0EhOWb3sjCsMr0IYcYgjeQsLNuSrb/9T8kdbaxSrfUk6xlVpWRrva+7oNhvks6LInYKGJ/f
hP1SBEA8QI+kJB+DX+GqtLTlLXkLDkjS+LHRcoivvUNTO6wIuEAXvOTF6HRxWPR57kKGu8M5T3cQ
Eaw7xYpQl+W1X4Tq+9gc+Lfgc42oeGkgCsY0HkvGp/F3/3LK1nur3iGbVPPQX+ryWXS+U9OM4640
XO0z1mVbsGZfT3cYxPvwD+K93bhXAET3Tfdkk8zJbwuux2W9BEMNVurV3PUVMQjY/wwMHjdoiLXW
EIAiPWka3JXGGvv153Xu+0WqodYG30a41fYjWydJqgpcIvfDUB09jqsGYQcXvu/Iv1bIzbcosbcL
jdvQwuNLfWkjlaUHtfqMPlMzEKn8PCfQCUJzrl4dF41ZV3+j1hN2fQ/FqDHWWqWayA2iBwoagp7b
HvrBXxtBbP9zKoGTqFvMaUameLro6UoGFCJZrfoRrTDDdEjuwJY59ECd0YzTWaE4oLF8t7oaY63i
m0lMIeHlqHOGsFYTdqo8Ezng3FG0BX1CdFM2CjzhUGykcEYJ+1fTJbSrc3N9MANHV1BSJZmdrQtj
uvAr+HxrJWXJSPbioCMhgNjpZlr/9N1u/5e0WdAePHtb8WOT8z2OwqcZZMnkwh32jUomzZjhAR8c
jUuS9mPe+akj0k8CJVIqr9A0GVsIRxpMSeKSp+CF6CCqbvbBCgNpokLiZUO/HAnAUcYOPgdOtfOb
4KYTiOOZzu3XdUKBxeU6ik0BAymDkAmQR1mVl2pDXurtbkkl9B3ACMwikPv/ivv+zI4NI4EVOuvm
MFmtnhGni0G329NLz3Ez65o6FOBARwz9RiWv3Wdss0EhCaCi30M2RoQ8WjJZ9CtYOLl7IovHG+ld
DRqFklkmDtIDj1UO47jD7I5lPUnIxrzztK/ThfSd7OeWhHzUaMKpkpxvLxUnC0rs6bOyK3CmW5qW
KSVWrWXTuuRxh5uwa99G99v73wN8Gy4a9FZoeiB6IFDjgrL7hfnnV4cIzZCQSqaEw4wQBB9mDM1u
he0lh9qvBeC0IMVLU5EsLmdevEZ+5a+Zta3WVBzrZXasioWQNhWCAYznBOhSXqmp45WfGUhA5Ru6
g/y5yZJmxkw5kqwfxy2a/P9fm2FZFpX36ig0Bm0DKiw0h7LBGyBe6bSUiypGmaK1NiFBEsGq0ch/
a0KC66jJU/Mmzc0f56A7Bk+MCUaSLLIFlzczuy0bcr+MO+lKB45HB7s0HOcWRRLHYlezC4AVsU55
Qg+whF0wPvWjKuFQiLkDUirz+me0tojDjy4slT3+urS/TdN04zvnppPZkm+E+Jf2huS2EW8zroxD
65lsOtDHv8XRTqJX+TUFFWabQW8OKfePmOhT3UjrRGMlOAQdvjIjPFNBzzSQmOwTw1tO4sTZ/snS
Pm2PrIEqc/ZRTx9ImtfhuymCXJTAmXudb6qA4GCN+bdUEXFPHBBFs2DYWR5DF2iE22JRZVs3kY3R
18Bs1E6x9ao9sy+BELJ80YT20/La4KZ90X3y/sjVPIy1dnctwR1gYVvN6U3r/h+aPS/qOGV9DH7/
312bDcBa8wcV8nJL67XqwD6NDOSmz71aQEY/ha1GI9FracT1E+KQNTC0bJsxXHl9HKBCXRciIzrQ
exH2i1RTodl15D4TwD/B5oUPKipO0OVKy4x3F9bC4bKU5MOqgDZmmlCazXTzxPMo2KH4p6+7sr7c
x2DSxj5C53jPHdbg2lU6QdGchbMlnnpzP7jEjy/EHoSyLNlLK6OK+C04HmZvs97oTpE4TBe+Bw58
MMwFMIRLtYbKPIp80gy5xjZDEMnpT2IMdn3Pt2kJ/l8cqFIDkUOoBugdHUmyKLy00RZyIZIENxfi
sgzbpXaH895kk50+XjWjvr6CXA6r4l8s6NPfGc7Ic4taGZKhhAfKAfsbopb1zneRxSo6PG8b+UcS
knAcxB8xmDJ/sqTId8epcGHlznKyOkEXAbNj9cEOgI0AiCIbP9jLotD1mqLQJmbEKayl5apByBKH
v7SC0gMGsaoEczMM97//hs40Qn8hgmwkIXtPOvwSaMCXuJxrKAP1dYEZcM22w5apEp711gp7DuFC
uJuSLBTtJY40wLLuU363Fx+hbAHrCvPmiduPILK/ZyRvpBtUF/uKHVnh2SNP9rdn1zFkjwxMispH
A2ocHN4qXEE4ksS01tF3D6JkeW9yvD2ZdCucPMmzRXsXSNgqoC6hhXNeGkna2H1NmpSne3uzoZ1y
aC0uKZTkEXLR6uEx8krgkZ+Nka9o4Nbm+TSphOguPSTmypVh/vtk67r97VuzPtT//XN/DcK87TT/
Fr9uirMbL7zmrh0wo3MEa1C9VrbT0aiSFruMeju3E+u/nFmTVYFEWWTVK7gaCwIduioEPH918dnz
OLtEyU4Awb15QMI44BNRMzqd1EgIhLj4UqOFmTDQxX7zIXnWK9Pim6WJHLQSClmoArS0ju3+S1gG
JZw8P8xXFuu6S+NZDeU3cbq7CdMnd9F+J6/Qd/Leznaa0dXh9b2mJeIHncp/ZvMkR/jVRYNwmXo/
s9NXbhaheQpnL7ALjz5u82Hurs61DRcngNuYt4jRryJ7aMagAdHwDvWA7UBLXJhJgLRzq5XAiCat
MMCnQ7aQGMbVPa42HxFADRTLf8yCXVnhW9dPmd57ixFydZ9IIUgOEM91p0HLLpAtf3yQhSmFT9AC
bhUdn7HpxwMwQdDDyiXutlxvDMfsBS0AQb3f3JYvocx58q2iNh8akPvE1spm2q8GerNg6FOlO8np
aa8f3yDo6xXpGLPh7lFGKyVkRfTfVTSvP0f2p8SM/CtIh9xo1ToDr6jPUY4M2sizKHPzCRXOoeFE
DyxafI0nQ1g2m9VkIVXWhmuks2tJRvtb6/mZxcjN+dY8ua8XhQtxxbXrFD+kY0jbPK4+xUS6ujGg
FAuASis9wyqTEn9JjTg41mtjdB+PdVWaoQDEw2ATuD4wl3nsEroAqMyk7DdUyc7ebv8f+ebR/c+y
izJcsHO2YCwSeslfbmqyzW90REWKglkXV2a7KBfeG8Xm7OLW93j7GwbvQYXl0by+Lq4UIga4MD4m
iO3Xbd53BOng9uHgwdU+goHmKvOPcQkkWucIZBzcUsC9vHtyoLaay27mGVk6u4Wxyd+zJ9TdivPG
R4qCqw49g6FA5+QlNUsohGyaNETZlN2MYNq+lGnImrkztD668H0GGGZcLN+w9GqOzd6QReF0bozr
AxfFplUlDZ8IU3sUwQbnlAk0KMpdWopn2zIaRquApTifvPpSgO0CSwH/bwCJs8hI31Jpk3CoUCni
Ex0rHJpJRuViORPs1jajRVMByEY3wJwUBbcBxgJpf4BNJTPRaWQtdwaAKv+AonAH9WNJ0tERB8GP
X1PA4H7RDfvLXM8NJ29gFwjcDmRk/MJ6iXkZ/Tw6LFKKttnJNAHG+zDYnNFxrJjXqf7MDICZeHbi
1ehapSJHUiOSRYkfY8HuyF4YZU66KMqiWeLBJXkTql35aSQAL37WY+9d+bHHs07LgvTU0HzuBoiW
seCYDQi5qAETMs/qcw7izDiSkQWik0LHrBQYmRPBIT4QtreZMaH1Hn8CIxjrjk/BaMa9ES0AanaO
iTc1h9P9jMZHT35GLrSdstg9BAo3cIVNtsSzansS6EK0akO3sOi+kNej+YmrBNjQj/OJH7mt7f8z
s10ybD1TiatLJyO37XG8HGcMiqlYmaxtKExHNSruPCG853f9iZ+D23811SHOKeiXmgaqQQ82ImGm
zDpSMxr2GTlMcF5CgJE6Qtr8xvQ4QIJyJB/n1VgMTQ+py8nYUhG2q6y0z3/NfTvUVqo9aJLLnmlv
gtXVZIGvQbsQKY1Q8avkeY9/TSYNO8KtqlAELoX8qOsIAx3VhPPYtYovx2iKpso+u3sCGrRyhNsm
XMmu9s0UUuFqdsNRHYdWQTKIGAOFp2HUUNCqOUf0kgPdRdsN/8aG1MbtZPDeWs08gosmHxNWuLLG
4dNc5v26KP7eAMI5qaEp+HhCNeC7Z3z662WFjM1ST7mwTcYIw6NxEz94pssqyQTf5g6nyHt2D7Ry
VdBBSwvanhuzhbIMkaG46O4APR44RfRlcAXqEkJtABClIL5OmF+8F+5SiM2TpoesrQTnF2fn5hzE
9Mw8rG/VLvsUsMifxcX0bsTkdl0A67uUpKs2VhwkBoVazKTPWj0pnXcO3KHEunuyIvZ4u+XznAvm
3nG7mppwGTogsJh1sc7UChLNEsSG/hmTK7X+0K3dHzCi8OFN0IIBDXqpYfPlVH6fFthIt2hWO/gf
bmK7mqWBwtFR0yHhGQK1rYQAhM5a6wcYqNYbh+bgWufH+e/omw4/ll0zjdHShFtRWyRQ4GByn6T3
xX82FPKYlsmvTfQ7uXfGekQqLQBvZ9E+643sxNbT+DxB7kkwveXTHjBkZvXrIiOUtr6L56Z7Q9al
rhBWW7M4KFauRAKCxnImuf6B6pL3Af7961XJ7DgOy04AyyKJWEGLrP1FpplEHpZ7o3JQXuDzLuqi
DdGKznh0Geindi+mow5xYb0zTojYMqm1KErQ6A3nDH/lqu8i+T4w6pHrFw+bqsgPIve2RoHOeUVB
A1of/46XJ6GdHGpb6WJtnsgdTOrK/1nRll9PXmojbXwV3bsdpiL967fmlDn/6Ij6Jq23kQpcHpf2
1tdfTGEc8Rveh0MrIC87X2EwBTTply2vfJGYZ7w0Fq56+dA+vTzJttd7dPOZYLU0SeghY2wccip8
4TQBDrC0C9WiSHP/CbuwK3Zom3IShNU2Vm96P/RMoi7YJ2SCvDBFEEAeo9CN8+WVlWbsvVv52ed9
PN2m3m53iOrR1DtTxnPdCZJ693aljW2rWeQ7OTdA5BcMcp8YWLorUTo2THUdY3r2GWx/V2Hx3uNd
gSagGKoOtpFkUiPUhYu9n3qpcSv2Wf88Fce/1Q81rhSuwS5RLIkiPzErksALw9SYKeGCxNRTj+eT
RgFQ0QGhk2yZ0UaYughXjf8j7X+hEcO3e4f6eA0KTHlJkLtNRdikqMF9YaJtgA0di7FXjnR8qsmN
v7X025A3PS65BaQuY7cLaIXE28o2e6yqMwKCCwc0IVL5IhKdIGd/rpXxb2RTkAMJ2R59agqInZk6
qHZhvkWSTPC1AzXVivgsanjSCbnhzIRIk36qRqTk5Evgsi3D4cf2Jt2NExAx+oZeirnYc6a0bz7H
333BVufsWVxsgunaoMckwZNCb1W5BMXgvVCmCk+G+tq3X6mSFJLxYaPT5Cw86hsgFiydxR6ePoOx
964Xo9K5k0k2Gr9/656bgvitfNO7nVpMiUfP9VQEDjA3uybrySSbfCua3qmUBqSuXwBCmQ7uo+sd
iMIrp9xW35MrLPP1Xwaw3jKREQq3CENOj1krtF3dhav4hzQ9/vZ3XqrlhCA64a+wgT8MqbCDnYgO
03M83GXaRJ/DBxicFSVLTobPqdmj8O5qHtPzB3bzUW5sN8ElF1NJC+g6RVmlx/UBEgzL+BeWfWnq
OdPcD+MG+4OUzthbJ9pKmbd+282qYx9Bb471wKFRBcQjEpJ9OmcVe7HRU/Y2p31SxdI3pIdmsXlB
osB0zRuhLecsru62hQi2dO6b/bvdSZ7eB2aHlHizPCgQwAhdIkXYQWRpa5LUvwSRnlb71uIAJ5X/
+1GWhWiXMwZdZilgVukYgFyqQ/VOiW0jJ+UsOgcjH+QR2GOoWoEl+vyxI/Px1D1jbiXgIOtGm8lE
+V2GKJCGc0jhArDRaXO3iXQYj4WxQZwHdJQqSe/6BSWu+9K7qt6mS3ixZx4egFMEzePTvIm43i3b
AIWtscJ2JHCTRwGaGIwF/uemTuwYZJMkJClBI0Big+1jD0Veml5WDeIZTqK+3XudcFqfg1box+BT
NN4DSiTvaX1EPWXz/+ZgyapWvhNIqWlhvZ7ddi5JjtthqXcY4yTXKmXMKK2YmXc5ivbkleVVCGY9
cNLp4xPa2vpMDz/xjOg4GUKRQqftnVST5BTXUaSwXke3bar3qg535kYwiFx/9n7acAfmbP/6p5PL
WLelIMvYlFjJJ1vj88WIm7pXFT7E/WaMkTf3Fw4X4/yQrX7/d4+qvLr7jUacsyxLn4VyGXlLpiX6
EZEZOGnFVwnmczMoVf+vIlVo8MhezRohMKzWm1mdodo3RU2so++NwCP5lwOK56oQYOT6NBmb9m/j
piWZa4sWD63qerzRslkb484MiD0CkFmr+4G1lXGqhFveuwEVv8xHCAeteXnBQiMCpJ4nWVhPFo4V
UBUTb0iCTvws1VjMUVHSGwoJR/evCALx6Jlvmqr9BmKDbbl9fcqqKDsvpZcX1gyUgaeIf8cHkqXJ
1tbaEivo9q2IcKzBMRzy7uBh1H/N2pQmiXWBrRHkL91O2P9aQ+LzCtGDy1dZE2I+u2HSmy1Nq+an
Z8uS9d00Sxczr8XxvN8MfZQ+0yWT47jejKy4M0rbF2e5ju0P7GUw0Zduj5iaK3uLV0Ke0vY+OJ62
+TgVl4CMk/kuuAg+HZIzpFgPN+NTly5DFEajN3CYztKiSzrvmPhLSY25kCnJU1Jbq2GfZxiUivs3
/VFz9hclH7IsPkENRWnhuYauZApd/jNfcI0vJIZAaZ/ih3SJRK2+ddgqXMHjL8mKimkMQM7nhqPQ
0/XKJMBv7c3gGL49ntX2spT9lXdD2hmc8vINudgGJaHf7Qm0EkE6kyeTeuwWt+h/sSKeDCwHTq2U
DJ1sUAJbb9L3fsnkGud7S6dafLVVL3FQQEnF1JqXWzN3ykWLXp8TTtn1CehQJprAy91A3v0x9LPc
ZTb/ufZZaEVQeyTaM5OYKs+ExQERFj5RqrpV4rrHknvHqV+R5dy26Jr6xqIsYl/oNqiByl3xhDfV
nNtkEqXQNJxbir/7LGoE7sVDKrgjWXCd8BDMNOxbg5w9LrG8niZJNZQW9FeuXWtYWLagJE1K8bco
OsBqjlJDT1n8raeLYi+sfmAGHj0n+MxNtpluZ4ohTU9/VcwCfaCgFfY4H2XtcO52CRO+ySbRz6o1
K3Y7s5iO5pDbZbyoP5FoJjdyzr21M4a9/cx5xT/CPE2psj9BQRzEkFzLl54zkWKAmGMnqXsCSC8I
LWqSt3ERUHBGfxowfJwsYQiO2GPTZL+/XMpGHPC207La4JkKUmkTZyfIGDKJkgIXJ3ZDcgX00F3b
7SOgdDOW0kMqscK4ndNhgJGz/uAaETRYqLDtJUPap4jg7zb46/fWrz6E2lvG4DQgtuQGb8Gd+3BB
AsLPFf4+xfCs9mYQRVCG2GXDwUlkuLUcg7Ti/TcyAK568aK/Evu7mJ6c/ERmh1dx131Y8eqFQCpx
gzwV3z6jI+2vcJbJX/TWFmLEhfDqJupjPLzU+a8bkwoMKKgng5UIBADTUFTro668CtVGojQJ/esX
GWoxTEdFhuOC5R9FjWuPxkIlgMWPCN8WozgodBIQk88GfBoGrNJrxyJ3yYMMeYSDb01sXroXiTuT
GrEQ2fVshC9KsKWvyu2ApmDnDRvC4cMrK8HWb1yumNsrn/n1bl/ahcvyTEnOZ7ZGJ4NUc4+K6926
LKoCgBxYceMnkdTPWHsPeONVjEojysodNDQo2RjBix1oLLobJZbkuGLVSRNtjXGShKRHJxNxr135
Cp4fme2QXUQ46XKCBDNoXxyTmCAnf2QEqjmNpoMXNi2TQATPNueGhcOaUIQNwdT6cFg1GbleYVWP
7WS3cEQ2RqBlk9ZAYUD8uCfrDM8TnT5Oy40j03PxNPgCmO+/dCVgZ+JhWlzaC2TrlHrhvizOXrFJ
gFtdNbRb5UR+/+ZDoLvyulrXfizPlYxdGO8tD71PeHNnnSiGnXK88EgKURHBTW71bc1AdkPfMVX1
oMZsB4q5W19YGy1eqSPkWGOnEH+ECGuFyLmo5wvRwsZD4ZEa2UCXjJeDTIY+PvZ+D1E6B+ghPp0k
DEr7S+sznkaylL0xq+v2utnWfdL9t0MYE1F0CAIc8UGmcsssaZxRiLAd4P5Vb+HCAz1O6WLn58ie
Au4k6OCnpKspAgx3a9d30hbwiwUwXVOP+F3hiRlq3hpaZE2c/YmqqtH1Brr7qGZCEJvQv74nbw1r
XXCewWec72lqamYFekvrwPn+/TyxbVsKUtXxDwMPOxfKRmj+P+yyvnQNS0DtXXkGtIfQoLDzKgN5
ZrA2AiLfXLqgUkU+Ge6d2q0QxGjF7zQgt2Sk0QUBs5aU4oc71csQEVkqJ6y2Q1tpk1O0MO8v8BOp
bQ5Jj4hEjV48X9zA0sapWiornVh6p062pfKYRAZrj7pnfpMPYvqMXQKpdkFaqMHeZWJJYauhDuTZ
BqFFaInojmF62DQe/IFOT+Wv3DtFC497+BNJiK6RoUMzNJGmDEev/Wa1t9xJ705Y1YZ7RA2/gTM2
/M8GHtRQEQT+/BCG3wttkQ8k7GvmIzEi9w8wUdDYdMTH1OIp3yrD9OwutZ12yM5g34cETKU9UBnp
itCXOS4OV8di9eFtyIGuoJxRGtlAd3BVT6luPwAv4z/J4xPbGlFZxo+phHS3jBMwpUJpS/DLxHwV
trIBZa4bbZTF3FTmctocjagjowGZppYhfi/SmOtKF1PrAxMutt/dPvehGPbyJwjLs9UXSvaylPWU
jG14iAvL8WYPTEkAy7dweAZSo1gw1V6EIr3ELmMEXWXfLuOmYo2gIf+THgjPoj1+03626HjuYSr/
+pYwSl3CYgXqMqjRiFRqycVHkkL7KeiKZNb/nmobrj39hvkFRSBIw2WsaJHZYzgJi+3ZTiisLVUf
azAkMkGTX9E55BjwdtQ94TNxVQQzwZgdOxeY7NWeqQcxAvF5GeMXo1Zd3Hsi8TmNvUcaELhunhSC
6uCaSjtsHAmBuUnYXCz8uS3ro02gHN5DIS0qM7uoGVErkPV3M+O3oW1+LkMBcdyyiBjM0LOmF/w7
LUejx8AEzDoa1yuDkzzVETaKg1t1bfsnxQi+H7WojOjbcJ9c1SI3TFxW/GC8Fs8fVs9xDQTIdmf8
rzouI3RUjQyDO6uzwSTuH546hoKF6FaC51EAH2tqKR7T0xqLyn4oOyIak/GD8UuAtbJEy/eFHroB
vpgrYa+1YdRxXbw0AKCwaPDi1yKC5meyetF0EL+RZTj90Prc8ZGN5elVTg8Vw+mZFn0Jzz7BSJpO
U3No3T4gVs0pPpFRfy2CBGfIginEQ2t2JNDzZemd8aCD5XP4rKV8i7o8ojRUFmg1Fq4YAEoda1EJ
vqFR6WMmJWKURnhhHKWuMagDOIQK2At7/gP+G5ZgZE1H68z8k6YJ23oSGHE18VwdIJItOaTd9Vm0
MpLV0bo5fwBM07AlzwCq16GuHuGzx8irn6qvkudR+l4y+QiPyNcvm0/NyjiCw7hnsNHvNBS54C+7
IDDNHniSb/r3WSDu3QzHK+jDtFIarx1EQ4zM/dpMnaVsVT/jFweaAggfLhnS+4SdHUw59KQJhWvd
0Jk/WRAxERO5brrwtROyA1G8x3xAerqWT1/JFzK7PtVohcHICfqlQKVxk6bAzLIeyJOpx7XtyvJy
36vdOVvpNGHaewjUrdsKtd/A3KSxNTxNvbNWGrCb8O0EpXYa0xq9llqQwM5tbfrduFfVUkDQTMdv
G9nYH4n5/UXC54uoBJ6cOXpSZdUvsAyf6hwZG/MTzzJlLmFeHNHM25IKNFh5u1Ot0aLRZZZr2CyI
4q3LEzCVm6e68vLqOooW1A8C1swkEHzNWITRb9OQOZDRFCdnf/iJRa06GXCGT1D296Lcvi9RW6OX
MDgrgUAGfxdG0l9udvaZz9D/KK23tHUu0SpT+EpHIzB9Q342QvR8OAfMewqNhcxSiKnAiBHVRzuu
K2j2Rtm6IUMF29udLy5COwFAFKwq7PqHTiS4FHOokSvk/C2l16fMtPWZpc2eNIRRRGMsqib14Sqc
giZ/vJDzYWdcD6qXtAtLkBVOzWEvYemgzkGCvaPTPJczoRGK5Dv+MhcgO3b8EhPGCg3M7q3XDOKN
tI6Gh5w3FZaJlvyNyUVcC9QzMl4lcZRpDtKnsJ52qCwF3KMxH9k0s+TbZ1UvO/SKnAMLcuWNBFlC
MrZgUw/B2Wog6PLkOQy/ddB/OI7/SsA09eqO+RAbZ7O0ZN8vKKquhiNp19q+OgOTHiz2818OzHn/
OOKddLI3OPMCLbui5zPZ42+5NVGb297luU7hnhSiaoRsxO4yTkPJ4orqEYw/+0RVb26QtYrWaw6V
fKAT8LFjhhHPSo7PkWGsbzBIqXOJ/yBtA0hvb7oYtLzCKV0y4e0dG0negMC3CeDxsHXJ7XiO7S2s
r3kQtxn2vLvtIQ9hBcETLuJVzrcuh21RAB574T/3ehOoHbSrKfmTYFJ/H3Hyiguq9qukFqGqNWPO
4YQw2ROjXu0UoJSsKDNYS/pPpTMvh1Pqx+Llgh15OBrSvcG7z8DMiCIrcx9IIQPINxRyRYlwHPwC
nfId2I3jDNs26aFA3tgh4eWxmxk6C5f+CX4OFxOaksNKgNmhmLQUCkXQPuE6tSJHaoFTLFAiFyo1
lJWKF5Ivji2nvrCIdKVnks/3drg+Gw3GBbuM3D0sKqFzO3dvy3pQWirgzRFYrYXO/C6HbR1J5iJD
tD6uPFCk08oL8Ex5fp6ys2MEg1kBc8gswovTZmbjxkACVlPdEkTjh1TI+h8hlrF0+stJnaUxoh6t
yNBxeV42crdDX7laZ/G1ExzHmb2pWd2pBevmVbpcFRxmPLFdiqjVvGZn/qI9yI+U9IaFbV4h38vF
en29ns9bMdFgUs6P8u9IaY6zrEP9ND9KuhuTYATB7j2P7wIjE9aF/Td4FRwvnYYnyr7IA/wrYEac
Yh+3p2sFjqPzY4qpFtCaM3QVpUx9zf5bc71q2YqHT7vmuDEsRl0/OjWuLDTVH044OlEQCMNc+QjV
rbvj0uVmFFFlSISjOJoG+gqcLfE0j6gIt3oKWc2NFfX2m+ZsK8YWrluPBIJt3eR2JRNxdhhu4yvu
BlsjSQ77FpKe24Cy14elcE25hyFxYTNWKkmZq/xvB07RWwIYw1fdVAmTmjU5E3B1Bl/9Tx7rqwKd
dlB9hJjYvWZHRWGMOmWto7N89DyDGvUeTtty290wA4pUnQ8tKQKL6HsPrSN3QqUys9W4+mDRl9hk
YvrR8GKqLbb/ynHN0r0mKlTz28x0K1pOS6FIfhk/oIFMVKav2wurj4Fg2UbNcU6+Sz5WAca7EDFH
WG6xqCOoRet6mxSwNGUZNLlVtYB/qkXg3JTdc3TGEArdcMOIZsBkOys4/E1VmrhOfq4Itmnxk/uT
NIuQf8P8f0zPbH61wnR1o84ahMYmcx3DLL/dO2lFQVfey7HTWkDyuD9DV8cOHPDQZBefaQzT3fgh
LzDiOYLh4LoFtHDiLZJVQNCoIRS2mME1zPaw+zcPvz00ykaLg9xStjgaTVG+dXLdLL8TpVE3Yy/D
bePtNMqDeaSPsyrpn/IwPBWZd7ll8jchTmwl9qlfRMts25BmlwFINHYZ11pn4971lI9dpWIqV5fn
2l3vWkXaHjpPZbw6ZTtGIA4ke4FdAirD4c13ksPXEI73f8841adS3ygbziXb199xP2LKcJL5Q0Jg
BGw2FiFBCoVQdD+dYjURT3kCMuHnxoO7zuZfuoo/G7T+R8qfDbJFQ4KOgEno2MBsO+Jm1wirzFit
jUYBs9PIthuG+3wx+1HmTs9WSqMK5OPCJeY+0chOMT4SK2LGH3AqXjmbv2Aq4wgOTU18w+WRHHmb
s15iDCj8nggcZpWjDAZhYc+piZEXdKN6Q9iar0FcBFetK8BchgIgfidISmqxzQPEtZXK9Jru8V+n
ZSM4mnh2lvNkQEoKoHBS8nBU+TfDiT9YzQPl3Mv1dvy2DhwdF7ce5rI+d3XstpIQKuZTGEBXTan6
Kloa9N5oqREfB64Xz0s3tTWdi10gB/60Av0JiK0Av3UccZz/+j0QsaM9im63V7e52lW9yhbPEAla
gi8I1zY8JRufV7lj93Mn7ZlUnIHHvAqK96Ex5N7aDlukrA1p11pHH/T91CD+HS/SjnJPx4QfXc/l
HZ57zn7u4iGBoaZiuHlDVSbiyUVJ/y0xYToPIHwMRDSZ7p8nV8+zLrp+RsSHsSfguYE1sfVv5ks9
XTQ/1Pv3m+gcdePc0TDbFKHPXI6hfUc7DS0PAhrxP0Q6WlNlXoPPKCHbhOJ9gQ3HLdhmLqKXw1gu
Yg94Cw1mCTeE/FPPE1oOLUPuXIt7PyS4V1URRH3mz0SZINgPyhuoUIi++01YL50lH5UbqqBL/U0z
Z/W5TsonfizVILujDsdb091AKMfz/MPpqaaT1jayXhY4Oi9TwFw+jSNhURvWFTeSYez2DcLh/Mct
N6aFm8lnMKvy8M4Almc6/0amJImUM+l5epoLzMBaYwzUTvXYdF0wsXw1KDBah+Iw8nMjg7kKathE
OMKzEWn5VHUpwHaokJH62cwDL50o5431OUmUqpCTnj2C8EdfkU6dD1nJsKuqHG43Po2Pcwjdnsv+
1P/nWeKRIufyYakhJxZmR1rz8iGxM8AJxdP5ARKYV2KDYbJK5+vMQkX/eRlvZcIq3aPHBJ8tho2Q
E+9vLITvAIcePD6nbjLU3bOF6dicBX3ZribP8+EyPJ3lJDRjYZ+dtvg7hsMk+fPSiHxqZHz0rL3E
Pbpx/TstTvTGhwaQes2xO2cg27nfBLM63oM4WYVR3kEG1T+8XMP4Y9mdb+Y+CbIg5+2RYmUMtBkc
4VEOMqDO4ZY482+Ven5U+j/cLosBykpq0Wxaj4QMRyecdLoo6L9uEeBM0qOPfV0qTBgDQLoQM/UA
Sz1usbZnNYfpL9es/w0xJjf0Oz6XD6RrA4t+gOzPNxxN6vEoG7+PEbwLbjFfnJxvUhg2affw6LFT
LYFr872854EW2dLku1O/ZnqEHsqYVjfy5kh9oN/vkImoMklt0fMtoaJkEibTlBqX5PcnBjac2CnY
CrFsV71TC67ZQeSl8xI3/nH5ui1jZezMPJ7z8jJo1D1Hc/7LAQiIqc16J/04TD7zpxgFYULU3RoB
FF+0aetK+Z2AxVNB8582cgwlpGaPOT9RvLAW9QqgJ7s9/KD71SwpyIkt4Rh3aW+o7JZQIC3rgeWx
B96JVomooHxpw91N6HGinYyAYy701SsCKbm+WFe4pOHHRYtdrC9F3PF+t3eNYqp5EObWWGGTacAF
emcqChe/yZYNE2kUEfEzGhTOxsB4hwiI/Y5/nCgKZlp5cdt0T6U8AFPZFHQtGJpVmm+xyvCi8Sj8
+aGBSzTkTLkblFVQZrjQq5Xcf7RfYtl98t/Zg/W77CBL1RGE4oj7oQj+BfhfADPTbAtOakQnfT7V
b4ugw/nRk3Txq34dcE0HCM6Eqqb2hOvpErhDE26IoC8G4IqfaPzbboDFJc1JHxgY+JO6Ap+MqWI4
MsLeMUr94CkpREFejN1AH215wOLBdGoadXkwC5WJhacYLf8OHtasG7LYOKvUpvd4Xoa6bZN/8InG
EQ/IdSr3DvUpP0pQADJfbRORKtWBHeVd3RrRAvbPpmRg6z2lBD0Sd3gB65B1I5h6FoUf36AldTci
xLLb3QDQLPG0+wE4u29puS/+n+NNEvRygJKQbi9mwdlswFrazxvlptlT8VQAam99Om4XZR6ykukz
gEuT6XSFVUtiHCaLXl5TeeZUKQTT6lHEIRHA0zZzTu6BfFoIlicmKchXT+1igznV9AHfFDkNKHqr
/Rq4fzym2RPW1wm1C0cif3BoDtVM4pNHgh2UBnJgaflmsGEmLLhR1wgWByEt4cw0qxXss4aU+1lM
SkppbKYzG9tc2HQyOhLbR9K3uG64KhCMN4DrdlTN9VcxDBDgChW9oIQ8OcXpWVlIrk6QIt/bbPrN
CaTHEcspdOoB8FXyyNEkn00Ioxpp/uJAoG9M3sKkNUqpjWAgPQJH40EIQO+GXHQeyVHN7G+egEYo
Trkan/pCapv1Tcr3HmWjnrKPEJulIF+8BXmCKMlCZcs13wVJWKMhUNSXEvkrwB/NcpKFk3HjwOtG
6ltd5lvoJSEALH80Wxsujg3xACtrc0J8B/jDms3DfkbWeUlejjuRvW2ZnTAtaOgh9ygPilMuL0Ti
h9SM65j6VwUG4yI7HmaqyN9XkUm4FXIDOA13DAGSDM3jmBMCgbpjlCTy5I3XAzbY/y/3hJhtka5G
o4oatXCp4l8AwFdZjcNExHE917H6cA/L4xBNeLAZXmWUchWKH93PUWjm1/buVML/TuwBMy1qMF9K
OqYSB1q7BW5sS0FSl3gFxMJ+6QMipgPEBv6FMTwlub6PHuuAVDZTcGEnTC6mmtaUDnB99QDGgCEj
trw/1qZjTNrL7BB/etMm3eMu8Wxz55UJY7W4w+ytY7kAgbs0Cp80veN61S60YqT63uMK1EHqN6UE
AOuDxvVcaqqk/E/9ICTuohv0BUbUWdgsPTQ1kNOUT+RAQWWJSTsZ3L6fzTP8enS8Srbgvg0IkBQk
JNYj0WSOWcOs9z+ChzwQKlzDnE9Td+cnzLEmU8VmdcNSDBPr0tUldURGxfzYURZn3KhrvjZEoXny
z4VjY2SRpTe4M/EhMoXgjyzAVh6bv8YbiHl68AS6LlDP57q6DM3MEF5Gvfse3fMZVK+u0VJC+Gbw
f9LvQl3RfHikdQPOjZM/xllVTpJvSXuOtXShiEh7jJRccGB1FBs3tBNJ0zf098/zFKyzB0o5f4ME
uPgAanG9jUXBn2MkELvsQ46yFHmGfvJjx/FVXrzQscOKantHAw8FZsFtL452rLDJ3YBMgWBiGx3h
x4mGb9gsDIjlNSjkIv+JWTQiAjXySWdVGiDtVE699zF4Xz5vSFqNxkuL4InUv6ywf1bu04bZLt7l
BeYktUWjbbSLKSIMCpq/wrg3ixIgT2lrLAjMDXrDqxHnb2qSwR4JF0VSJq9nDDRJQGAY6uRlDtO3
VuNWJlRQ7PoVAwRP2vsd2ABBMkDlNIRYJKeHZ9AyNeMYiGK+iKbxrYQzkDvpRHa3JTpn9M5UZXz3
+ZEM0huFEgRckjM3I4rEjzdKXWT5WMr0raBB1GRglzPPpl+ioETaFIRadY11sACEi962059dzOlw
0YeMPdyO9ZE0rFYt4eqoUosk8bLS00p2+xvQugQilApTmfafVo4njE23yPT1JReq9Xu40jJeRyIz
afsr/I0KZTb+ibCtiwPFc0rjutlEn+8Y7UkpRTXLo7bLjLVIkLEkqkz704V57ifcs4WvtIcSOxOh
4Xcbzg7GYdirh9ojpIUxV08ZcSSlwViJf8wAftR9bX3+1Cec/6BiZ1yvhjDhXNxYE5Y9I4TG5LrQ
0NKPwLMUa+ldW4J+DOkKBEsiYrOc9HwP3RHbd+T/OpyWgQY6OfoSFzFmQjXSBb5SCAXxKrqFtswQ
6UmVgedpC5txZfQvFnOTXADOaUvgu+Qu7MCc5RQ04/1wKpVIo6cjvJbkB1l0a1ymPfdki2VO12h+
lUSttKwG3WcvxbOLbK20FpmmOteZ+Y4so7pYsbJ/O5jQG+ZAfOYH0Sx3Y51uHmuCd/TBP1fmegRP
wfTNN82u6L8EJ5GQ1t/qYcJoaNg7guFGkcc0FQO7eX9L6oCJXNxPDWmEBjJH31RAOpRQiLHPzNLI
iQtQsDBqYI0uzMH7moQehkcMn8/0E4eCiCYuneQvK011BzcPsE6WrACuH4BaPyAq+W2VCabme8Ot
EONsh0i6agiMTLP0fWlyO5uEAdvfoKliO4PNKyFRzDjfNN3koZFo8hQ3cX8fDgv6f/GjRg51AJ9a
UO0fFmGzp+9fv65tWAY0mlAdiCxRiAj8fIbSGvsWeg8EJGMAIZXiKX/j/YdpEktPGyWkBzFu0hwb
5rHyX7caCtKyxJ4MvMP4csYvUiKzo7w1b6wrvfTf++p8b6mFinc4cN7TQJ6xGhgCS3WcfrgXt+Tn
i/PGDwHIsr24XBHptWJN8Cr61R+w0rmiBRx1yrvLFTIVmFxLmj4eTJu9WWIf8MA3eCM37vpuK7hH
viBlnKH+m9L9v7e599HLqBQ+i5C5UGXZKVtNH3RmgGJKhGB7DElpA89GJFkhIRn7Dz5l7N7wLD5C
0oB5iybF+ZBM8IE4kNntAW97hfxbZeLRjAnsEJHp++1goO+LUiqyJpsozFpTRkpFqNFLfUyMxZUw
dw4Ku5xvmlEJLo01UhlKs4OTfsHh/9IPMSzEawmcizMuDhCLaoa8grMPnm58pfPWMwpwmiCycf/a
4BXkpgiie2meWhHB86WWId9WTPotkuQGpZ2Nh3nt/Roxv+vL98c15LZEVPdSF2YCg0PLXbB6DWXk
nHqN8V2lajqC4NivTJSe3ASOF3leCpG9WVtFp8ybm5wUh16juJDKuP4H1II5Lrd1YU26+NNk0JKY
7XgBX3ohxIMkWWXQJWPWUeR09bKeywhAzI+f6q/xAWMPAdAT64ide5+JYO5mWQNKWnDhElDjzP4O
CVOoBY42KVir6Q4u7TQnQFyJCNPjqWnPWApWhOc/eBen7NXIFUQDA5QVSvnY7KeJjHFocKBKThin
L20EoypPwZt3G4vTMNG8DgHDSn2c+kYeMfUnX0bPWUkHWfXazZ2THjY2xWy7uX5lX5wvVcN5bWrj
Jzl2qfw7XFZgtludB/SEdLJWf2oTzdPoLCf4Opgeij+zBW3vc3p8dl27gBgoz6gZ2CngZ6GgpPI3
hk8QUcKR1VKRUkxqNeF+pONL54DdsLo9ZGyMY6tvU8+G0hibYnqvPrWoL6RgwIPV4xtGlj2ZDXrP
BaZNgo6SAIuC9fPIhOUP/+o4fJ9TpsVQmhSFLoPwAA07dIlqIl7OxB0hhGPA5VoSJHfl2qG5QqTQ
Wm/qELVGAs7dYCnerNshyJG8RReS2v7jZh5FkT9tS1w5LrzgT1kKGSJYM1GOFh+jFewEwZme6Bma
1YZxKGjZUMh/Q02gtkZk2lK+NBFvG3Divtb/ujYbxIdtCSj8vlPlz/Ku5pQ2d7cWuWvBd2ht2nKx
1BZj8R1u2rf/1O3PFdEjasrRZvNVxSIo5vEzF1f3BU3bLTVahAaQ9L7x8IUpPnD+IO78EtDcBPmj
+HP1duVPjLP/MspNFuTiwNTiq4pEhPBskXLP8w6ofRCVyImFwnRHLtcaLVtnp+E/OxCckd6D9WY2
FcHiCvH2Uz6Sn5q4/xCAg0Z8QwDuRr6DYV7gJh/F5DK0lBLXv1E9nrDHlmFtcs8aWxZZlWkXaTN+
M960l9C9AZK4QDZL+SYGVKzz12HzY1lgiHAeGpIi6b5B1qczPg+Y5mzudRighuT/kMIEt7tpvgrG
sQhtuDGY1Iklj11xc+OkyqnCcBYjH2Lx2z0zenJMQIy/jlqtqhODi+gksU+kdaXwBQ1uTlRJRTJu
LAYqYbAc3F1E+UqG52Z9UMIKeB/+Twop2JihqUPYesrUq5SWtYTK2ZylJ+wsRYgF+5rmx5Q4pS4c
FAl6ZljT+YVTx8yEVbBcAGv2HXg+RDYQ0HjuzgFYJjKRkEjiUJANwbtIi2j14VqBXzGeD0A1+s8d
vJpzPcZD9j1dunT07sAYiQCCwR9nyutYPmRnYwXnZYzPvEkA0XxyWzWW2cl/DEx9xuyL4D488lNM
6dMxEWCRneSBLDS8N6PZBkVQeNHrDyrujsvbdbhxZsQ1yP50BG0tE5HcJXdA7mSZLrA0p1YSzB1X
jOzwpf6WRx3r1+eJro0YJS7VIbGmssh0RBOVHrCbtg9YTREYJoveEYBCqNzMeS2KXflnF7tZEKdG
GDVmPORfZ0wXaAOoAc9lq++7NTlPVu2/2wAXF/pTqXYBXElF5/EMSAiRrMzDJoZpM3U0Jn3F7AcO
iVhbJ3I4e0kMWfbVc+kCY9DSa8er9mQXf3abDCc7OHrWyh1utCu0fLH8A9p4W3i+4Rbv2QF4NbOm
O1/dtVL1q2x+DILpC6H1vOvms2vEU5DTi0lVhuyhxtKQORAfWoz4r8HXn5u4AyNAcuXyNulomi4a
oN6Y9YGPjtLAOm2yQ5WLnvIaEscUcqa+S2uoMTULvWuzMd/RScj+4/aPQyQBI/4xYFezMppNFs0z
AvX9rQf0OHmE4AjOyBH01VJl6vjk7ZXj0aGJmWfiQWWmXZvtUpgP+btZloy4lTbrsoJ9r1QtaXRN
OLZJzocrdvlAfFSEOrdNan+aRdS6yTTyjx3epwBOJ4MpW7kVdGDqbWGOMtMPiVmg9SNTnlqJfdGX
Qan1AlYTvb6G7Bidi/a9pfNM6coHRVsxNVE/Sphfyy/fK/qv0R8bmgVCPETkhD1mhVkfXOdmovAq
iZtiuYBYuc7vUGfHGpvVbW5/y8UYiay8zoqWBZXKx+YNI6/btlir43gN7I8Dw6ZvvH6XJuoR14nt
c1AMOZcvJYgM1hIYVwiR6tmba95VofjP6lhj2HPWd498IBLExjRZDVLq8kFcGd7bQEhVLUDByAZm
utAEgxW7yVatR/X85oIQ3CtJfGHFXI4FzwzQnSq48MIBkB9jlQ7X3lyDs91uM4ptM1uVvyWUXJjv
yGrDbAECwZwI1x7q3rNoDAEhSOsb7zdDbbuhd1xz1n2th/oirV/L7OpRLmGbgZ4og1/mfRIteGjX
q77wrTeDvNhq8Gv30fo94wKq/CkYaOHZdE5MlfPiXLvktjdlDkplUTomQbolDQZ+olUP7SVfLEDo
XUpG5aTnW2VoEjecz0empwCfa3q1x9MuGfEZ/U0Zo/I8E+kNnfCL3HwbEmclziGPlKh1jOWop1J2
8g/Uj1u7x/t4ptwG+Tcz3YH6JQ0RaqWLvYe6UC0FTC84Tq0xru/b/L/g0XckVYW/iHCCO37hQw+Q
OZlAhe9vB5ckvoSIUI7ubL/eaOjscs5oHC7DlIS67JT5zQxnAP61tM6LGY9G6bwNvHKztR4vgLIN
D5mQh4Azn7B4LfhWfKRR4bwy2qts9UbseiGr4A1hsMMmV5Em5nQhMYZxJxwH6TfDKwKwJWqnUxam
2NVOuiS8l18wXoPtwSBZT8fDPeQJP+Op694aePwhMBbMEIlEAibHWL64EmDpN3/69nsyzDPRJwBv
kVUAspj56WPX/w7MRX9h6K2h2WlSuxcAbuOe3cP81Unn5S04/mvGi6Vpx1qCEu29iVIa7cl64sSz
04ek+85KMC1+/2WjDzxLZc1z6zejsur1NWrsgwhQpybLcMH+vKQ4nb3zy2u5loNi+Ggcxtc0kJhY
pt8CqGP0XJlPUBJmVuqxudLiJ4tjxewqB4uBRijG0IbOhb0x9x6hryPNcJbgia/FjoFAqlXy552g
HJ4fChaS2enSE61agUj0tN+qnDT3BPohenEDRJeKw/9sgh0IZnYHM2MOQmzit40SsbtcK3gutmc+
qe4Jovn0yjWEHet5luaBjjSR26M941igkU3kq7xkkd7tcEoPywtFYjUb153RBQ1vSElaaVxqhzR/
KRu1HPOgeswGTOejZfnCAFqi3MB+uy4Hd3iExiiW2cmk1dWy7wOjZeacI7R2h6dHpLWAFh+QP/VC
UzqiNC0CSZiKYpgc6GVxX71G64mXxGCRFs7RUftnbet1uH/0oE/wOBdg+HrlOQJNS6F750HG5wfr
txjvYeqhxfFpQw0bGzcYDn6XV+9UK/BsBKCnGXhXdujOJJHX8MfaEXUd4wy2dR3eQg2OzgcyFxqZ
ojNEZ9qhsU+2wa+yDVMVTUBHk29DAhLYy9E3z4CqV1swZqplTWG17KrzwlJxkMUWnqU70HuxAeE3
3Dx4SP19ykx1AdToiQEN4l7dPAJfwG5hduUmqqHXM/hSBL6tPm6UeuAuO3E36F4vB+/Ovwe7XZ84
nZCVQLj9BjdWJ4Cez5gbw6icXOyT4tJk8u/xB9NCMb9HtehAwsWfqqj9k3aaqZbGz8quVmPK5a2a
RWRlP9Kf3e4HIgpMaGjdR7meEOSub9KEbZphX1hF/runkJ7hB8ZXcVuAyNc3wWBwXVwKOkDsiXwR
mwpqANocZ62PfjHOiiEuN30OS+IIGiOAdcVN9pwJo6vDFcAkj7IOpakwRSPLMp36w5FoJi5a987g
z8lZyPDPA4WkmxUf9D9KxMrIjP5GdAzaq/SPuIUTUdk480v38OKDKiuHCssq1ndL6qf6a+CwCzno
GYnthk4/Z6W1ezhZQfYA49QX2YkS0V60L+5UdCen5/4UVNIqyG6lerEhC5t/RIG0fh5LvCQ859JV
2oom4U98LOnn3K9iQfely1EELFxo4gW8ADQHMUpq6yxkF49ic7auRa2RvVERY66c1kVdND3kI3IM
w1LKgxz0gH4lqnW4zq7tsNRpP9T4z36MKYgiOgyPUkuEzcn4jQKu69fRNvtxc3xBFy+gnrakh6xN
iZ5+YYs/I8RTpvs5jWgYUdCjYfV0q5jmj581LFq2aO9mRkJjL7xjlITdk7TurVbhjG/dmcwSFmbT
aldivEmd+hofWVgzrXH03Q9XsKQQuNt/VNzTM8hZaAuA5LQdWiolG4+1QcGMt2USqXN1N5pIwXyk
JBgFaMtp3qek74+pzrMEZfhxOC3HzMep6RTbUXO9i3VCMtEMelox0hem8STNSIIiupoU5glM1inc
U9KL8QMc06nCjgM0GvFH07Zc8W718XA1IRZ/XE9THgY5//is959njnPMQNC0gtTxvAX2rjx2YMZi
rCiR/in8JMK8KDGqwp1/vjqDbBCZRWuOCVzD60ZaQgt7RkHn8jum7H7klPS8eqr/kv7xcflWHMBC
xjSXgovgMeqwO8ssvA3VddpfTnd6MKUy3QLFVdxuPlvTEm18LHUOS+atImeQJMU+axEyDHrhaRsB
ZfO8U0x9Sv0EAxB53A/z7lKA1Ee9HnYXLiLaeAtw4bztOapUvnZJtJsk6JnKdEPIlGynKM66v3JH
pko8SXNFkewYFHjWgSVcfGF9+I0CiEl3G3lQ3F6tEihqegDyBzyBzWsoZG1xr5JQ4MAoO+C6UcOJ
hKuP56fQ2VN9dnvvEAclVSEr5YTwOGdhbJwR1MC0y+Q8dxgPqaA40jPw4lwa9a5BtFFecyi2oDDX
00E8wH7kzWCAoC+tx9roLIhFMMK3kvUIoIfipj3QpEzAwAl50CNDKjWnz0aAgvySSFQaGtmBncOM
vOakVl6trm1gt61RWhfiwE6ZUyr0XaH6Bi6LwE+VsJNvyQJVNVxCsilQgS7Rho0piCsQbYZblWc1
+kwGX+penxAP07t/r/E50iZHkB13+cWP0XJ99KlW8zqkODIQmjS3TzIgir1CPlTQwd4o99b4G9tR
bKCeUzhK1Tn/EOnSjTOTt7vKlYQh7VW/qQZ45LcZIlzUBSAE6vNkVuAw71akH4IpkMPjx0XBaAUQ
j/IWpWumFMqZzebjxrkDm24lHtjRBsHOoRzdcH3b6x/qRytXqtCrQt74Jsf08n3OCU6NgN7QdqTy
It1VQDIHAu5SLSYb8EDJD45Y4zC3tfZV+I/HhgcF/VbpdYgNXiUz58xvqr+hKtpjt0RTDayx5LNS
cp3bLtA/a0btGmMZ9h1QUArooZPz6AOiYLrNrAusRzNMbl/5BB2A/2wO1NCbWUQGu65CB7h+wqmw
iImggyc5PvLbkrSSG7ITRn6L3a4YugHZmqcuoXFUsuWddNMrgOgAYGm2zryjgThRhwKmLdfpfMxY
tXlAA3BQbaqnw/qSyIj0Fi/pD3pECYfYL/PTT1zDA1NKMDc9QCZPaPsRIlps1Je0hqmhFlAEoCRF
XBBmObro1On0LBRq9/ycGGMDUXQBo6PAA8qNpJNhAYYePST72sk5/DDmUsOAlm6/HGQ1En/kizqs
ch1gsqd9PNdLdf+cB23naYCLRyAwC3vGGFIzM2lgbdP5bN95shXrq68mlRjLXpXbDliCjFH+RfOV
npW7XHU88I173IqNqEcUEpeb76XqjeZj/gqILrenbkPaUCdApuWjbbZk6muuHCxCbuoiPg4GgBtz
Hn34wf/au2VWmNF4HkYLZCfieLbj+osilEBz1/WBksCRUsMx0FZnUY6VtkOyTMfvQmolO+uRQ2U+
QR39PJGUG9xO90/9XdWMPBpWHmnal9MU0o3xMsu8xHiNEbb77nb7ueMpnERRDhINeCpVwejDmR1t
4JsdQIKA/hkJSDaz4hMNxFwBCRhYVNOWiqVptFiwl/y2mX/GFSPDN4IMBIaBeE1UO6Ah0ItSwpix
Jb2G5Avv6MGGAbcYqYZuQn0ZpOevIVo4WcuJ/KHTv6gUJhlCLvYO3a+ed3UzVee4VZq/1l0q7HRK
mA9wIIbTM45biNmgpPGKV48xdPV4UMPYmg9byLLXz2zW0X3hyZ6f9vO0YHHy8hHOaCQLg5Iudr8w
CW9T5JYISqGws4WE41i5e3X9J8lc3hEH92pZj89e19PXNlHPNTaSUYKaPZNJ4M7pS3tUDVk/zF0J
RZSVrjVlPyjzU0EvdPg1fhaLYasNfdMLDZamX9k3Nrojg4pCMW+FYaT3VyothK6ZKsMDzKDjMx5g
VIZc2cc1vW4BOILPga3fKJtdk5+MezubPI6HNVGHOom5sA1FMS4tmqjx3Yeq2+euGgPbRXTWBCBE
IjBDxZn4O0OfcFyF/qi8AmKmecBV4mAuLsdmm1/aJwRTTyJwoqwxjiHEbHGMlyo8PA7zVzxy01Qz
vhWiWt6NRkaUP5DgfKsvNcf3qFb9uS4+O+ykPIsVF1+azYNqfYlmhQEZdEVONlBgzje89nA48CVf
LtRQd1Qxa1dkpWk5Njk641kDewaatWZRG6Enc60QpbjM7+R8pfllL1Yl/XdLcDa96fNI3u1dO2E8
3vJvNylsD+7it7v1hYRTfKRHOGr4QPe/SMzabIS8G9xd4tX/SUseoVfy/05lMq8stnhLugxJpqqf
Kn/miS7riiP3weerRzoJvYzEZzicSVck5uj/g5Mu8FCwrNt5+GhupzvXVjIgs31WbfN9YY86I0N5
JdndF6JUH/28rXE/WB1omgOhM2E5wdvhmErI+pHr1yNU0jcyYXkqhZ5n+dSivFlJMDz5B9x5my+y
f5lY2N6/TSNMwwESyE4sS2jrsu20wnHu+vQVze8RlVs5kM5eXMP2Sn054GDBfV1l6e2ty7HIN4o5
xKZ6BcaeY04BdlFSZtfhb8mGGO5ER2Q2fw5MTOtXq6NqgbFhCBroO6VYpnjW+pVepmHf0gwIJwHb
7ILr6T9tqtN/wddI0h/aX5zfP1rA+OhWfgZ+xw35dHAB1oEBPHmtjprT5Mo5+O/YCdoO9rPrxMyA
iuK7lVYLRHPZjXeVT8mDKJqzpABVH8C//oT9nyUUdaHblTRfqeV/61VZQT536E0CrUs8C8FbqVjW
WsihhiPexVb0aEFh41FoUXNCY/4WmJ0tubwCp08+n6Hd5YTajqRjBsQ/6JjwGkwfgAVoPZMMAt1J
srBO0jwgvL0a4zgcqL5T51pGShR02+3gBIG41wK78q8RPa2cN3KIpaW4ikYTO9RIpDOIguIQ2JM1
+ZC9DeeGErbNWxzfPhFW/GJyHyHDxmBjuEK03UgMZZUZS94n5Nl9UxgtVLCC/tjxOcWafQ4QNCs2
J+bAF6KAMRu93l9W5AtTYFVZYGVL+In5KqtwGWJMZl+JbvJ5yO0XwiZPxPwMZ1h06Qia1/wgguWg
YTomGycMkQEKLydrq99DJq0HDvHTRSR93FDS8/UBpXoEpLC45mi6sCxGp84H8a61uJ0a9FcBsqWH
wpoMl26ApqLyxYLfO04QWLagIVI9o1AM0Kid3sWibe3veUH+g6O2yVCztl6kpzVSMhK/yAQ19a3M
NUFIWKYm+GmcbpUWXMSzBMosAIcJxSXi4ib004V7b5c4Dp/20cc+cGewU/U+Kw9GU0BoVwaKjr1R
a5iUYs0s1IwoYGqKgZbUW4++zrL99rShXE8txj5p8R1zUQUlzA3SJqVcUhOniQv6Bs3RzZiPtMKh
lDuQ2xt7MxoskidkHsYKDMw/r79eqCSBO+z02T4pECtGjp9o/4tMxtULXjx53hMIxN+UCpb2aD7S
zHXuEM/mqOucxYpyezY45/HbAljsCzneOiKM0KObMw75ibkKbda/tD3I4QYj0OZLdyyYfS7d3K6r
L1Viz8rqvbHE/98jc0k1JReRV1iO2+9/ARLHj7jX8e76rCjT9TLjn5cxSKwy6j45fXBadRvDkUrq
X+LF5KB9aq5HOaI1xD9CI8zrgqFOkfk/zpS26/ehlCloyATetrnKOnaykgxnMQRY5qCgOncww9IR
f8eNZhN0VFpwgabnu68WuQvKvqGiTqBVVcKKBh1OtIl/qB0mzzhtCNuKGevAjzPaB4j+oPr1sUBJ
SGC/nuVufAn/0FK63lOOILvy1hlxWJee0TnOOndd3VLCmPQXoV5zIXVI8FtYch9srSGc+8hv0pRt
TzoGGC8dc7ZDgQtC8oFHCNY4dHw9yHLKjswExgdcCY7ZJOGeaNVZeTQvR4uYNbf+cS59X7amoNhk
Wz3U2qnTeAzS/ycLwB1QTKMVb1IgfjbIH+tvuociB1u/cIOqWLEL76k3ibAs5QGEtUiKUCuzp/NB
OfmqCKsFO2XamVV+TJqTakUCCcMHKIUFbUaW/AV+VoLzHQ3o3d5twc2QHOgqE0pxoUkXUZl1s61y
B+ZUPvcR6GYA60EBRkndw80nsz7mlv1oU2Y0ix7GCFgeHtXUlObjjdy2zUtaDGFUqOfojhZ4WTca
WSfmBEQRLSw5gRt+UT9Ss4N767+pIKaWF2g+R8A1h9bWcOI0pu00wBpAmPlib5/0MmOjr3rqYihQ
CzkF7sBZ9wvgxfFwqzehSvIAxwRGdeO6zTLwiMpEieXPWWwYioz5HBYnhgRyQx/8R+Sc1PS0P9s5
hKkNJhYCx2MLm8xhpyheqFOhWOJ4TQqWkq2feITW6QmJJfbXZc0hfXtVs/ZI3ymmXUCFhw5npzFx
uzZ69dCm9OmnKFXudoc24wSQ8ywtOdEqkVYrRA4Poisiw86I5quo+98baQnCzEP4m6lEkeEkxAWC
5bUgpOU0TyEEUDWqjtCGn30BL9MavnmWlexxm5CfonMQkLjZQlJQl0MD6eHpy5VrDb/TiCpqklwJ
WrozCGcercDlv0fqumn427xON0tujLxZeniXrUam3IL+48pgyesfcddqk19NZREAQP3D250xLl5V
+jBIW278Lbml3XpjbmoSXFnrC3CjYzHT7SUhk4ubFtl1ahvEQ6S9K7UHCIbqjQQMXyLvlEcX5tq8
iRoKgcX5yWTa0qiBfAmY4wDf5GryHqB0R9UrYNhsnXHt2nYZ6EPhGaOU7xgSwtJwOL0MfvG3eFDQ
Q46KptC7J8NG5kssJXTH0tt5jsiSs/7a8u/MhSOC9xnHvJ6kV8vaSQx7Wo2m8Qn8yuXxKHUiyinO
Ya4XBks7TPUE+uZrfPvizbTgbUIBoT5nJRiI5V/sl6ybu20dJOf0XGHAv4N+tatiSjWonLzJAFDd
BuGMlLtfxODWImHShUDFqFraVi9L69RYNlk+B0Zp2ZF5j7yjdhz9tfID1Itzn1JMZav/z8Z53Zui
bjnM5QguK2TiKAuAzp87zmpqwK1qLAQqa4ewo34JwAf5PEEwu/8ioIFTsH5WAP56T0SJE6sGRhvF
4ROiAcZqXUcyPix65yQZuTijzRf0NP6S3dKm/8ufLqkiA/AaujG/Tetvmvjz92sOmTIyNj+LfO+b
E3UO1ZT32kXT/UAKB4R8P1qa8SO2onjL0XlGpa0bKCrB8G3dgd1oHztx1SpadRgED1qOz3/Ese/q
138gPcVu1GAPzxsqU0VCMx+km4w5Z69ACPbdzvKsUYgDXQx4vHIdTfRT4WYBH5owPxxAGzpuZzak
O93eHPaAkgiyD/Y039sP5aD7tEgXR7NkA4/BrJR6XBB3ZN0Lr/yFB/u93chM9IXf/hhxn7FffNIf
TamCSJGeCh6wIUWdBCQvhvWVQXt3tRHM7zbJ88iCJhtB5+Pq9dSNl7wrREDZ9JmJLN0HOxWaO0v4
Jw5EwTGmdXSaVZKtngDkVfYafDKDyx618nhmFw8gvGF39p1vcS5DClk2xVidwQSdrOBDwdA0HMwW
dtsRdH5Gr3O3m/2pHeEn2AEwQPK8SvNoQDpFvEoJsqbyiAbEkFLHD5YTa8qE48WobG02crSYFjvY
j8okrX/mlzI1Lo/sRyFSTyFUqGvHplPtHPWFav0+E2oB8+crp2JPo/SRh9smxDiaS4J72zNbmvf5
DVffvq9ReRd1w5YWw6Ze4ZLedmHJ9lc9oUmCV+FElz6amiCVHgtNggsqRUgzYqN/m545JBw+On4T
ZJWu3XJkJcookm43VhsMSu7Ebgj3ntkg6GaWU7w/Dgmw2Em8wTk5JN4lluO7Slx1W97ZzAiWqUN4
qxA2ySosohtGybA4SjwOxlqFQsw4nG9joRd2OUWe2dY2YvgflE5bSCtVJE6y5EDBOJBgrD6NzETC
RWNlWy/oaNjmK+fxVvjMQzG5RtOsIwHz6dDw6CD82F2mwydVlXzHUnf5IEx+EnTLms/ZY9INlyV3
PT2JPcd3+DBFzSf59ZaNFg5bKxC+OwpkuKktMgcE4G6jyV78M1ZfxqSBHJENUCeRgVzQRn3Edp1Z
XbJVByLNhhqZ6PyBJg5GuKa0/hk/SVJlMI9HpiPTVABuhQ5Yo8SoMfgEzzX65hyeaV+oMpkLfNcz
mqJyIVSgqy51HNzTlOtWKp4yk3eBGLf6tumETG0Ck1SJXZMvapcCIdU6sNhLqIypdeEiDT218awB
T9jTsU5bU33nfgCYor6lUZ8oBD2BYHmyXcSex2OK1rfbyYGVE6irrB2G/+0nhWAm8SOnCXKhoCpp
N0GqznxqaRitd2RkcQmiUcwoBezk0PLrgxyISvJfhnQksRS1QmTfQDuT8F2CFeQ9geCyw8+OatG9
e8bUdk0ScFEmPisPIYjWOA4Cx4Ts4hBX6YSaFw06D/OswEGoezPHqYWCLQ4BFJ3rpGG5NcNzJ+Fp
AGCIECurXY8U1HLa2Q3CIPBd9GMlU3aqZori02WfYkcm4Fj5J5/Zg2Snl7iHhcM1ZW+6/U+woUh4
MJqz4s+IqaOTAtBerDH1LUY9XSfGHEK9+9t16jyXg0/5ISHls05c1OPCoqXdb1r+XjOAYYAHqKAb
s75cQqUGoieBqQUTjYujJEbvoHsvpe0ocZ+Vrx8RQ/n5pp0tMOU0asVCL19iwGoEUDZ9Fp3Pk/qh
0xfXJegxKGsK3V5be1Kje2cWg6t+KWcJWwuHXaHsIysSrhuYxMsS9vmw7jev2AgqCfEFu1GsNzJ5
Rl3kmh388PoQ2s0KuuoJn0sArwDV+wyQc9vtrb21w3G5waMYjOdHPBZKxpjMgNzLPKGtXVVE6MSw
P0zXEf7Bq/pwUZvHDY8rxcjZ4+Q/PEC9P+agoaPfUqvPzRue988Pglvqbk+QLZdJqgtPFsBJOP2u
ElOU80wcgDLsFvT2ls4oNcg54lBLkYwv19Mu2AGf3G3aEQTEGLaHC0WzRJ7kyBJI4USaRU55jj8n
MDkadbAjk6c7tOBJf2G0Jp4zWJY0KWiaQfB69pnbb5v1cbBLQDPCRvnFT6gutU19OKFbk9+F09Fn
A+5XoUQRT7cG9rpjN38+eYctyyVn0cE0An0PtnuBZ1OoS/NJeyQRmm6r13Lk/YHD6TydL0XpsjXI
gUwCTo7zVy9qPuXlGEXtHuts1y0q1Y1TzTnNSn8NJIACN+R4LsEDXJlN343hXcyaSgwcol7+avBN
n8BXadtYIl4e6mLNaz8zOTG6CWE6UX72faf6Nb1eIdXYcaJBWxX1b3fK6xlcv0P9X5tMJSItve5g
EM1yWeiYyZPVrYCRHVy4CquDakwPk5Ua+j9EmvWc5y4LkA9Wo/nTloHF/mZKTSgdRaFu3eGurEgd
zLu/EfnLf793MT/LUQp/nQvc5JYg6qMdubQZEmp9hgjblRw4CaLWIbY+gNdsJjejqD1vzWTz4hYf
2L0uj6c8rxKoPdrgZKRwyHs0lCkx/cbbdRG1V2YktOsbRHBihuVCexajFT+zCHa4T2NPhe8jiTXt
b+75kuhkWCAJwc/RR7O8OronlgcE6J/x8UujfjJbhSDrRetSRlNapkTyf0qDbGPw6ipvUIwjA7Hh
WnAO2Sx7mKgKaO3Ft6f+B390YdBJ1Bd41SZQXRIbri4OFRh7BaQImGYualL3fWvmWnvMRfmXXfUs
73Hy7y3xFz3aoExjPKTNiCqsA3trJH0LHNM9NTknFL8bdVH8fov+46aRyLgdZ9t/ivcnBgyMchfa
kdez7QDdq/8Cyx6NYdflwgbZ9DVKNqeaDznxH4IunrZ5TC+O2IaeMKcpcwNPHVWYa0ennFlJgX1G
aE6wIwLs8NHmoAtx2ceVHpERE01Q9oGnqy1TQdq19cZLQ697VpVuW87u+4rAAmaFLXKbGPf6TRj/
zruSUW16+WUQsIG3kAYGWg6iYpbAXbhE19FyPmyEEVPhIyRhDZR6trVA39yn/7xfHzkpyLL5sW06
hZLhb1FzPv/xT/xBVaMP2f/82AAnGHq7awSAur5hPse4W8QBhmjAZuGAl/2DxeP+uHd4IruNxYhX
L29kcSAVtRLli8WZmTdSdBN/7yMkUhgvTs8r/hTyZ6Y8iriUmavAlXhL9m/xVb93M05khi0gJPHA
+7mHDKv2st7e1/jGkz40D7p8sK7vetQ9kDZUdq44qPFY2GQG1CEwHF2HebQhjfNrSopYNAFW9qJO
hkY5Bb90mSAh8pjbN2z0SLqZUdTKlPUoAxzQ9he4d8pRf3wDt2dsZqXy01LXa5r1QXw2PjgOuT1C
BDQL/fcDnwEjHpLGIz22CC+BHpg6tdKsEvbU5IvvEIeIDvgz/dtw9dFcIZMT9BvS36x8A0JozH/I
ymqL9mym809qCuYbgxzGh34tVg0hsMRqeCtFx5w+LFCqDmzf5CgWYLlSCgFVW1nI69g4MHyE6KSA
tzoGzxL3yI9TMCg6Bkd3MnKTqQsELU5S0wVZOSk8tu5Bht/empGVbgGnAFqhaJHbMlZvPVe4Maa9
gOsh0u2DTBpYijhul1HH91zBW02wK81tWsI1Q3CAp+zzK/UjlmVgoUGmgMmf7+vRPWG5A5jkyX32
T4mfLIg6wWzKHdNdfWSxIiqgYvSLP7G8HzhJN/HU5fQ515tod46Q7aDhArruSbloACyuYILv/yLQ
2PSrRs7pi3uVT3Sc0q//mo3Qe5D2Y1lu4AdHzcmx6nsGvqYgH3vxgJCQNkCw8USTOCfEphoUkuIl
90vKSKCv5sjvtTWePfjAbLGwZflq7s/PeuiPY+hF+5HYOgfluEQeq31/AYnGcypMRXmdIbnhmqS0
Mx1PJQiOc41ZMP4Ig2VljRs5mkjcO2JRHRIyL+meKclqRX7+rl3UrFN8iEBbBHJpFJuY7Dj5PVe6
C4AyeN3S1XveyWhfelP5nHML99ZmYlZDYUQRghL2QVDiOs6ANQC0TzX7ZcoaXXvFfyEz8JuEIAwH
yUNymSflrWDQ5PMNChIky+Tu5HGfD39vunKYbY/3XT8PzuqsuVrvdLGpITtBnqoyV0o0DdwV92oq
wLMeTbirezRcozYTpO71WAk+VnsaNPJlLnSXSKmHcjoJYTTWm/Fr+LjzN9zLiJWheXuAGB7kUyWJ
TVJsXtCgcFd+WGhj/GaAP3nWZCJfCrKZhLlhBEs+V9FqoV98S5ZyD8rAleIk+gZCraPOInZxQim0
NTnYRTy/Uzd6Bo0HHb2MYHdFO4ESiQCx7KbITjEH8ZwBURjUMgB7m1GL0/dz+2gOBFWqkO6RODiI
xQ+ptEV/fRpvzct1wyG8ncdpbnI2Bw3nRzAUCE8f6IGNA9HSzz7F+/Wge/hMdW+xm3vTkrVvBrHJ
qrunOdQGm7bl5EFzQSp3Y5rvgxgLN8iJ1KxvEIEum8TXBUU8DudCgTZFnxPoVZ9z/cqEWV2r6dxY
UiMsHmR7pPObGElGXMX4JGMrICNn+5Dd81jhrbw9z00l+Dim/Zb0weSr+mm/Z8RkE62R59WAf6cm
NzasSqgVUTfqEuLD6/VShLpR0mZ4CsvkAfNjr0quqTLuynJ1m9yCi2dXQCoA3Zru9CHTzMCWmPHB
KbdnxIZ96Xv7mH6sOrGxsBVl9CwFYUaVk5jy+2NEMhSZ1N6wphFLZluY5N/hT8gVzN6Z6igXjYbV
6OM3Xajn4h8npP3mMJ3/dbhNyP2HaOt0jYB7xScK98ZcWw2CzDQLhj1NSbmsf5tcZK7Hvf2JBy3E
cLO0klMjhhqF3l6447HBxhlDMe7hrA3h/vytBCdrk6G+G9f33hQ2mnvdipBZouWmPFUXs2xuGDvJ
MTIrUNzgpKMTMVbFw0HtUBljB7B8dVboVXIfX6q/D7E+RiQdIBhl3pv52sKJ+XvPJpWsfY8czF5J
Jvi4opFH2nnF4GZoeOb+GpzE0F6f2w1svtquf2xtA2wfwsAenm2e6ih62NpSsmFJ9ghijXckhEKk
ue/BBKN+hrDm/+D9SoyTuY9yJ6nej66WPGJVk3CtbS1dANYs9m0t37lQXnTMW2YNCMO7ffRsfhza
9Ql0wbTmp5XSNfFkUd9nR9d4wF3+EO5/kgljGxfL9sMdiR0KbC2dlhdZwOAXhKQ+SfvDitVXowZR
80UNWd744ZNtf9WN0He48nlSQ0jGZm+BiU4EnNRpC+SDUhkhY4Gq0s/Yk43C8XskuRJF5L5RzDEa
pdSWPHvr9LKK6k8ZBWqAXx6ATJHVeMMapY+u21Zxro3mlnC7S8ZwXhGc3Kv3rW7Gy7BaIA1D6WGL
LaqQhoWs/x1ytCUW/6dpploKV5aZ1IkYySeb9A/Fhe86t3AGNYcx2hS5lM+mIyL4c/k6wjd6AKSF
vG6DEbF/29Rth6mvpMV9J4GCxu+d0QJkxjBTnprA2VuUPhhxi3ThOX1zQkJZHcYbsiAkhyovsyl7
v9yzFXbo7bYuqIVtqD+LZqnZ8Ktb69bx/y3zN0e/OVxJ+aaDPXH4558gcvyqLTBXe0jir2jjNh1U
qhPhH3kvcY/G963KF3UPq2h3uWkfrDH5Nhh3fKZ8LPSpFGNW12U68v460EFQFgHXNN8rW9aW4E7z
l6+Cy/DqKR45mlnhS2OShvLMjwfB+/GlTne0fDhum6l16NcYnKWh7e0deOdI4U9iuP5w94hs02ys
Z2MKkTz3j4dayUHsJP7tYboB2BDkDRpFer/0sD9P8flcpWSfjtVJy6dEORgadBJW3qi/hX9XfEz2
kSZ3BsnzROyKB6e4wh82VSqtvrFUFgJrAZY8rFbCZ46Ma54Y5S2/RO/WPuoYhRWQjld0NRAyQUXw
NDsk2IUqhfw8IXGqM7KkzM/JQzS2mZlt125YREshrRlQDEjHhB1wMXpcORItjytaWldLZRQvnBv+
H3mTYAIGUtHIOOX+fQNF3Oxa71Gd1o/y0+TB6wNqQxNE1aKt/y+NzE98BP2rhIP3Fri0apovWCro
FzPtHE6zjO8piqdzUORhX9gQ48UE+rJaglkVpJIgC3Sm8fUu1HyTCFGo+646vlmK/+Pph1q87350
h3+eZp6/HmwpOVukDFIRoOI9TOMlc8pX1Hj3oz306ufsR/56MYWz1+WiwnE9IHKlgL+WPe5+nE+i
3EiXjQDlJjBuU9GeBusPkWkOMjVQloTJt+AXBEE7yDA4N3tARUPOlZOyNPQCPH2iqvsTu9Ien1UH
a9tIlXiLB4JGD8R0LPIf4w3UpKhM+rLiadXdL893UNejPuVcopymQiyglzNdFFLP/xcT1QSTpBuh
NtRdOsIvkBI88lQCQyc6K/B64KYbwgeMs0ar2ygtznjHZbbaLe+AsU2wWMLkH6z3tGOqEZElGqVa
QNRoj78QFeH0gATlvEN98DtipFC++DjqOfvEd1XXj2YkE6rgoj4xgIneayFatvcbH4mWY5QIP00S
42Xq69AZq4AA+B7EsCt+Jdv00rt5RmfmEl8zeik+iVpbdrEIpT6T+y/I/3w+N76Y4sB+u82HcUhV
FXGH6ZcjexoJOTWkvIyBhPXsqRqomS/icCHiTNnCKWlV/oiEGTFUsO2bWLsHTnH22Y58Lz+LyYzL
4lhU64OwBK0zhkchQ4k0rjTYnu2MoM+yiDarjd58bWhM/Weles4dWBA2d2EjHosgMjWMYjftM+qW
ukBrxF8rAM6s7UTrTiKMMRtDpc36F8Uq0Oxp77coZBj+YjJNd+7Kxq+IBifbIoQBCepS3W36Xqjb
P+6fh9LYPOQfCOmfdXYoMMwwgUMt5Fr7rN3DMvpIRNjtCR7apEldDMEKtUSpTxmLpsRd5Pkay64J
qoMj2AUZyns9v8l6xrQX32F4wJ+soDyoK70ScS7Y5JvxxKYp6Hzhr7rjgmjPQClqwkfGucct8oRo
YJGe5r66AixBoMgJIDqo5i0YP0yH7Y1BHmuQiOx1nYq61P8ATX7NDeW5Uw93Aq1h7Q7+4RkkC+3Q
eFlJm815jSyLUEnM0U/3AeodSjATGCMQ394+gNqKwbnB2X2A6si5F3gS1K45eY8oCM11JQEmCtgJ
VdWlI0YRDpeXwhvAx/Z9wTGCMye2YYRhy5jyX9CUerfiBRRsopj2qOZyVuX/o7Yk8uCH++DogUEA
2TDwrLCYcg3tadOH7vtVwPwn7j0O6crgOWdmNCGc5M4he9LgxtJ2X37UWi6HCW+28/QFhVWlAu0T
JiLoq35yA6bxBxS+5BUM2OAFbvYfRUCdilvLDKm+VbYFZ4ZTbQCkNzYyrvFXrz1HUgDxW3TUZ4MU
hBAGx8xjOrItGShjOgywglYcAFCyo9SLwmc2NtaKwH+tunXy33fPNcRMQCaATm3++kpmY6rLWO+y
xl24KuwWbiusB24aLGMSJDCVZhgG2FDEgN0XjY4MTRoCEzUhOxOuf8L2NNQDc/sQMO8b7i7dKmbm
e56uxHkzkUP5km/ZE+NKnyO7i22erhOlNMdOP8NaRYPl+wqzoVUUgTaMtu1oaTwO75ioLG6XIFjs
wvaSQnl4jsfTkoBqgswmJPfFOCnljBu1COXS7x8xNwyVka+lljH4rFDrtWf7pPd42TGe8MjFLIjW
lmSR3aa5Psix5rjq3T10T9y15be9kmwLnGDOVuHis+QaeVaCPOSgDr6+y0ryfOO52mn/bu2mlnuu
HY1RvxrH2Xb/4Z/3f7aOEY898+jJ1uRMAE+ttGTXq7bfdoQ53qCe2ImAHyGGjGCqP1kZvsHJXnBr
sc3Vh7Z9zbPtBff4IHP3TOctp+KtqPRIe52LRfmN0yqQvwzHuicENpE1k6f61fOEflpVi4enGtW1
heqMj9n7D+3CVyi9uEXVii0H1xH+9zwEcabVQjgSnOH7MnsWBXL+AQC3CI3E75dCAVnTnYPQ67MJ
lrN1H4poxb2gBXhfJ0L+X8fQyLepdiN59Jthrmn/m6OZ0s6ffOG3x3ztk7C56kRJEps2t6TGQkwp
HG6MZRHeIrhk//MTELETN7Qwb8zX1dhXLMAIyoNq6OxEnzRwqNe6CWH8VIUwCJ4+DklY4gqsn2Gq
L6C6IGjQCLXYQ7DlTGaQDt6qe+kpAKJRWcjg+08ihkuQ+GYj6UXeTAfJKAtA3iAl7CfUgQftXR8v
ELHNP0lyt8yG30hXEynS+WFOOzRznE34WLLrNYie4/pNYFcQtffK+cCbad+tnFFoh1gU7pdsDeWW
s71pjo7zXSWCUy/1ECTKY1Nm4ozb26tm1JPabAKUW92C7DrDi/EQ7jW989XkTYg5lbYasNzKCzch
wzE8Q6xOqFs66v8PZ84KYuvqFacG4IBngWSfIuWmmmX+/htmbm8l5uN83IYXA7h/aNkhF46MCQqp
OK7mZraaQHog4VaYYTQCLf0Aex/+TUw/HKb6FbHKKQdZKov6tQeNT5ofIAMwwjiikqpcZGsOoA/I
t08F7avt4Src4VGs7nDL33b/YXa8HHtYx7AtMP98Ew1z+iqXKWxsK/7MDigROD6TXT/7797DRjJi
8PwJTXexmrQRJkFI4mOwSubCtTHPaXrdo8lw13EvpxIQ43KmHAQyCk+zWq852WCOppGl+M8tXh3F
JRk+On3bwh2lH2QOEsHCY65zxiI0DU/plBNg7fOJL3RexxAmVd6T6LwVl1dR2fl1vlfuV26vHSkB
80fhYhQizAoOFyN7NF3IKlQq5BqGbOMfPRyx8kBmUkm3zJC2/ccTP4Ej8tJ4RjHHuimRIt4Rpslb
DX56C1Cg7UonsMaqZrtAqBp3+Y+f2VutlC7gDpqSG/9Icv+zymmCEWClrnusQbjGX8WNptIiYvVz
GeVWGBX78eyE1U+kATa8qzmTcV1ulFeBtpuqCmhMQfpZkS027QUcIkQK35f/tNnWs0VtaRu6VlXa
WIHYKmR97LEeuhznHLyiR3nZ2HEhuFm9ozzsIsG1w535d171buSZ15GOgyAix7WhUXIxXqsz1rMF
OgnrNhrXxKRnPUKO645lB8upD0I2qJn/OvC/TcfL+7FXxq8OhbnuwmpifsHfUsCSy3aT3qMVK56u
MU9EkW3Q5s+is382ckLyNPnFCYoII7hEO3do23bzvE/9GyHjRTI6UZOIx76B08FhNFq5bzvgeAyg
3XInuU6LDXAXgz3Srj/lDm5yQ3ejWu78MhjaS5M3QawSz0RDVY64FTKJDhext8qtkC1dL8+JRFHs
OpziI9kpzSHWi6BBmFlbGJ2wKfE1egxrowlsRTHcu18qYzxCfMXsBSXJlmXrd+NHSJb/aERPLqhY
aFqJkbdpndY660H7rVf8ejBsnwVqr+wKJ+zWG9/3oJSv4LrtUhhc5Cv0vPAXGhdcGjqSsT6SeYSN
lc52MRDQCMxlq+R54KPUX1CsyYe4NQJHHOpUESWdkjn18B2eVDsmnhO59V5aAdeysatabJrNV1ZZ
3QbO8ibNgDKQXAnq7mkFN1tbJtLPpS2wDiTW2wqgZFmmdwuQq2yD3KAac/G7EKndlO0YOaQqYLmw
MMlmWWn0N+HzG9XOqMZUJhW+ooqLy6X8QAevkg3qdOz/0OJ462K/aQtIMVYsQR7x/vjrCe41gaYP
k+RVe6f8lZZI+KygzAGWH3iPhCl7HzmN3L5dh6P4xeso4uOn5O0kXKmOWRSPuBDo8atEbLGvbU3H
1zm5PaG4ZQmy7ReKAFDB0XbRb0ZD8JOV+whK+nQCADTxuUM1/fIgSCzYe9TyR7FYw9X/oJkLaGMO
4yDvHbKWpkgBRdgX8nl4S6ZYjF5kKjFqNo/Tua/WfLrsOqrVfE0hgoA+rfAFuXTWbO28tQChybv+
i8Et1MfCS7KbxjvC0bch6+as/D5g43qg7YuFaMLHcpsW92wU+ApLDQ+FhnRaBEaYQ01gMSCpVpYb
oSkyyIk5H25D6DnNyTCEc+q3H0NsJ8TGIgRItXOkap6Z2DS/PsBixxql5bGZUFZmVkw8oZ6swAPl
0z5jNSPR9NvyD0Omh/Bk69/ppFzmGn29tS4ZOptUkkUSCA46L4u8JhL7MzenlrjVwTk0aOHeWb01
QM3xxVu7m6tIukeGiAMeBdcuNu/WDSwe/65jkwYUTcg3j/Hv8BFhKBWNVTRostzlp8kCdY2GkK8u
j2pO+GSNY8PwZMdSlasM4yVK/G9jx38mXW1xDnpcYigU2Rw5n8FFA8CiNBgpe57DI6IuZ+wDbciv
LkxZrFLWlxmoM4LgV8CfdIyhyZNHegclF0SSLVSSTnx9MDe0dPGpgeCBHxHbdjNcmvTCguK4DOsp
wXXWVK5kJNTKlR7yVVn5svaZPpToWKKQyTCn8hvukDzCnQgc0TPdXk2VtfxUbpJzrCemX/8W3E0R
mUtTZBiZKoW2n8WkKdeaVgff81gp6joLoccPUKp8RDYJg1j9t1NkztEyvTb/RTOncgGeidg6Vbmd
hNdp6s64Q42Ki4ecdiQbQi2ZV5JxkwP8ldlM/ehC+AcJZSD8zzB/dwu04vQADvbp5oAF77ly1bBc
OX6VgNedEIa3XuPPLxMwvREl8rYjcCyfthaoT7IU47jf9vsJEeNrvzijTL0Vyl3jJS3FWw9not60
o+4eV6U0PG5BjjqP+OogbQaap94tQEJ5U5EM7EZzMVGkio/8JH+ytJVLYMbn1Il1oEbG1pcVnni7
Q0hZ4a469kurJjIwbQWyCaaZDKGN0ZMHvYgA5CZJKSp2/2wHA4oSXH1usmf6ss5WYGtdzjp5oGUF
FLb8fSx8vNpZBhvso7s82aBINvRAxm6VkT++MC7/CZk2BawH4l5/eOQQRZIWAQDGW0Y1qZN0ZC8g
tUXRe2AJGIS5f/CWrppu8G7fmS3soIr/LNv2UjAbkWWZPp1JGLcoFisvG6yuuLFjg2Ct49cRd/XP
XRtX3YGKtUMjMLRIpJK8ML185nWXDg+vJ6t0A3/CvTBA8OYoJi/Ksu8TdjduE1nIQ3vs7AjHPHpB
zG3w3yX3U3hKFerw6rjrd3ACb+TcKWJK4KsXU+Pz8poOz3jI5qi5EfjV31BUHVekxqt+xhS/H6CM
n0XFUUpsPRKTKebGy3QRmHpI9QK2T6wpK7nGXoX0OkRVChV9xuo3E4D608uawx+Wdk1rg5nQmVoA
sBHmSO2opKtmU8L70G/H1DuUjYByF3RA+LlkAiOvvBgiB78lmnNB0HmeacjLexqkEAYiPJZCOdhB
LYeYnctKGR4lOCI1H4ovPnq+devQ6jmeIzXUggqnFW4vAoXT8ZtcVPwUrq4Y6/zsEgdoyPG1M+lT
3iY3pV66S4aKfb/bcChARDFIWioyHQZYrTQMCxgIGhaJr0yYSytv//rGotOxqJFF5hTEPo8dMyvH
QW8TQXi2ymDCAZFX4dMmtVTcYkTOPy6CpMrnElHOplHWpzNPEMk2FJz3MU1T441fwudhXqu7CAPX
TpTremf+RBvMmbDbx+OpLKkKtofrkHukEPFscZYxz+drk4jlRWg4Z1X0DwAKO+XxfkCRC0cqg8TD
GlbIrehMTPm6KFnmcsTGA9BFJHIK4NsPeBRFPJWD4IubjVLcmchSZkVLEYU5/zfPLKb6QRok8pM/
Q3OQZrdK0om2ioyIksmnntLhMzZpxKCWmxZr8i0tBXPV1SlticcRMmKXdjyJ5DP9c2Go9/GF8BfF
uNxOMS6lIkI6FEmMFGGOgDbebLdzWjFNXNfcPZ3UlHyZifeUrsptPGlJkUSaceIy5UfaG5N8ZuCl
9d0BMvAVEKHjipmYH37aicx4zsS1EOu/Lo5tiuOyUpf3w1iCiw5etbzWVHqLK31hj8qpm7Wy16mq
EoqXe9MM4OYXjRnoGqzIgoaOKSEIU4IjJfOg2nhdMPIH/ThDdsQT+AZX7w3X23Vqaub1TDbXkPxJ
KwAh3PuArLJ7NQmNwhOiZo8RzEM31WzwELwCLrMEZ0m/wHEwhxtZ6fDA9aGAZdjs63o+Ef9kQMEi
RwMxuHooQof2Ej1XgelzSjPDNKj/i51FpDLsrcLVa4jztKHIUoXwqXF4UvCEBTBz+3nUs2qM0CaK
3ey8NerwXKoMOR9VoGcNPkvh9FX/X0v1AWNKtm8TIVfGA8FqCbB/1SYL7vQH8KJo8KFtWq9PtVq+
sU2c4xQSMnewvZXohFs9f1Pgx7U8COQND+r5EkW1gaCa1/W1+7kYP9AUoLqmo17s/TrRkeiPW8Gm
DgUMVeONTJCkS2D5ygGqKt18CT33KSmzQE4MGjYP0BfTkcFLtw7E1DW+B5QAnDLW0EDU9tdHzSP1
AFfeGnxidsgPYsM9ZZhnVFYK50OCVDpdm+QtAtRfWz02ebQAIFI00cIgrp/zKbyF5DNr4nQXiSL5
q0S268svJfr+lwYGDcpPkagzaEXFU89CfYAjlsKMk7PF9CO68LplgRGx7iMd3xyjuAAmfZTVfasl
uoIaiQ5/0sSq6uEnzb78Gotg9zX+B8zgDaIFUCNbhRODI2gQbn0CU3TEC4pSpm7X2TyAWCUiibBf
NL8AZeb5yJa2DHW220emYTaW0F3yqPboNQYmNS79wcmVH5uTfzQLA6FdhQJ2DrerZlN5Z7d3kX4V
M/Mw26x0YQIKNhhRRvfQlMkMAfMJjXPW/1VgSCJcqo0LdgvjY3VheQ0brDRB/NiEoXPpWtVVojMI
ehOK35Q4YkiOuikL4K7m2K8DSLzicSJiHq6w+i4jTQDuyBgMgR36vQ0AIS2njFERVrH4JSm6v22L
dvufuJRA8SQzwpVMVfhLgHRjNZarSYNl98MwnfjTB7YRNLCfJmAczMZ96GROcdOJB52BQf8y9NvU
32Bkw5sQhkRwwDbY7NvNJpnuEJI58KfmIf4YVHTQayXUv3vl/pbRXf1dlcbhokC6gOhvE9kGb9ve
gtRU1oK6tD22JcKR4H1L7uGH65AkzdEgYOdsFJCFkaVl7nYtf+65SroSOvuANKic+plQUE84y4dQ
jzVyRPlPB2zp9zWqmI7V/StcoAFU4tgZK/1dopaiRZMup7eIUAjsSpPCnAYLfozEfR0ghNh6ADMi
3MGu00kN93w17bRsjnJC5l/hkfoDL1nEnBoIB+sLJY/Mu4+0LFN69pxtCK/p2oYQJIs+VzV2mRYC
/v3NgfsemnSCR4cqbsmQblD55Q9rY9bhnezHDY+8+t0qG/m7PHs+XjFzoTUoy4C8c7mZyXlLjgog
rLp2w31Ou0d+zTXJK3Oznu1AgYAcnqgFuahTAP2fIoYpHSIgTf2OaDiNBeDl4w0iWTRzVk+ariSd
0wkQxv1CoLCrcRJuI+Qkoy2Jg1Fn999zUVgGEpVfGzlTT57goxVHf1mBYAv7uWZEPoRcu02lee3J
VSHL7HM1vbLPtsBFTaVFUlnkgdaLOfx8oVzBqgfXZcqTiwMNalk7V65Q8HtQz7PW94ixAXztxnIk
PCc0SupGdGa3deCiTkHIFgf5x6YgA394W5GV/XTfMAgaiqn4MHnhPoymVLdyA3i2s/rPf54QNYRW
Ex6ftZ6DlaJWs2gznQpxBogvVuZf3Zw4uBgsI3F+g49zZHk7Z9AsgTA9KgCdCxZgnHxRFixUsuyP
mzF75TuI9GWMuRjhVBnE1BIZlhGSWzzVwElJeEBdtj4Nb9I9I0V+x0zzOJfnk7F+1ePeY5fWbocv
gFcOPQwZ2C7M9NmFJzG8FCmuAe18+cQ9TO5/f9iNKCpI9A8iFTATXlkn9EqqCWi0afP9SSXCdMq2
RfoRVm0t6EnByIis/KIWIUVyiK4gGRedWgWXo4KVCfxJSg0e+2Lt/p9UPysy1aMrRAVGE0HEyEcS
ALmfPSGq7jOr0IcYuIJQ3Yrm75JpTkIB7VC3kdPT+smQXMUtLQvP13K0XyCVD8pLObQInFHuwIM4
mESM84ZbLwWSd/61dFb+ccPDa5lLfdvlOWNFjOe9pN3SyphIMshdiQTqMyDaVj3J5t8N78nTbBN4
YWN2RljnOa8/5uon7ekD2b7n6fpuB0BI2L7h0ouW/uuLieD0waCC653cdNpHvuPbp+plukkNXNpz
mo6vd2us/N0dhwGYSFl+hC7Yg3svyTzg1uDu6rVeFRQS66ODWT3kPfmBQlaoxu7duahzbMgNtKdk
KNnO6donbOhf/AMDl4fcJVBBZtrG8Q8qKDXyxUH1neHhliAZ+rsB4IqL1jn6DDtJ28ARFmg68nLV
odl6WQVBBwPpjbc/qtl01EhflNrwNFp/jDIPqjWtxzDG9liS8p1scy+kr15GCixuaNN90qo0jVPE
pjuaIFzN+ADiUP4Ha4oj2N6VPWtD1Hjsjkq/MWsLfXi3VwhKQHnKUz8i/2pRIkh0I4W2MGCzXgno
FWxTkB7EsYJS2TVqiS5FqHMpbeve/vGRC24gWcDnEizhyBFKUARTCvskz90OmceMSrEzvF/h/siF
WVlp0i76WiXIBBQVGRbePHx75VOse3nLlE9N4Pnvdju8ANwTkiFbr18Lgq+liu2VAi6cx03HJsSa
zPcAowi1ysxldSDTy6lPS4bjdwZDjiGlQX9GpthGliKYdGcUlt93zQRuPpHYkrbQUg8FRLDqVz9N
FoMpE5F35REWVVRSr+yxsWqsD255DOQNXF3kWNbqFEJQzm79dXoJk33DMEkJnSlzwFmTo/guGtX3
eq5QsFy2VHfFKVdI/RiDIx64zcnrMAAWTD+lIN2Ri8sVBZVR5ABcSlyWs90+1MyQ5SA2XI8MnscU
fIdLqKY8WgDZEoZljsdBhruyKY8mkgBfcqau12/Qe2gguCEbvny5OYtXBAjw1TiFZ5nBsvuuUGOw
DylPwY+fKGxZ8rMO1ReRXR3pYiZlKgMR8fVRqEY8jkWLjkx7/pJfDrIyLj+fQ1L1MbdKCcYHZ6/r
kwVHilBzle0+cAMFtqpE2UA0Sx+kD37yw6ju10XeXm6qyGyAW+XkwFz6HZLKZM1tLVvJLBUuS1KB
/czXjxU5U5vYPAOL1lguY8WQtAgQnsSIRllBcRvxs23sAvNRQYnjjl+rB/o6eQcE2zp/F8Cil4yp
K9RvXvXLLtl3LK4MF6cKchAsohFLBMndo590wxD5BH8MpaM1sXYP/BGiVuBwRhLSiwFL17+zL3vg
TzrFM+zSxt7/jSflyKyNfHAiLf/IRGBy41PKM8ovyh24NVNY/mdP4OwygClAkNKTYJW93W1UANSl
Zr21swswQQ9kG6FrG1KiGH7imrtGPqKJgrsuegj5DGg1EyKX/F5yUTs5ZKoLC/UrkxpTVK/RFPhx
yNcIjoX226AVwt1de43aG/SKcUtdeQKeE1Hwex4pEM1yIZsCCJlOD0o33Jnw5lBOFfYuUZ0ws2KG
YOYiHLjfO9/Qlex26KSnVGKLLi9AG2e560xKmSXQoWoW6cyIxcvloC/0Vtgq61lW8167CMAagn6V
1/yJ1LvPHdhMMtpqld6gtIxQIEOeJ/G1DFDw4uYUuVrKarIgCqKvnj+xmFzMUSpSvypj7XXO+Iq6
fdG062gvfYC3d9QdtRVCmTcrfL/NHbYLfiRUAUVaYKFRfU24TjSAVLup4HqFIwV0AdcGHOb8kxde
EqlIaDo9MalMPbZlCuUfP41FddRL7pKlR5Is3SyxXnOoBbanT7DBJzyHOxEkDv8JKokaaRo2jbEl
la+6AITFeVYRRKCwUuNMSOaHqnPZju5vVr6CrpS2Dmo/8MxQnPvYPB8jcyTeaMFhCJKnxD2+5YAd
WOfE4HdHFYOd2kcY0aLr7+aV5Qmw8H9k0xcW1p/Y2Z2kLKwf/moBOhVLpWcheJnr5tLNtxB0LZBN
uED7UVCb+ma/5t32y7vtM3lBYyPS7Oo/4IYwVJ1Fqpgzwy8LrRRHaozTsU9O6e8676JsSzWe7AR6
foJFxw70A1xt04RRF2xE/qKx0kFG08POw5tKSvAvbzOU/h0znZtcJpP/8mFVD3HvDeO2csZATiuE
eK1Z7t6CsWAgRttEI1+UlLQqLPc3xZ4oJIy0i7Xrf+4+S4FSpxyYMt1p0U0qARRgNoG59jc20yo/
K0+VjBkWYD4kUBuh5OBittKbOIsze9ThZysgnbtikMCTYme6y980eSXuhkg3jU7cmX9Z5IrCk6sm
/1Nf2Tx2+lN5jIPSjQOtL6/gNRCoFdM+pzeczrRyyQmFzu4kXNYBwZJlZzuWJrDlCIBHbZ0yQUh8
erauZCqwlKDatLlPiD1CP5VfY1RiQbOQ3rPqHBKn4cYagiHrxUZyzXISqZz01W2HnuoBmUQhvTzG
7R76bakEkHdU5NVROXl1ai7fil/Z6SKUypYPwwKaXn5oRwKjPFhf57Tj5iIcMIotayRz8kufIx7Z
BgwUHsHSzEwISKeKJ0KRZ1zBOeOVeGcPjp6Qyj9o5KPzOMNDf+MwOeAFEi+36X38QyG2mIXlnry3
1fTONUz/fKy6FQ87gfh5VID+L4npgQBdfieGeivxOjRwk682hyT8wLcdaFitJOXsuQCORkmGVXDi
6NAvnKxIUijng/m9TQWDV5ybVic/9/EfnWeMXkD0HcQgdIvjPBkxMzZd8RC+z8q+zaZ2udK1BoRx
2EggUvhDjhVFAmvox0guwDrX1TsKfqAxyp6rnQyua8IJTTiy4Z9IuvEJci6GAFoDyasGEf4MiwNO
1Euwcqp8uUkotKTRFxmywszKuDndi/CQdR2MZ13x0ocF8xvlWzp3Kn8PsX6YyH3JUUkL5b/2FiCY
cffXJXLQ0Dl3+yQ/5dEqewGpXnF9XZyaa4hXJLbAPThRC9mEV7O38JEg4P05BaAqbA6QKcfNNzFg
JFEFS7DNV7acLQNE+U1D3U78HY71pwTB+1K7gfmYjZ75nEgk+Z91FpEVb6Wiou01ZGD7TLPfHQJE
Yw9j5FXKVOjRl8fF/cB0In8VriD1vnWF/RsP6rVcYFPoyX3rFH1qqwkLx2SoN4yJujQcNNWw2GD5
ymiTMza2S9sc+YAzkqgmO3fj9UO7mnJO0fxn3hpRIbZKT93bBaKTU8doBVVyWBwRAIP1AnJ8CHbv
koRE4yaR4/mhzmB1bZ75pHBWq1s5rsuQpgqUdUYqZHnv+YIuoSOZpHYnYzyB9VH93tfWgPG+EtyH
ai2yKhd8mfBD9j+/u7IUiBPa4flsAODTDer8LIX0lurTBi09Ucj9sFk2//HBq1lQoOcDldZ9XPJL
6a9wTkvAMMWuaS//zqMJjV+5iAjxJH33B+pcG3WnG7sRqFqc1StghpYLI9TfRmPf4q2cWWHgvbG+
sd5oRqYwICaaXcW6izwRIprfdIPLy3VmDbp8/21uBO5fiKrPbNTKtu9MyA4D8L7lNCb+bGQQtN9o
8XQXKNN/hBxSeT0N6NMV0vukNSLozNr2sakKBHHqe2ZdZHfYkVlfFBelvcZWq/xx7zqUU30YPQUh
iXX9yI47JW7jykeP8bwsQ+Jxpjh/sQYONhBzk2bS9Tr/91P/IAZTia8h2ASlx05EGqTtuDQxqz2r
L4dJjbsRs2MIdMdnekmJpaIqPUBYmhCzTOmQaBaE0nZUPGFEqmh5IOzN+TiWGbgZ9QdSLutFSKx9
7ZicPWgDCsaYaqu/5UM0lh8mvfnnO/26c9hNBH8CEGY8XzjUsxpWTTKAjHSpoDcGINs/jDO/Nuuw
lvM2tJL22ptFB4fJzuUhYOZZ4c3eLOz7eg+zMGB9SVhaPlQrrD2p59gJNFrUyai+Kjm+4ONGZOzw
D/ZgX57mI4/s0KTOsNRpHooHzKctL7vSfPBIhlOGzBz3eija647JNQ4g/X/TE7vfRZpeeXWFOSBa
WSeBX9LKXxDbji2VuRmycYqx/OXcta7+u1uLvpaG1b7HPVQnmw+fJrU93MkXggMqoy02jA4eHNcL
pmNiDiD2JXiyvRlwfBsb5+9csWS110viI/mre5g+kTpL2eyXWOtK6cGfDwyrERwR+7I+RAotBezd
RH2gVP8fqE/FBLZWxcmKep8UbctIaGzVpceDMNRRyxACvqP3VW8xVRlyak0S4MMlsW5hOYbjw0mF
YJ5ZPeaAD8+WHKVn7vGeDpYwgx53P2FLtEnQIeCTUt4oRhzsHSKy/KkvXHjIxxTXbpw5F6ZRh8ZQ
X6Z3uNXOzeHXQRrBbP2jD+uZ0edUIb7XeTCNevUVchuQeGiphgitkex2Oqf7tj3CRrlaXQhSTdxY
nscKo5gTsUybBhcKUWz24izOqyUkA6zEbm2TFpnb1WTHCx1B7GuIC7bJYFxXC20mbVel7rhEmIBF
Py1sWnjZ61VsKH2d2W5/9Vu9YVEZz2oZCRs6HIRAt+nbWdSM5C1uYz+XlhNxf4vPbpF7atvhRT68
8q6j1jCg2oiEbMVKNGpEYBDVOLBtABT/+N3S38Bc7OIQhlBM3PirdyQltqOu7t/WptDX+IWPPM/3
z4ogtscW/5O6Oq+K/uCIHrW6x7kegkQOfwqK888b77uLqr2FpeOY/vJVUxRIkXPIkpvxldMoabd4
mWd79O7j+1SB6jOcHiIs+Mcr4xdhL0z6OI1UhFyZdVHD5XPzPoy+TIPGd7FGbFLSwmNbXOPkYNWS
wamubowT9t6YSRiIqaqC1Gw7WKabCBr0barN/1BHd6YeUG2O69aCycIq3WQ05Xnhdnn35HpJpFiV
q718Gxt9VYZ+piXal+bxjgN5LLjEzZMR5ankdci9mdUd4etl+P1r9ZsdBW1mcjx+SymsOviEPFDi
graqGOWxj082aIrz8h7MKEYHm2PBMzP5LcWEfiQneJzNOe00JBM4JHUHUrKVi7/RvynEzTsw1/NB
rFGb3Jldd0judO1uGQRdHJqEmMR9jQSzzLLGCs0GV0M+VkqwfXgA3C/AeSBFgS9VQ78L7d5wLhIO
FmQC9GCl4ZzwF3WmOJaBzqnlr3FE7B+YzKjr/+Psox64nLsDDmi/qDzxiVvhyFPwKSxfgozwturz
aPnJ+XP5eTdE9q0s+p+PSRLp4ct4GosD4zjX7kfb1u+CpzP6ZI9X4fqpzw4QHRq0wh1KK7D8lift
hUei1h58mxwcTHAbeMeM1z6n56GSGEs/GBO2EjROrcAhRlv4Tye27Te4ctCt1Q1ptN+5f+zagRXA
LNdmrTcWeKz8jYQdjrrp0P25EjK7a2kGwWIAKN5cB0MZkw3hGnX4qm4ZV1l3dGmZ69a3tfhZ8lfI
BgilyEcsyiEimTi8CKkXJUy3eFPzVT8ue1bUCl0nD4fhs2GilgcBTv363oVOc/Lz6NZIgD8bNb7W
VKcBRWvdvoUZSgQwarf2b1aNdJT0IXX5IyQWrC+3IdRG3NfgyvHb5ZEseE4Qw0SJo7Q7jaKKnHah
85cgwWgU2VZUu6YmusGt5H0pmYXL5Gj+xN3MNe/g8y7G5cu2C/QbwCSEV7VuYzGAoO6a9FVHgSyY
764CtoEkAjjVjtvJqR5YXOiujtAzsPhXzgFyLo1Ny5iFQnOT1z6fLHcPy+hw+jGsBcaTr9bhL10o
YuM+JWGNIIeHzCHvG1NtcYqltkF15z9O58VpjLoxseEtngIsjZrmUsU9p9Pc+fDvGnBTrQBdKDJi
hMRYna1L8Q7UBTmb3T8RcJFGPo6xDR335MAhdwN6AoRE+Jti082TRD6Rqq7N2kf4L6Z3JZsvUKLJ
UQGbSVxJxgisrSpxh2PaK9CNdjLqmdwXRRgTs8TqLcXsarB2JG+ovASJYceG29rG4uxfv6fNX8So
tkDG44VfUCvF/moMh9elq0fQDphRE5VLYxXOgiUjf3TZyZKJCdhvLJ/y+8qngq6AMGxRQWDsJ18T
FnfcfnD6n9BrslSapGEnYUwq3Xd/uSan2lqpPm1nSjHAPSVvooCpsepm2vLUa27NQtya4ZzhNN09
ZcQ6TeqnVm6Cgzuo4v7SPqfoXMH1FvoewLoKkRzHvf5wY23OI4B/qFnrn9gez/kAF4Va3QMPNjyJ
Ugcdwb77OeFxNgOBQdb2LEKlYdvnH+0BRWlNLG2G3KhtuGKe53b04fpk/vb1Y7w9yqa44rffgoev
VBcH7BEr2+yiCUeSXaS2M93e1+QkAdpy06qoUTlhnjt1OSsuKriELrRFy5wtTicqEOx/ZrcJBXLf
ix8pLKskuB/fS6sez2Wq+Fhnv59LJXhtJHC4p5aBXHbZrEqmyZkRQSq22jm/PxE6ck5dagi/FJw2
53HtmQ57xS+CEdCMe+dmzv5a6XHys1Vfc6KcZALMjWDqPbcLZOiuLcJl6CkkyAP1BGINb3oKgkAC
kBorv79zLMQ3S4sSptYcWsNdqOLTUV84cs+WUTngJnvCAMWzk2XPfLRaZr1BAycDDACKIwvzqHk8
yiUFgcHX2+d286hrmAIHne472fehRzLt9MIdzwLFynJ7x/ScXCwpnB05TphC2t5X/nozGGpO+Pw+
E7d0xzaDwi6IsY2jkaS4zJEMmC9a4UWq4B/Q4se32eCWAxDUUCL6RB0546NAjRvL8XG15U3D8wZa
h9QrlEu91IYR2Tzt4OFvb1R2Yd/xW6mIXjZ+5vCepvivsLu7pns/YTXNJcbACQGnbPuEOj0yzrCQ
2XIX2Bq92K6yoGDjnZg0ZAJV7ZYubvctW8oG1fizBzZSipb58feLN6Yhx9755EbwC8TAQ1/lj9bU
XKVr30hfKMbDxE8QJX/jy3NwDPME2mW8UGuqsPx9k2pbmp9Lrz09LaCbc6WaqVpmvJF1BR3Y0y/f
Uy6ZKxRW9bluQKC7+1JEGAzq4GqGPPhJlAcJ0rfhgDt9dDBxoYcRgFUrBfj6U++ih3O1WhcJJxVl
PNg/OjnaWC24jtLvS2jC/jpX5QB/g2ayOvPKx18FKGnPeIiY1JULs7jlwGOym6uF+C3eee15xjqF
MGrFa/vw8CPzh2/oe6H1MMubZVO0Ootr63cczk/903IM5YDsAgXazsdKoD+sDofo8KzGuGVtcfzc
ieQYvqE60BrSE2fIRhDDfS+MwVOeQLp/Aiw8d7TcvWsBuw7Qr+TdivdUT/H2yIXbdVjssmtotIZ4
TQIsrI0jTk0gC/iYUgxadYQhxdXa//BJcFp1nSHqSu/B9YSZCiLtDTFscTK4aZbtUnHZjV1sx5Lf
AHOc6+iIWFWkHd8ustA9NoBoGOXyguzsBar1oVZ+OLuoUyZI4K/zYiBSotxvnpJFY8FUcxXjvEGQ
aoHhlSLxcQmomAT/6hlZFgQqKzn2GSdtTR8xYexFqXRp9X48cBORTKS7D3dfOLwDgM4Ld0Phrd2m
1BHV/2VUOPsIeooDdH7lOIzNWxKfZv6tHhE5Qg6nBe84quMlV/PbLYMTILI5+rQ/KiXBxGjTm9SM
gTr7VZuodbom8MPN+C/I2/tt/rPJfZl0jlKUk3/UWdSekmfU9fTRr5iJlQDjk1UXzeI1WAzJ8L05
50l2czlJXpYMOTLycexepb/9TuO3tJzryiZik0t1hzH4t9XPqhLy3sEnq0nQATTt0UethHg0a3VG
Su/rszFfOWEQPJUIejdYnzj6lgUEiavM6bz5A37t2HafeYN7Tr5l9T4dD4hsErB94P4VqZVpB1M4
XXZMN0gG++Na/bhoZHjlaQpRm72x0CwVZxYjnGSc2Xv/gZh125O38CILkkF2uSX1MtVtfjNjv+Yk
U1Lq3xAOg4vyMeWgOOoPiXHL0LFdrvR6j5/PvjSyQnqIU4nqc3Vj/3k6GLr6oTQ9f3vAH4COtWHg
Iniv4xJla/QB/TRxuV+EElnx+UDm4DENIhEaWwadWmG6LIEEfnr9w5Dnf3yRzSnZ8kdNE30Cb38q
2/ucnhqGyuUYvg9V8QTI6EVy5nDf7Fn/cihqxqq/IQ92haUOignfHFmDKhdSn5zvXtlMGeeePlvt
yrFvmoYAK/YTE9v5nO2XMRAWs+/AZx8GCA9xLDfeSTnDHwqPRdsCUaj4t/ReYtX45hzdhhCKWl01
QRBOROX4lCyu+NAyVyE7byU8pGMwMDGwYvSQ3Nu8UQULye+sj979AWdt7xkTz4b45qfFPymaUd8H
4bpk25b73KpPihF3jC+9RdoSREGxEcpOTcboL5I0YaRscSXQhHvfNu7GVO0S6rAIRA1XBvntYSpW
L444ua4fB1MYI6TT/knxgW2FXJAQAHobYih6TxeqUNv39p1vfkLUQipDsJIBb+YenZSvcRE0RopM
gZFfu7nJEmludFDRST+eVCmmOuCHjIf/63iQBi9z63MiurAZ48rNjP1SdZQEa2c7wzdqiSceio3h
yJ78YTizYvyNwSOR8auJjQJfJGCzRMRh/JmHtf1vZpwwG5Ps0IPBw/V+adG3K+nI+ARepM1vewu9
PsDkmpEJMNa7t9inCjD1i/E0WMNMw/TEPbdUvaJ9qbI1AFreXGd2z2LNJySsUr3LxNRFTW4DP9a3
UHXIqaYzu++Xm9u99qIYn1SeJfnKFHCA2rdvejBW2lJB3WJLJl3sPfpVd1Kwtvj5ZXXERiPPLilz
H9mDC4PhkyHDZjqirbckjrxr0rBFTm3j2p+QMy9GOk+HQAJL0XPp5l8fuhOZVakvqCiD7m+mCTkt
IJQthQ/cHqWExWdH2T/JQFkgWJUVtuHfwqrJiHOWanKJvfyX8oLl9S59y1h8Kda87voxGOosvkac
kPOD7GNHiwOP+H7CdAmnaojN//xyK+mDSR7yfQFK3d4DWc/Smk73NaPuyqbndslYOD0s9hz0WHoF
uTH05/opmqWMsXzS1dtU5qyqlviEHAuaKluTrh2o4V5xjz6Zj9t7WmDAF8kyhtFlX8SYTDgw1CcN
GzTEf3F15x13qdqVDo21D+q6T2niSDh6mn0Z/1fv9Bjt7L6nUyP4rJyAbTY55Zgmpn8YXYTVU38j
Ym9y2J1YQqjM65r60upIBapfxn8w6sEE5poJdMi36AKSYPVWJb+U7+LeLqAT+QyiKBM1FXMBbXP8
yb+S39Z4O9VszMp1ekdsnWSU21k/4Z0mX1ntTUFOaL23150ATMCs3WmwLTETQhkka4IoVw+NFhNL
WU57hUTBJWKeL5JyKi2Y/MJdIQ/SKmAzVqsqSmELMSaM0I5DatikYhgisWVhSQjVhlYRyuymP7jA
OkC7HVQRusGUaT2cyIcUPuy5TVdk/M3zTgJnMSK0RcXpwgi3kAKTojB2kPHAW/mLc+yhsP7j4SpK
Z91TqDpcQy34wps/slDUkngtbwe9C8O+Yv7zqpzuwMABl51cz5Zrucz1i+IMjqAIYWJ0YZMpEYzA
I4NQ6nTOD+CbWwj3F+2OMBgbH5J1cAm77JC0kAgtPWl5Y9VQukEprA4anMODTNF8eqgWQwS40fF1
LF5uzp2xHG7oyJsu8Nsev9oKkQ8S3Z3UUAJcEWc2y20LpOfpQCrEFcAlG2z+luSAvpDXVidfX0iZ
HvZ9DOdHnNOIzz0ZZNIWUyE2c8DGJoK0CxCHnv82D1c/BBkc5WdvkYBB4hmIPsu5c6HF1wjU69gi
cfppztKjfZ5AVdSqdYTABYqnacpn6I65RyRv8t1mbZb5Jcz0iO99RZtEG0PBIjJ6auuvljuRLx71
EjT+HZEt3DhJ0z7Xdp0GSrn159W0r+dq0SKKWb7LsTfNVaqKnPp83W6GqNECNEYqFL4UGV60DCSr
/Gpht8xQsCBqywbj2OmdsVcDyKG8GfGduCYGUFiHnhD23LfIdljHousoz/PA+uABfvNxTq82sWE+
edlCXG+RTV4EJdH4vdwVMduht8IxIIYnGln45Hnj19GLGepNy4TIKeq3Jry0Nh02MT/NVXUk4pIB
QwVcggz4Imr9y6ThVIxsHeZG2v3EdYkaPFYAIoHx+kMR25LYoJIP1GfTUmY2VtbPcvxigDkdApFi
JOZjcaTtlo/e0VYY+IcfuJcYxpOZr7G9XGUNAR8GpaZaYT/Ge7ynbmm830bCQBB9I5gaBwxWkxdK
ljtjWcc912o/hv3GYZ1Tt7JV9nkBbMqfcHqUe8/dcx5fZ7g6+Quu7IBPFTaVp0mvC66rUVYUFnnN
aAG6FNpwq8ZjQtr3gkeD2N576UdgL28h+L03AE5/+TkazNGDikyTjJyz8f8b2cStte5zcMx7rV7m
GM2gmKMUKlrUlQOMg0+Yc1D98sPVqIdjGzxSBZaY4kIqpuqyaFwoe+h5u8Irtv/j7XR2iOqV0pUv
CF6vUwxoKhB7hTVQHa3V0x2uCmXfmHCP8nfTZyT/2G9uRu3phDLNtrMXli2KHmh/55d3eGs3M9V8
unrps6lavqXLqU2fPHJgf9ZdR69BTrrV80Hcrr2orz+NxKZGaTCkp6HkSQb512fmjz1d7paYKSy8
Qyq51p1VlkKVYCQxUi9t44kyJ/2nK0RK+Kyrm9HLGaI5lbR7DpkAEw31p7jA4rvtD8Q9iK7jJELU
mEqMMnmh/JJkcgo63v2LFHxiTU1+pbCY4fRHoRl06jsFhFpTkWOhQjvi6Vtjr1gyZ3Ea8RI3Unqj
mP39cDrU31vY+cq/36vEqxlnts9BvtKzr/h6HrOshLHzW8wk7Tsdn0N1XGsq7Y68JZGd4r/KmUpJ
4n8pkG1rJTlld8FF1KqJbNvCYQl7mFO6cjn6j7L0oFl0OUhPjWOfd5GNtGlO39ibIYpZCbVVNuxD
JvvuE+xeCucGT4si9Dho1LlPcW9Osv6Ogybve3YCGknOitvp1xv+JwEHbuwJdV6b05aLdIaj2+Rh
LT5SW/GFwJVo8nupG4kN9ac6VGWS43mrq+Z21/F7bpOg3zTYW8pjBuxDw/4x4FxjxOuUGK7M73yh
QmVhRBBbPN7giqFjM3+J8hF+9R/LyZfSJ5mdC4d12/vQAkQ7A+SYPFRv0+m7pxdeDDMzmCOvRyLW
WArpokj7l0NMhx97gNHnt495Ijk0sNe62IBjuRFjwQHAGuHsf5gYXtcundVoCZFxFtJf6M5rVHjA
m22TkpsDkt9ri+5GYNoBWH8Ijf53m5lPTT8Iw2LhgQkDA8FE8YxdsHIrSJrkr3x1C/+OaWUOuSkL
t4Wj84tgDgNAl//LHjfxcWw0AD57ak6LACxqvZzqM6Nl+LDCiSH8DneRWtzqUaAvqxeJvdbkeXqa
APe7mr+xeEIcCatsolLsl09HowbZVmpxm/a4V/1Gl238cPB/0/IwF38Z7VX88xypqFgmOYVCfo/L
X1EQX135Ssj0qYr21dAXKwsbfq9k/nPPtcA0OmprtHrS3+weIJfllEt3wn4S3AUeGoU3nW/xLxow
lYe0aNgrWP+r4ER1XuZFsMWAiioumSVXFJl2VodwzLLTz4JZ35u9xZjGWZskDVa0CCKx56WcUp3P
euYCxnJHWXpQh0cxvbleHwxYucWalACHYM5kau811S3Z/j7bSpbpxTKUV49mCqQ8SrikvWpYS3gy
uOLFPKSc6E5/xAB856OAHCOCi0TOWPDUTNvWEf3vanPb9oO0jCyoap+h5v/8C+wTa6rSqxVYaTOQ
05pIC7p4zoOUDiUFrtQBt1rpZsEbp/P1MfEl57C2TUAAYSnTbBGsg/5Y43TR5huY0rmN4c0on1ip
IDRyPwRNUWFdsnZljmNXwxMuDnz++VG35GUdDEeCL5n/+OAvZwfIyMaulwFHX6vsk0pTJNEKmgMH
SQsvfhQfF3DNEKHLih/6DiAnOuF1ipf5UeTxCN8em0WFba0zJaTB8SuDhOM7jB7KL/ZtlUOCuISn
b7hj70F4MlajH+0s4fbYSn0PxSyvBRB4m2w/bB56BmFKnUTTAjdJl11RDuC5/Iq2etr++iNC1kR1
y4MS8wtKSEL0I5lN9x5hhnBrDuZzXw2jEPcrU56meCnPxs5p81PpssrBLbaQjDmyaqG+wI8209XH
hHagxLiiaH+gcSLG+NzMYW91D2MRSIkknguNPv9IbrQdrKVtqfZuMwKdV9g/mqE07AL3TQLmqpdB
jdS7MnBJRZ6k5GwVHIuK6mC6yZ9D3fPv8UcGU2Ztc+UfyqHQnmrCNMyUpIz29k+pBTpQUUkbRwzk
yUNwOPJ/bpwAWgM3ujdQ/jvp+98zaFNugnNNbkJOc4rAG9xAWrXUHIapV71j3kW1/fVSIjzSBEn0
+tWB/Eif1o0zLNHxsRYWTvnYdQVPQMueRPevFrI88g3EMbiIab2Bn+OYqvWaBUTg3PbwmBbVIQBG
nRGoEE0hFpjqxem5VQxkVzR8WUg/uDBmuUo2t142Tl6pZVXe3LCHXh19zZ5IuSk53QoC7J5WsNV9
r+kGttaiIVLpfh4U0TSp0kfHqwYeaXr6Xkh1JtHDErGccZQGMjJf0+c8EGFEbH8tNBQjPt8WHehA
EZppw3kaN9aiJO9ahenxYJrNt6w9ilyi+YubY+trek1kJNvFLc2Oz3nBxYdzR99nSUHbz55OcgZY
+SNsVvo8ME58uI/VWG1kaAQLkD/vpXVqHE+3gPKZ8+xFuyA2QuJrv0fkwqXlXhhFq/zytkJSGrQF
r45xpH2R+mpv1sh+bUNVj9qDpM+9Sr8XYkPX4pAm/k7HOftO3wwvvX1/bdYe66c6t7U6dgCWrW7Y
2dJNTkIhJUFiJ0YuMsvVke0fpHu5ja6UOz5mt44lla+aOmOovayYqzlI1uxiJ2Z8qmPCyFdJrEk/
t5JYpOkzsm3+jKZvKH5kPWIVeFC7GHTV1m3f7eyJ1u1NC9j0lKL7TzDcYfweq9ZR14iWEkBsykwk
OloaFV07psNBjG98jMFGQBRVIQSR9/aNWu1BkI4JARkwe7963J+t71oLfWqdfjAGbn5srMK8oWtY
tGT/y9taB1mGy5G2FAIPgWpPTnGHqHKz5mOoft95ajBk16K8mcD2QU3micO/8EoKFcncDzdhgEg7
ZFcxVDb+Uz1mUQomY5Ic1Q02WXFGPqCYzCIKN49MOxctTmAxp0FX08+1ENFFwDCsqA80llkaoJDp
V7jZo1JCVhZud0FnU27IFWIOpRWZu77VAOrXbGj4LrZFJgXaghdonU/3kkoIZLKHznCAbkpc35dK
PzbiEx6b3w+iLj4xj24aocA7sS5pzNp99bTo3nyEW5yAlSrSJtU7QdGIQawtb7hWHtWNZXofuMDT
rPePLzs8xO1rgNMEKEyolvjm046qGMuPlYVop5L7u1erdXJUqZhLeES5OqxHf/mwnyl9okUowQVL
DElBpSXWlghPNS2pNL7BL8/3YH6PfyWAbmZSjsisNGJxw7UOEWjWNCskWJGHGIVTIj2hztHgi7oz
fFUJO8NR2OfwIq5bB35OseQ9GoK4BNiNyTBesCsar7+hOb0rp5PBvrxNS8BYfKVJ5JgQHrm3vg2Z
yPxlIUTi7u+CvKFNoggPEvuKxPHdaF42l7vmv8ySDT5KnHx3azkFdvTZnoRS6zHOpjXcibLr0H1t
cbUj93F2jp6Mu7eg/pR8gQoclQ97sHYRr7Es4HBURfsWvhgUtt+Tc/84OglBW2Lx1gYtg/89WFz4
03/YFi7VcKgIFoUkEG9dGVY0qR7lehD9H1ffOfMp4iM9fQe6JBNMQdIcoIMvts9sizQybUyyvPfz
1/7PC06mzAhcUxhtxvzlXt2RoA2bVJyHFV8eLQtMN0BLBqgE2Ru4TbZzHhWMSPsV64LxJj0hrAjo
rg5RqzrI7xO4XrO8WBjQL0Pbkw2Jv1GSsYT8GBqpwLoIzxpp7Ig+V7kCwmkG5CsGX6S2Cm9Bs6B0
+rEp7Wc0aOJLLqq943bic4d4Am0JnOJkXNBP6kadrvZZ+lrXMwfPOQiQ4vYHzEUcD0TBgG7DbBEy
Eeml5uMKnW8MIbaRWlERCHZEdaW0Rh1RU7HuyDA8q8NwC2MSTYwmIzAqNzNYodCkw0lprT0q1nQQ
gbekMhPiDlubVPFSUMG+nltO1Epfla8bXtZscfqpR/I3oUsHvcg01MJ/feH6uOpskzr71mOyj68F
2TYcWA4oZZFCU/zkKJmYFTDmgUrAGHNVdik7RoKzgX+TRfUR3XuLUST7hCGoejATRGqzuQbgvaaQ
/wtJmTx/q1lX+cFdPjwMTR3zlZS2LtYKNIUlRJY4bY2VwxNH95Q5khw1sr57SfF3Nj3G/pxipfVi
R7BjirO+FHLgMG8+Z0LOfLXYcSGU94PmXVKyszvaRc8AOiD9MNUCI01mqZXUlv/PfoVpJXkLVYjd
Cymni4Qv1IEa8NAIxhwdwZr6TMy0NUO1Lu43nPr/HJuhD0ityrian3G1X5aOwF+H79ymbR42u+uN
38aA+w3aX+6py3HabkN75qcgtPpmCbOfw1y4XoxbiUGOcbkoO1vi/8eFxphsf+Re16MGyK2s5hXH
vhoAERkgrgxxn3Pz8DoTXJi1YWm7kaQzYWY9bSvxTUIi6Mvk/uyvxkTrLCPUpGhLrPtJdGSTsZqV
jSBOlOTahCnzH0DN6MFgmmbggnVs3vpLNEAjgPAzqtnMdKbiyrjr3CYRKn4M97BW7SQLL9qqH5+0
62pGbuaWXVdpXAMn4RVP/O5jowCXxEIJ6q2EWJLPn2OaQQ4hrUAUYSdZQqSqR7Os4e8kQGuV9A2J
qqbV11BfaNbIww/QXnrOl6rHnTU9itA2kQckkVmRBTeutfvUvD7V+dX4kwtiC2+/URDB3vC1F2Qu
N38oazcBSiGx1AwKhPIGSjbJdsvWH+CpaOYnzrV2NpF5Nhx3q5Z+8WvN1jEvPtzwTsddkVQHPdtx
ucUacsUqk+d9ST26D5GUEnUEbjf9RvdNu/ORkfFr5YcexObxoox9pr+CWw94e4tS8JakSKY1R2lq
Pb2W3X5mRfa2hXmYYhr6fiNCsX37tm206yes8q8QQuCZWR7l3dr6DPxGJD98UzlyREVFa26Vib/n
WMJ//72tnMK54cv3WLpepm+PvMre+yghkoCQlMo/trKpDOurNE/Nt+FR+YZAGhnW2jrl2y/ufT3X
hDRG+YZvoDboatrAfgOPd9NLbrXjrwDyCc0q+pMBj8JWH62oh5gK41mnsKuAPNmPCtll/15U0u/+
lknab3k0PXW1pLixfJqGHaxKToV3PzrbasYnym+xZ7gyniAqb+6v6U46+cxKA9MOn2m+2/tAAyTn
ZNfcEk/Nu5ax3xjIvIEwMThIKeYTUL7diOUKpetNofMbW6VtjOKM5+61KppBpk91SZfX6kyk7EUM
lI+T3h1YiFl32jZpWDXMZxapSQReltZu591ceM6rAFL5ThY/CnWwDpwWWkb65wpB8E/Zm6x9W5mS
rwDtTg2HSQn7MhIC67snX3cvzNDKveewcpzTjsIBBlVbC3xFffoUVoNKyidHD39l+wO2JWv1//ic
jxPbKVKIkjSem5ck79hrDYjdSIfY6HHWR8w6NUi7J+wXUHfQqhfD8CRTkGEl5LwKDzAnKLbzKMXf
mMFy3O67LJt83YeT9yWOxYMrukYbdkmwvPzywnKxSMv5R2vkvrFlWXWzgB3wlX3dB1DpMhW2Bi5h
V/EUsTirZmQ1QG2GsQv23SZVIhOn+L44eHP65qwZ6tfSOqkww2Q3wnKoXWuBSMJAUVOrAQp/qtdX
h1u8D5DA0XTYJIsOMoN61K8F3BQXi2P8epRykHrMT0aZrMWh2jiKhPD6JIXzeG1RFw7VcPJ2WUjf
M33axbdMZRDddkVCQU2rr0TNi9V8t0VjXumvaz3PgJbxTEi1JAlwuWMqjn7zF7QV1MH5Xhk5g/59
KIZ5dp5T4o4OINAc/V1z1fcfEGjMVWPlmiRMXmvo/t+W8RwT2CPxBdKGSekEgrdkwPhwbRkN7n3+
3y7c2YOCDtSxNq38scHEz5LFINccbSnIJA6xo4UsOIA3Zsgn86vPNkiTgE+Xke/nCzBWT04UsI3l
Ks9wZCJZD6tspOae0Ez4+d42OFfRa+2B3jdJG3ZrPniNmdziYeVu6cnwHXlr33MFRDmBaopwTP8W
whliamIVopwH4JNdNu86GZxmUGZxit14phtCs4MtJQPy7FLAvv9vKxIYvp19aGD9C3OjW2C7TdH+
QGGtIyFVlXcsW3dUFz3XinetX29GpyXddPwm0EEpPL5zFxl5GflRHzPA79uJyNywCByErFJig535
NUuyj4zP3Pke3lotsVcBSEVk/FK5P68D0OS7OTlEvsVQ4x9i0RGwMnZVQg+SnHEuUECyAz74Rqbi
9k9wv9kAkABE++sAknvA/3wGXjOn4CZyZiqBdUMtQN8lF9VsCjPeGtrDehVjzKzBu18FQcUqwN6Q
DVNCWqEIyh7QX784F93EXfdGoKeGPKBXud9O6vHNntUczzfli/fpbL4RZAg+LEImt5FryDHDUrCz
EmoiUK/LYhYXawT0eCxTGiOuDKoaJpgs6WoOvdCMG9zLtxzo/81GGaOOQUQMrlaO26gfAYIx9aTC
u2eBBXAsh9M5fSeCQggTMpOO43bwJ+vOPKbV0ypPptVUzXZjjbKEhxfu2st33Jud1/9mW+pL5xUG
n50fvFcRG370+FB3OUkgcZ55d4Ouw/JpI/xoNMz+VGP45jSvQWOxZyjRBLPRbiiJY10XXMGegoyu
tLpHNLQx4QjEEG5in25V+CokO/SuPk5Ig1HRJiKV25lhuug/+yS1pe5KBBLpVVz01jaJWWuKYosO
PnPgIeBI4/JInUGhcBxSHFMGWKzcGSpygS/jF/fjDLpOzttCpzxCLgUqrT9kG3Ja0FFw8LP8YRY6
WHvw0ElcACbe8rIQl6PyF+d7qKMsvwN20iR2w1Gg4gH13ZVGfq1d7XqoH1NE02SNxkE5r6HrDj22
ZbYhflzu/AT3fX4iTM+gVRID41omBZnzCvKuzuv/V1hAY4hkegsfkwwh0TeAFaYNF8T/W++Rf3kX
wFodn6HgRvBZ/Qk5FycSyuMWh0woUxuhYGP46fMJMbwf7ZEl9pWxsoHdbrJ/bsdqJy7kEp7k1thK
qiVWUW1F198gB7J9YJWkm/FcZjt8G5KLbstVBrBStxHYtdreFlgxZwV+UmQreeUFKXSo3pc/XM5r
1TvZl0nB+FUb6k7F6z1b+HH/NB8LfsqUH0QZbmXJn2WO+YoY+/2WFNPIPvaPXM02yR1a2zz3bFRi
dlti4PetbZBE5c0s9c6sMRxzKMx1sebQstR4S1FZXzavUXsxceMLSoYaETqJd/rDySGEwqV3aCvv
4lO3Mf51Eow/ewtqxwM5iAx8e3EuX/3AJmlyyNAoVvQeKwvjP4c5/ANB/YdGr3Bn/JE4VcBcKpv0
G/BpI5F+JF5BbiDoUpSeTfXKEkoEIP3RTU30+D7TpVI7SOwCQKlxJY9oA9YqjqcCpdM7oFn740+R
Lwtj6tEHey+2wjCsm9M9NSnsq6rtXB/HPwPOPMmIt/lI0PDwqYA8vRxKvSsm7GLi+8RCJUR8ZIZ4
YZdi8FL6LNP0aoK6pvl7FPov+20rlHtVmcBRpR2vVQIDfupewxrg92QPhfkEPMGddzq05KPP/Ao3
3ov5KPQAdi6uhdHhWBbp68dZlOwJnH8dVnycty6cntfzQ07/yT2UXgb9rCsDQIVvhU/VsVNVukIz
g6L6gJLMqZn8xzCV80vqSojuXooF7fyslEc+KaMytbKSKQx/Wk7HbaN0HhfbX4szowzAszY/IH6B
9ujp3nWoeYk0jxfo7/pqUY85qRnU/2J8nME3Zxe0rkv8xgkzd2q8SspBVyJKqVObncD4wTFrcNn8
FGxjKo5vJup3D7LeBxwmoBswFDZ/Me35I2X6438WRFkAY3oD1GQN8KtHPh1MdBm5C+kG1yLdoCm1
UHn05+EuIbqd3Q84XJmLo+mkN0Ua0npqqqc2ldakS5ZkQLx2aTM8A+lR0mUpzr+BUXFjiIiliMKa
ZZXqMhuDaoaakOsfJ7mUTot9a0iH8hN1uDcj5wn2Np+IT4o/Cf0owyDe8KgIGuJRULaSpFqVMz/1
tm9vSLbTDAhsKPCO8aZ2qrHqrQlH2mlTsKC06e14G5S+4/y5Bv1ywjjOEgvS94rZKZZM0U6PYUBi
9Q47jpU42J55gaXRVNghbyGUatwx3bWdozDz6MZNPyNMIbi5uydxPfyVnNYzWpAmn9JNlVA8THo0
fb3uLFci9j0JMJWwr2S5RYj5j1Ix6dK34BleV3G+GgDikBIAh0m4U2Esk16TD6Eep/TqmThAV/uD
rH+F4EcDoAFDNL7kj/DTm5pgDZ4TkmfcB/yxflLG6Jc+SY5UTYP+bi4h2nJxr6QcgyYEnCRD326w
7JUyibi92MNy85Bl8VJtP3XQP1Qj+6a0nGOuphaRIVRCsY3aq64ZdlUcK6lVjgYgLd0/tPmwq6IC
kiTvjid4OdrlpIaJEqh1KH4teFVlen/ayn2P10qugY/zIzMTnMxuSuBRRHFfdBx1ZQK0je+zBgMD
ahOPLRjTF/xrK2UmiWZ1CbBvCk7juB7swxb4+YPyGujXuBlfaylmyU6tXE2ebetKvK8/vi77C9HL
DyJHwBr7Nqr1dOdnTsYRdyWkx8KhjCAgadNUKyJmVNooFLIAtjsN6L8yd574DUXyfqMHzNshzF4/
wsRmuyAUZ02pfqQ+Cnz2ICOBWm67zx8eK+UmtDsSI2uwc2YqMaH+ybO8E+sX+z9WKKef+PYbUh3x
4UeR8JOY5myaHNRl4PaurKJleUe6vUmA3RYbj8bbdC4kkKdHpAdV5Lv1QGn1ZAYTjtSX8jPckDI3
Gxxj3iJelGZOQbkMpH8650M60BMNobtpHlNLppQ7e4Cd9czfUTfSQf3YLxlLmsJ5/WqANTLn+TKN
DrJpYMzqhzHV+c5pn+AKhVakGO9pWxHmK11O6FKkT+/CKipquYEYmjKV8bH6TkqCQ7dA1AFN2YH8
RT5xn0WDGRztEgDXpUGEY9pfpCynGlbn2jq+zGYq47fKmtaQWv+kXC79ntyRvw2kkbt/+MUfCFGg
06oScLu1uclwulpMRqIoKbedWfbwV6r1Y4a2cIwc833a7aLVlNfkmCW6jkN6PrZdZQTO3rFf0Exa
MvPEv2j6+reIaWinxkZndKiiUk3G5XDYsV3TOUvGWNfAMDL4gAwZyfOIB4cIiSYITS6vIWLgpoUb
kk1zBTCyzh6JZQRxLdngNQFgzfAoy9L9m5g0+Sjmx0f7jzUHckPKKpBKe16iK6ZSnqWw3rU6emB3
JIHDZkl6cLsE9y5auCkZv1tjqGFFdN++5ZheQHaQdaVd6KYQlE6FJlbBdnUCnndRg4XBIIDUTmNW
1gLvYtTgcAi+1pqxptZo4zngaNWhG4GlAu6JhmA3W+jI2VwYgllHDS+gwlgcXZUtUwwRSjjynHOs
PcNfu/kuW8VSPmClz0oi/BiAGG4Ul8kllvODvFtQJylTeixVrck5CDKFRzakUep2jFpYCsEL+McQ
9WTbtl3BFehou1XBe+8nm01MBfVOCx27e6bQhi2RT7T4T8R8Hk4Tl1svReSyIiW8GyKG22RbE7p3
o8jYFX4EdtvuWdY9SrT2nt7P7Z+eX57QImdKAz5/95cqpeMLsH0samBro5BuRqSWN+3AA4ebwgfZ
5qdD8/32AqlNmxM1Nrmx+Ohld/sDS1Sl4iUeW6urYdwV/CYvWvAG8cwhFU4b72ozbu96JQ7f0jee
IlXn+jj6qCzGfrkmviBRpL5ES0bwhznaBhJA5cY/EW3PHP1kB01h4CRrhMlc80kIXaqcLRBfmdWk
babZT3fmdxTEuPGbahfcgixH0yBrdlrROGDAaBQvDMa8DwSTIWaJJ6tzf7v7xkVkS3PezC+ZXpRl
/nm9F4Wfh2er7DKrSJvv5RdYRtz2QY3apxd0GthFGLK+KpsFbMdauNqsc4C6zBj3EIT8O+S4hAVi
4wNB+fZwCVhDJlswiFAROnhmLZDyU8ETJ/h2atOGIj/R1yvXnArn+X8BX732uwTs4UY2gE5f0jVM
tFSLYad8sbsvgkpT1sMcMDjeY2u5i6KV2LnaRM8KFm8GrVtnN4447XZY2TUA8K31RccyJzPYGILb
jpXFUhlvxGr/4PYUMjrixH2K3y6jvmQ1VgxuqgPu+04dMf7T8lvrjbMcQpjVNFAK21KhZWjMs7Wm
8JhSHtZYbjn2owRznOi4lj0N+gCzn7ZQWSHPtVRJojhbqhKIbaJF4TeESy0/KNFe5zdt9QReMHGi
aO6JokpWNNQvWES6vdA50Kfg0DoeuadsoBX2zVIthvXjMjmPy1pjBihWqJrGwlMPZAgy1wgx9wlC
Qblw1d89H0kHJ1N//s/9fr6lpO+KmRtJdId69spV1cssfyWB19waSd0EcaITuPZsOxVIAodLeD6y
qXin3po0YpVUELHLEieJvGotdE8QwfkbrrYMRBZG3mq86VYIxeVS+nuOOgzR++Fm6OTmbhpK0rRG
sNXJUf2xX8/WHj5nJez/GiglgGYTKVGc/sLc+HlTYyTmvMSiYHUckmBsUn4sOEUR6BaVjM3gAZ0R
STU13+fVi+mnIJNVNVfmej5wBEQeR5AJ8fIyWPlKHnJ73KiI4DJzeOH2CXIi/GQsElYIPSlY4u55
hLHsOi42nzUTyDtAeS4uW7N3OnLa8sAKdzTFwSgJIAtGjPbdv0FX2X6lWJkNHzC0DJM+njtxEmu6
EnlI0iE/iBD68mw+miu8iWBvUEyk3QJUjBR50agdLTDi0HVAy6+AJaiPgoi+GS++wbgnf0DQWEs8
nHdxmoOs2sA12P7fJNllkawR/u/8OP9/68us+K8mtzHU1MgtKK9rhcNZcHdHevK+lhbPzqPtiBLS
7j25v5nKfUKna+P1s5uf3WjwPmv0ZQHYRZ9VGraHItAevY5lx5vgYPMfdo1XPqoniS4X+gKWp054
0AzDo4sRxb53tx3fQ/dpLUnS2Lp4hyG/XOTUTE4LVvu1JIoTTBGeiLn7TKGZFQ2yT8QcZ2gq7azi
antcjWpl/idrwh5VP2zjFN/uPE+Z/qYIxVt04bpwq/FgjPDhT/x/ch657OpirkWoKvTdH5MVmu9F
d01OqvOPVbXh/d1JmEBDeQiNQNmeyPkNP9LV7MjYG+8jO+FL7r7QmbM99OHkJ7aPuVOke434YXhH
joD4VTIMv8vUZh4sOP2vA/zWZW6uYRhiVLmP09ipqagwBWVpEr4hzA5cmqcZfcRohb5jEvAiVOLd
d6mh/3n/OP4Ktb1AB/VE5O4VkqSFtNh8u2ZfuR20VwHgO5nxXAz20IkoQliL9fLWtm/CLgljyBDf
J0IPpUpL1sIfh1haSeKsAtnj4kEgN9sTBF93FuI00DQjSQpLTTCLS2Rgur/ZKgXqcVL0GETfDsnm
8LKTMqpbwJf2fA7WJqaSJBFx0L+2wA4MBc/kDwcAvBiO+jDDGY2Hd3awNpBd0iXkDMd+W1QtOdRM
yt8BA6Zu/x6w+EwISPOTN3TL+1ZprVqX2Y5gCfQcmNZsgIIbaF2ATyCpokIcGQph9aFGJAaa8yPz
Wb+I3yl3y9u+onOvcYE1C9XuyZ6m94Kkxo2vmjfhbG9kvMhGvwLyv0C/q1u/r8NOIHIOcx+YBwIW
OBVOpp9RxN/2FdjS6d+dAnKIIR3Ew5nF5GcvY4X1Visv/bImozmBWUQkHFQ7+7eyQmreZmUWUf8r
aGHUOaMrvP4LHUQlzEACoV8mq6K9nOG3nL9oEuJ2gwiLk44qmb15a0qCE2I5tqAHPOVfSCQ0yfpL
D0iTWStApICgkoSYYxrV5Pnvp5WZrs0QmTPzYg82VDTHS2XNMZ0Ng15X44WEtLCSvAHhFqCqokYI
CXqyGsUJGcyeQNitxJxXIS3w85fBEK2v/K2YRsfWzNtoHwX8DRduggKbFdNGgW5dAQaQyNZI1U0S
cWHf18B8CCkSrkmV7350gP8zDOxB2F2UKBVD+xv6ObKVwl/855RDFS4FJGge7Sz7fF+aP48vf7Vn
zqyJcrZH7wlTHLPTbJP5QuJKvgLmMzC9EFrw/yTy0fWWLuqHGz5mTX9qMcDxLNEa5PK99DFyZJmu
yg/JZWEV8+B4agYwqP9qesA6eahyIFt5PeLfGJEMSFwdPfe+4IznBw0WtLWjtR5Dv7nVJRHT9qCl
/HpcAB2WE42BFUQLfuK0KO0W72vcs3CEbcZMmSxKXonQIKlzAzXQgeVaUSz99vh1th+1wR2a6lxP
kBnl04WlZlYMS+icHSx9/uirEfTZM8Kl2VMniRMLDCLiY420zN3+EZLtERE9WqZ07mNHD0tyKVJf
8nQBy2xfUMPvzfd+MUG4cwv0jVeEHH7IH2e5jF/orU4kAk7nVOvJnvLqIjGqn1ttgqS6OiYVUxVc
b/cVzvpNw0m7jpJjkQR6XXrZu1eLb88+0MCv5foPtjyYA+WCetTmBfHtykgqt7rX0dHk37/GSgMe
Wf5Eo2ZO7eaGyQppOLhZFoLEhUnsQNVxji/d6jSUaEii/ZDpsQf3ycaNTBgOAaD1cXHfA7RX7NKA
Yuccz2JnYVLnZP210xwPhI3w6lmGdOjPUQ4de368NEWPowEXnNejTBSM8hrs3GcjYo8OomdJPuuV
Hdkbyw/DG+CC0BvSovVzQG95+1nJ04E7qD0rRfpHDTL469aekcLecnKqLMhOr1t902Ve7+J+pMrX
Q1LxZRgwinpcICqXi8tLi71qOfkn45YeuDId0a2FbDNez1sQ8+ViznmZgsoIJ+bTdguUaOj8hSka
gaKaKfvchWZr2nnf3PYycEsk8VRFHHOEjDkISxRAmOtBVcVP57QqC0VmuOmCnZ+EeQuGr7/RK5gJ
udEg8QNKexGhzcCK8EwvlreZiD/xNJ0Lc7xdVrXbiPId4B7+SWaY11a75I+R6n66B2P1DInGwoHl
YMjLgXsm6Z/fN+0dDQiBkWFH60GBJSdysdu50Js1m6jmSby/2jjoeH55eZ6/viTwtkkfn3cmIKMh
LKE2HUN+gL0vdcfVucp7dFIuGw9g39a2tgqT+xSa86UxrALcTVZxNl1f8xCzk39H2MlsOn16+QYY
NlMOwp+1lHfnQ8D6rGWx3Rn+mo6lwC3j5mHZoej253SdfWPDhkdyPi6mz8jNuWLKdBjMrVey2LLZ
ShU2lbpQhuTm5WmEuEaOfNa7FJi9T0HnXM+ERAUwEwz6H0s5F0VobFq0ZEJbEonUvNKIChnmFQ2E
kt6iHu458ip574bMaQ3RBBEtPzKvGtFKvRN+JX+I0M0ENqVFjhPJq+sjZy9s+zc60E2HW7Jqk5wt
u6jgOankcOS9e3KHYhYydEmkxcPhXp5il9ql+MNvF+5SBzgAkEhKcG+/2EoYqLzs14HXPBDr+NsX
g7UZAQoazlT57m2LjpewRzTrHdvM0lVSEyyzcXYaOnejSBtq8+DGmgwAwhH+W7P4dE+AwtYQoOnI
8YSHhHWOTVhqZwLvy78AhFgippd9LlD7Ox1hKmb/f+q3zAHF+XOM+Qvk//r4T4VHAYk1JByF0P8U
RahkZrlQQeyO8pMM/hklfp1tmxYy36JGX+NfUJxCceX3ccWe/TL1Foy1Dge4upA3A+tmQmrtK26F
a8eOQaAP9e0wEkSirLsoz8ghGbywTaNmvrRJYsCdXtP/+N1u7i9Zd91Kui71s+/DBTN0dtJ27mue
p+YeuRtU4dVddjAq1NPiLgWr6hZHRrQpYK21F1zm3/XKlQW4EtL+D0xV2JL2JjIP1df62FJVk3dE
qNP8eL2/jdjsMLF42lRPiKPDwaxl0yHAh8IdDe+ZClZFvYmmGfTppLabSptEJEwhqewO/DyJRLyg
w/B3eSeYUvbMUAI+bXAqRVinRfuACZ0PInZTz9YTBZM1FYmpcLxoyjlGAPxniXKrmM0XhecJNXJz
IrbTwokD942pvNGka1HDqs/1IKxHRabfoFUr1c5zqd55SkyPVdsY9SpNKoDAbaAUtuCyBMz13/t5
BbpAKLfKxmUHgpUvPMKVxn6q6SglfPaEf73ujZ6kV9S0Yr/brYmlMYPuOOkgh6SZDiwXtXeg2Qw5
C68hKLdoG5cxxfzu9NOvWSomTswHYXp2u2Z6qeae1VMnB6x/GSJQ38pgRmaZgXnd9SAkhY0OaVVI
QHmNZFYtjeJVLGffr48IZc1EWEwqu5fn049VNI0i2OfdOnyddRqXBOBzkurHc63o4RTYsUu8cNAX
QWzWTdFhSiU4kZM/bRLc7C74g4l0PdXNx8CCHJ3wH6EnVhcukHePJKgaE9LvpYNvMAl4VqtxyVot
/f1Yoht5dgyadAkjEFAXl5TTGDFEvftxRgHKfViLaSpiEgLQ0xsod1YJA+Z3JLhAnZOC0fDcUJjs
LvB3lvz49FlxZ9d7ReglAedDfm7oVZhcnUXSAnAKX1t5eGJu3G8qmaFLrhbD67Djh43u4+3JuFcA
nZTLeSnjepyndG0hDJonE8FpPpotQhvngcUmhAemgfd4XALF0v1r8NnzHDJu/D4OrYIYke91WHLp
cg8bwJKnk3Gs3UEony4dRbEvEq9RJ35tcqndcHXXXnSB5xRWSJgIgU0klloQFkV1UOhh4LZ+m0H6
TFF8f6DeBhDVkC9tQIQ/sWlXeTjUEAOw9DxfA/fpmSufbm0U3bOx4qb+LmEJtAIpXmcmbFCQRRk+
XNh3AGVK4MPrJLB7qSpswo/F4A8rc8h4CZb9PU6tBLd1BtnE7Sbflt9nh3nmFdPJHnV/DVr021w3
4FcxtulEjRfF+NHUe+he3lHyx8fYDbalveMqjOHsZJEhfCqZKxCgTGPt+xUmqmjg4pveRlo+FOZV
BjfZXl+r2PK7YL2jNQYq9oJyZG8QBfgx5IR4OkWnD7lINbpmuGu4pptMIt88IlSCaGvbgDH7+oL5
9zyLxWrivK48ELFbQh/aWTIV+KpdAE/Ybl8CAU0kDAYfxWYzo8AVw3FgmNLHYesFjoa4E4m1bwLw
mTgcZULpY6Zzx2OOV+iXzEKsh+6VmwT1rANX/hEwhafHGmfK+jzFJ/VoYDLM+sBIHCIwCwi9FdQy
RtHyefF7p7NabE2Wui64nvtNXCYeQVWOCJd6+3K6HMrfvok7dEkX+fUrT0ylzjJqHLIBtGAclcB8
UucJkRxhBZ5QfdDkTjmJHhaOTpoz+qlMZmRgaxfM1rxKr0fSMVB/ITykFZeDSi7hLi5lLomxf3TG
2hYb6qrgNgzdKC5ykhOrfpf+WTMP14ArzyjDRFgiXU37pRKYb5O3lcpbzIhuaq32+X/1CuyBd6Sf
9F45SgeCl5tUMF87h35ae5T0VgmHS4yt0p5Za/cVFFi8fsYs9JbSQGqqJCAKb5YrnklGsaWeUIiH
xawKhhSvoSxvxYsU1MEkQ3gNskoR28yNmHuoC+eCXMLrQteXlT6yozOzgxTY6zEbt5qO8bOI6rHN
WTkhv5e94tJG+reDFSNTU8bJKeJvUGbTXkFGERg+nA/LItVDGRdYP7wevcyhSM/GJOIwRczvtopb
zFi3Tgeqr+4ifi3GwR4gX3Ckfq9RxqHUAQNGmVnUhDCVQtIlxsmKgigeLKGEwWiJOyNDGQQo1C6B
7cjTVXk3+CbnFuqlOXRFEWm/9xuCH9UUJJZbXJohOd3grtExCeKb3sUTWnqtCJk5dkWF2HJAoyFE
QhqOBg4SAZrNhkl00F/0eGf/OuTmshyMib0Aahg1oRg3DkXni5goTl8ypsmQxL+COSB+vvm/8PWZ
/Rt5Y8FelNjC8TSXU9z0tWfX9oqHZBctXs9MGs6BhOArr4AyW9qswvOtHGuJ3L4K5N0V/r3hRgTB
RTJWAihvhXXhjXZCJzySjF0ln0kVq14pAE7OgbaLT/F+MHYKW6bAD5tVu0/R+MHemAKygMwD2flE
WpkV4qv3M1Bdo4bxS2tTUH69fmI244epXZhh55bKcm87Ji7007JBuP0vWLtLqcYi4UA5EZlm9F6F
A5U4QfN/e1vIRXn3BJb017V6IMpm/1L/CINyM8rTynVOjCpj5YFHHpr5fiXr5a4aZGiw3byQDW3X
Ktk17T99ElI3f9EF2yBnV5j4FuEy7XG/rbLzEE9SN/Iw6krbg9NjXV6zQFO98DJwyD1y1cYDLMyR
fCwtNwwzIFxEpbWNXszKrSPwzY23yH0c/MLTB8OU1TBud0fjt2s77F8ZXmrJK11SBwm0WWXyq9/z
8exoI0g8Y/o3gJzXeKQSljX4eU3Cs7mvzyu4MjxM3v5qORQllkm8RoZLR89MnGHkVdRzj7EQxXMD
ZEU5dWJgpRb2ttp++h58dOwY9iT8wPxl/AyLZeOusFBYjr+kSzoMfpVn90f0EDNv1NZcOE5NC/KZ
hsxiHxq1VH6K8aSdj/E/ZySo6WQZqVxnaF/Ho/Pw9zgol5N7O4xiISekGDSLSDw7RF9WbEKSNLcD
IkY+oj2fa5QTx2eXKJro//wUEYEG5xX0d2gMRxeA7r/Bin/FsMsU5fGIx3CyJGuSqhJw+z1JUy7J
RzPIRYPbGWhRdZ3qS+vhWqnaOS3YoVSRHxm8iFmY6xJ+KWPj/eCVuoaesdIMLO+QUmJ/10J09ELL
A19KFcMapi/oDbJ2X5lbbbleHUxVRUB1cKCuSCCgFikLcn52fMAK97QlQTEgMdfvcoh8jSBb3NVJ
EGlhmzNOHSwJgFuMSn2ZfU5+QMYMbCJ0t0vDmt+hzZkD+H13vpKCOrB85xVCzXu7rnYj8v4MuaZ0
0+piBYS9AvyCIM4BACwq6yRqWVrF8Y2oPtr/KR4Kt2OUZ0iBpkpRbo6L4KAaCEuxWZVv0pOoplfj
oAxXinvoISlTBAdj/iT9x56xQED825WDCtB+uFkZbWDYVWQzEwhosSn4HabGKtoZg2nqmB0Z+A7w
2UeuTuW78y8kvrsp3Pg+pW561nErvLSFGoky3p4UQxuhQcAGGGL1sAh3fS0CJgutnUxdZTabsxWT
h21gEQJcBM1u3JTD7Z5WdK6pzvj6CeT8HSHAvsNWhOQYpUq3a9IpfMqDNMBL82CXsbrxEM+xi89V
Gk9pijKReeg67lOU+OjjpW2UMr7hYbs2yDAJtnNUGrJxTrWJp2Bhi1R+4g1zFc0LaIa0iIpDRxLu
Q9oWwmKk57h3GhFwLsRuasnDrswnLy3ea2eGHMsA765NrwbH/HqEFiONp2K04QoCVrV+yz99oPSn
UBKTEiKx1m4OYMEcNdPlWhipl3ZAU3xs8kP44etbbE8KHgkTaEdoCRBuDAwPhKyGAE+1eFmP0xjJ
xnkwvXYRyFSoUCc977UikaGtmdMD1M04/HyZ4AZITY19sxndv3WBsGyoFvKoJcd09oDTbD8tl9g6
kvrGKGLjKccUZ+K+wdDv1BhmOT8QzO5migsIEuB8CrU5YaxraKKR/9Vsx8OiuIKpQ4Q8MXueV2Bq
RfWSGBOff+GRDoR90mGEu/CIgQqoUIs3MzG+A/rBD5G4ngbLSOxzFvUgBDsxpkL8wTLhrsfzmMYC
03bA4S/Z0L7u07I9xJuhuSmhh49LSdqQSHP5yOCmfOZSVYHqw39X9zC7TZt9dqIK52BUxhrT57td
rqoYeNpRzBeacDFZuVYQ2JPDqT+PTh8cGSYgByDkOgial5JVJyNqSD52pMTtyZ42PGdb9oL8YbWe
ryxwD92TnmgjNf2BYc+gEw3n4H3OMBeY1L0IhhR4NmNZh+Ec+QNknoGnkNsPOWTtkCTwhkpii7r0
ceAQRRnDJBu/k5ReqJb5WbRZ133Sk8PNuot2Q+ZJMrGJDw928XpIFer+t4cpwSbSnARMOXGbYao3
tpVGav/jP9+XE/9szp05Z7w0IXQ9/Fnz0PYwUuaNr8vqWYCLuHzPNRsk3akFGRp1iqb5L2F2Gbx8
ePHtqf4H4O/8i6neC/nceCAs/ekzxbrMay3bHRvWyM5oqrPiPfyA70Lcqid/IJaseXe2Inobl9mu
eg0RVuY14Hh4jsJd691rbn6MVVXRbwov7j0eqARHPY1BEKmxzEXpmP0ESWfVi58ym7OCQ9EQn777
OljdDTVrVdpxG7tWxBa/9o87u9dfkl0CT+I/mr/rKENVx/S/da0/R+5me9e6wxhY50BgmsyB8069
AOilW5mi/EBTn+X2T/VguVAWmuATOP0Ik39KtJjDrzEQUXZK2Gosgtqw+de4rrT6dz4GrIOJWN9T
0P+sDxYmqZZUO9se+c/HPGu2jjz6qRZIGYzQMlZoO3Rsn8MSxyOfGELDoasSsMqXIv6dKpf+5d8+
oDR+Y0gjUW6TDFn04a4zSnFJKqpxRHgoWczjjEoTzdzS9+lKkOfDv1YKMrtHBprDRJ0bzKLXWPkm
hmog8VLI+GIxFgUJVumXlyidzAzVGzC0Jou/uhalcWxjTHigTWtEWUPLq6oqH0UYoAkJVdPb14Jb
BI4HP5E9IQR9o2h0xLnYtQb4EJmMPdex/RaQhHXX3kEpdDESAzOcRCVqq8gbjXgu7L+LWkrrRVeX
wbmzaGAqJpLTvKSAWKmF1fZ2F929j0pi4N+HOHo0LgA3gyXQCezgPFHn8uoWucW0eOCy/DFhHJsS
ushkvTyI1SDVXXYedt/PRf4K8MFqQy1NOmo60gMGBR/+uJuEeWlwczL7gUAFDMMdmgOCli0qN6ov
z0NfheIEv9F/HOU+7gLH69zHBAYuWFo2hC/KqMwdpqLHXVhATWvzjtEMQF7JQnvpqHtR5ipd9srF
2XzPnanOvichh2duxs+5qZhvp0f/lyDbbPuX/0lshBfhSr7VRVpSA69LyKjn14gnufjOmTR3DGiW
Qvg1eC7gh2QqEHIJrhQTCxNsV3lIMG5h7h8zFyLdd6Z/j9HGZQyFqnKK9h/xHwFmhQO6vRrRa1qn
Flyrc9WLHu/gcAcRgOeGTM3eWJjo0luJ3H4EyDxN4HQNeU7/lTLk/Ix4sHUI2FcfczSMGop4InfO
dPIQwnwwbri0dL/cPKdYSRv9oDLU/Np4KKylpcMtYy29oofwOwbPL+VQQsC9It1xL8IURM3BdjE4
P2cDv2K01y3JCFhYSw1VpItdtb6CECuGn9+3MDIg1HqU1rvMjVneBnSYaQkphZLTX5pli7RBtd9d
+3YFT1R2g/FuGU6LMkFnyITS7vUp3zSZXxm+GTgnIHeHuM/T2EVKjD7EHIf+38J00J/ZLlEuT0KP
blsa0eerhbiWAItH2rp3+WFfwcOAG3u/2vI5aOKVLy07EofTGiKMYWpGiU6gQuluRrrFbhu+dc1P
FqpCQmkB+bFIP8XFhLXiEA1bAnM35depRIhAZohcT8O3TtbJfvC6NubgPase5MJem9WjROxIh9yL
bw0KZiyzwNoBiZk1XsByY69DkEvZBoSQLb/M/eSYBCHG/kB1vmXC73mjh8S6uZZv6xxB7+StFrya
59Migi8kTnMaGHMuiR95q6hCOLV54ixIkh75m8EgvtBtpnRSIXb3g1DA4+m6f3jnIypjI/K4mg+m
xUxcyCE5jcee+03HmasQLbXYExSOjHTd1qVp63Ha7qJy6o2tGsQckj7TCbOYS0PgCOFTMrZlrXv2
iG30jcNfrOLbITRD0kl0eX1KlTWolXElbTYy6dMab4t52FsZfWHFuTPM1XkNKqyzTDtTA3Eym9PU
KaxIP0RrWf1qq2nUeGtnY1EZtmdHGO1MR/m5SVOGoj5wSD3tFWz20hHa0jMj+0ZgOOUg3/otwLfP
V8b7PMYKm8h+TUDv787el0hD2KRcc356XG8dG0Zl2cIKP4cp8m6fRy6VDBlG5h6/nzEUOiDwpEJo
DO0qmUMtkSU+I8KRtDRPLmW7Ak9uu5/b9TbLYZthiDLH0daeg5K0MacrupxazpvUV3iABi0yBHkL
dOpOGDXN8d/Dzsh9dHbrW2keQEh3jffGCdxNVk0Z2CxmUsiL+tGexZkucWzQoe1xp2gQ8cs0W+XW
5Yx+qMKzZccFC9r+c7VOi+5mxa61cprrQkGwhXRC3Ro0c0WQely6jwW0f4Jp1DzDhLON+vWATcL4
GiQmrxIlbOvLFeB/GKCPTAUGxbeE6WNkUH2fJxOWvTcPuu7h6rwxb4g61CnP5obN9MMHIdpaYEZK
RmtKWeIJlJwV1NVg2mS7w53PclgpZTuvfOywEFdaY6vlCWJ89RATaJxRJqHclh6gta+E74aHz/Cf
G5ozxS54c7CfPoDGtviKepwY376z6srB/+4xK+BCjmAo/ih10uvgoBJjatef5nuyAtAB2jjFMsTp
TKsnlXEqE7VwxENUGKi3/pLkYekfaxvqb9+9LtqnbTAs45ilaP6xdw0sAKWH+oHI4tYIOviqrr+z
Hx2Rr3c3obiob4hEIL1bTMFMuhX5mawgO+QMHeRHYWZwL4jrN5ibwMqkRXN7E1aU0i1t4iXCG85a
5IlLu26pOhgZYUIWksEq2Oog63d5Ud5UDWY4v2EkSYU7vZnGqTL8QLkXdjDN15rAyZ+qf6V/WnMw
0KU+IxgAqdzzXpeU6K84rWJL3lGGJCTMjl9ndRhgvSb10WqwHbUIyOwVQSrPTTh2kZIxllcDrjMA
xOZQL7hmCvyOKL67989wKShvUs8QfikWm4PeyjOeYgXNwS+inwaVcKbo2Ar1NO38mi8RjcBYuuL2
ktnu7I/+kb26Vj1NWtHI1IGgoOAZo2Yz3qYBJS9DuByBu9s52A/34ZV8fUWeUAlK/OUluOVkFxyV
g6cPW40mYKF8/OwzcWkGMIFWsHS5FB8DfVeXK3HkQbsORdyiBc/fwuJJLIoEyjy7gq11ouZMLto+
LeZikGt6PIyu7EdPigPuT9lbJb0EPF9kg68BAaaIS+oy1+06knfnNjOyBC6WIridNL82G9fIHt1+
J8OKHQEWZxtPGnG9rEexD6V523mO4abFY5fx1h3tjaC9LRU7XOGz784fWSijIguKgdqHG+MeueBq
/8RzUJyPmZ5leazyKzDuw6zMhVR8Or3MVMKKzsepAcjIVixvA10MzLynqf/T+/n2rc+KkT+oirqI
cvLGW3ijfWOEGISJAVXl4iAlHVja308sQH1kpozXEn+n31N6u3QgqQmJV+pofLTXcC25Egjy92KN
RCIXLjBJGsNiDvupVykGfPZnHcXYBqWvgmIRTYgoPHYfkPEtkG1RUA7EE0tOl/NEpEyI9YVqFubx
CxVgaxFwIcqkT/Buh4qXlx7xlXBPHioP7KI+PU3wfoXb1CN/qd1QspUAkHMV6Fn8zhHR/5ub0RQv
1FRY5ri9s88SvM/Agi7J7tE/RoqEQ/KqW87jj+RaIRoFQU9dZ+Tc6lx7K0WKSuiRPpvIHi41YADd
yQOIGfEr2ZqoPuTyvJPRUEBD6VRGVl3RIlu5TqAuO0F2su1Aw06kc827g3uWmBjHnS56X4T3RWqb
MnvAmW9Ram5JCTGuADBZ6lrHZ80Ui7cRamm2MfI4w08FkoKhIK9cDsEovFni/CRsKvRcou735nkz
sUfS/kAeCZ/YnOrmhsEgrfjbTuE8uIutcT+rwqn/SgIuGGTtEIQOM2G7I5+F8CCt7Tf9Ix+VLG4W
TRcp+2QqByEwtxQ586dTobpfBvnVMQxJyx3iczsOHi0weJEq7XGiXQi8UjAqEhXvMo2Vw1Ftfijk
1alnitCUgOqzkxowUmrRbIBGc5gQbLHyKfg2EjoPxMpq1DWWwCbMZ1ZASK0u0Ob2bcl63/baAMMy
dZ9aU0mosPJjsVI4OUgIYZVxPVCEx5k4gLTcvq0G56qDhNn5RTHDLNbRQrM+m8qK35PNubm/x0pG
3wloeBNnIrRXj2X44dL6y06E8B4EXTTvV/xe+Ahp8ul1JBDvghVukwP/Wt5WtmGWV70sj+j5ovvP
CFkC87CKneQN9ztzWxOUj/WYCmOVc4QAK8N1iHa23h59xywChJdfr9KP1oyVQfn3okbzgRYh1FhP
Jz67M85T+7R9ykk3+FlYqFR79xkC9XMYPogotTXyt6KXMmzN86ChYy2L05OpWuZmrCR72RO/g0cg
KFWx/T/BSXmPA2gMFn9fZGDoYycylZSKIV31STEDWko5lTCEjKmQ7hPqN5ptRMtouOEOdVGafrVO
ENl2RungqYrcRUkwZbpbc/qyCMHrpZqqDLzV+t+GHkIj5ZOcm59ONOHvZMMhTuDKP/zoWoZtQ4XF
wIBe2JbZSbrgpVMKxOv6aStkFHK/uMLGejgNxC2u3kLl0uzvEs3X9IkYPvZyTWLvmYelD3/OzQ71
DdWlAtineiK0CRdL9DIud7ejHHmTJE9pWX/PtNBTQeEhYrepj2GQOa2hx7S1shyN4zjwIuNsW9ON
PXntM38Mv73MMEHHoSpg+sfpx9CBDo4tOY+42bupKUFGUHS3SqpqjlOVzjfPeOrGkP/fg+HCAx3O
RYQ65xSR7E5+2PMqc9F3KMda/f5cvn7tvu9+lVPovti5HJtUUkXw/dDSDUFIXdc+3huFhGVK/t3I
bC/bkEk53buhr4zhBSW1cEYoM7qd039JQSjTDx6K95+iAXr4yzxmUiArQu2KVhPRxvSYAwtgY2m8
LrDspSotNfDEk/yK2pK0vqdilBZvUAMdnoAiEs9aAGxU2fQfb6fWSOY3mn4wcO0DtxdksONY10FQ
zXb0J9tfNWaO0bKtYk8vpZE5ykmU0TeRffgaFoEiruFlymCyu69JaQCGZoqKhPOmOACD6l5r5G1w
gcJSPrxF3Q9juWTuOSGHPaTMzqlJ7OiFDs+YNnt+Y8d+2TE+pjgDJ92SKh1pHELT9wjmmaoT0/8k
D/VplblUrJAwt/2d5QY73xA3ofIBR+NvuF9lA8tZ9TKXJbZEXmyQzB3iDvUMBS6PQ6cpKUonviCp
NzBlk2Ckxe9KP9JMBiPQqNzA05Ecgm+4tEj4ukgDgyzwEFGAn2wpKiM+IgVLizMPZ1VTNkIrVFdc
GP8R/xeLP+tR0dq/esTkOJ17LfvVvE7Q7QaVgxO33i799xAO67kE++8prcFYBwzXxSCGXFMiSf83
Lbg5X6rEwK8id0M3p122WZQPnhWcUAw3hOCRrGCJzGiX5DJRPGK6/d9tfMq86BNURIUvmv6ixz2Z
uuyu1N068Nkg8fQsfR58kdaeO4YJn45KHs5Vd3bAd9L0Yu/gjz/8tbLC21YyAAbS36veo8GHKFYv
OgBC0nMe8LrwNQm39dwwb8QnoDQxKJPH7qRgdRhvIqMMCapS2U5HYK3aEMMIO5uQ1WeJSKjuvAqk
4lWAfBixLnnEQ1tsJQVnsW03Pvnb4mp9q2BdQ7QFUw5QS6UxaaEz9FUr/h6/CH/65sul6qwYHGrk
2wAcdyf2YCipjXspingowvMKmLLt/r/BbQJC0D3BwvZX3TagEIAPN+whwm86uYfwCSRqgCLD6GlY
0zbFDiYltQ/vmkwaOJiId2s/F/klfI+mUAQSJYftgajA0ri57Pku6wb/84I1Mt2VeWBlURTTuTZQ
XLsPFrpIjJV3024Ha1QvzWTmCeopngG8X01esDLrEkkxrjqLlNh7RWuONbgpsgFc+oDgNVxMdrVa
EnvVO5WGAlMLJw3F25hPc1Og7+9/3cP+B86yDwEREuOfjDYgtoGRGChLjcj8RtalXrZre4jKYHqx
PS0T69bY5Rs8ahwA83N/kTcyz10B47mlxCeip3VnfLWWCANq3DHyLLb/n4wmcn4p+Lj/FNJlxd5W
tDhoq9y7IsJGOgolE0LkDKyKW+323oyJWAAez+EIhIC8XuUu8cxvmgwtpg4TmKRjiSclW3rvVcPt
GrrolhbTM6OtYZ9vKj+Gnwaf73h4IN+jzBMciiK1DKe5kTlv82ulMLkfcFdHwbuh9gS82x0J95jf
0y2QbkX8VnjtHtiSxR9Bnfd74O0w3bfKcdIIl2jiBj7jpRxkzxumlx03XlUNEaITdQTRDshWvJLY
BZALsSsIHXeCLThfu7Xhm35tXWjeUBkM4latdqTLV6+SW2LqtSDTdP34Uh77OkH4GwmS9EtQYbzE
Dd5/EMighcXHXhEY7FTC9LDLdSvcvenSZnRwrphNQKiPW4UAZmqYzAb7X3VZ0h+aNACH0o/f/334
Vg+8IB9bHT1NbuL1zwbX7s07+OpLDZupSkizwQIv1Qic4WfAy/eRH2lI+dun2eUsc9PopuEhupMq
G/oCmuEBuwiw+nl3bd+d4pIOHBxqdZs/xmW7PSMaK28KTr/qV8q6F2RWGB3ZybRpuguXkS/0IS6/
XLWn4cWrSgmjKhi7VjENE0Sc6cmjvY2re896CeHUSjHFg6WVtiiW8cVYJ8VYR5gh0hg3jMQZzLnK
4pOD9U7MIz2WL2J/yAL5S/2TQ/s6dsshKsZ6kF+gC/Zy4NT+2qLf2iQyRwyT2LggxPrzWOwGGTeX
xtDp7/gOJQDPThRJ6ANiVUpQ6k1D5oqkJwYV1vbH4azFI/cdvg3yjbsWWltIQpfUojWWfxcwooeL
PTFtywmcAgQ6mh/2Os7FTwbAi39+uwCXS+6kKWau0KrzFtRG42IQJQkUrHnUE9KRxxwRItpakVKn
B89TACa+Jb5Sge0Z3U5tue+EvoX6B2WhALjtcXv2zylnX+Kvnj8Gxqbnlo7gHpbsLacaCqLzL2OC
/gyh389jJ42no+CpuZd7WjiEqnH65lo4WbSzcFDwhx6acJGQQhgUV7C31jtKEnmeiKsI0VEu3vNX
dmfJACuhvHLa/qtAHRlFlIkicuI6poqw71zrv9Rx5LK0iemnuF0VFN9b0YlxF/961DGDNVrM69dL
0X9BuHgiMXoopDSzWmdNwZ9dX+lsPqgjGvmylH0WpEmWZsxakS+bWk8bkb2Dajo3O9EtCDFGL9oK
VLOdyWGotl+RuYU6fmmBVDCit3gnBli4B1W10Ss1z8PXcNFJCt1z+G5V1Y0jnBNTe12/jTSHdcwZ
mwpW265vVO+/W5M9kTILlHcKRq6+nD/jVXHv9ur+uzlbPfhXJV9FhVxnmdR75WXy9g6+kL+f12VN
5riFifp/RCJ8IBrE4+fewmcx83m/5LXmcMLvjIxMZooJReGI0XBLeiKP5nrkrcRbxJ2VzJ+aQYS+
GViSEJATLuOlhkfWMYO2ynKvEeOjlX+QwH+btkxLG/RTZW4PQ7XmDz0Se1URtCGL6YbdKhr2p8b7
IuX9O6sDxRLYRjueHwoLST4elcBN3xQe+Va7NNlwsEzbR0aHABBUEb/QU4BXlv6Jl/bPp9dZnHXE
CG2kv4qIhOq6YuA+lWs3BuK49NIrZvIC3sYjkH+jGmV0AI4biRxqcB88aFMS3Kh++jIxHHUqcszn
MZ9W3PieQdQ2pUv2MpHy9Pt3/Z98UBLhFzXfcBV50V6/BiO3rrgWFYfoykepYVVo3G5korH6t+Iq
eNiZUTUnvz09f5fIUGQBEeN8SooCrJfKKYIQouvFg4fEFFMAcjrXemyzZpzJgA41OY3siTqfKjC1
njYVN5KHKmvbGs9ArS/U4ZZZROY+O8xX30948xKV3UIvnPBDd5wKyEzUfSER5lUr0d8gJgHAHrk+
z6EPetsIBvg3VnPNueKH7Xhsb70u8M84MojN8cdQ467ZdBJOP3MF7fblE/o1s2eD39bfFHjG4lXN
4SAczM7atrHp0NJCsUCKqGn1BPBl/lcmTU4fXEFmrAqjK4lkJiOT+b6/Gr8M1/QlB8i81EI9ckAH
7+yrfYQnjw7u+cEpIpTyn1zCX9GAYNz7enjLRc02Ksm+N4Roc2sVaGTbgrlvWhhrY+MoXPLCRv6U
CWxbM9gwJrz7a0/5rQCYm0O7gEN2qig3L71n+7voUwWNB1bt/MplCf+2DcUcGpXHoG53hi8ybv7s
rB/YFcPOBuAky6quj0yauxLju0eeqy0UsKxIuDB7JzJONmx07Iyj1+cOq0FC3QMKEGM8fobY5q6S
Ti7hRP+drydENaw/GodKAsrVJyqvXDQ7jOu4MmjlbwRETHuOwNXHXI/k1HoENYE6pSSYub8N9MAP
JDe2upzDArPK7mffO5S1tr7k077NduYYLrSP7JSZ4MruocnygBsde0FlibxASU1jbIrxUl3mOdpu
PR/fRvMcTK9O0YYBWCeKwv5sRhOuZo2vDz1PLt+jjEbRjlxCwHcRjDrYzYJ7QVw0T6pDFEyyT9fH
+4XABlBQ/ioFWbYA6Z2UvfgyVULP9R1GO5xdEa1b9F6fXC/+EKGJKM17lKHXWj06WIHmhQ3Y8Ot0
F9PAghkR4jUPKVl4djo2k3eYQoisCyXdJlrGnuTYn7M/Cijz4rVlNK/WfmGBlbv7nukyTJeWNw4a
I4hjSy7idB/jI+2bYzgclXVjw8+RFbuGh2DjpakJ/pJB5CG2Qi/EiVL0MN9pghFVS7ax87YpAaKl
1i5d8rcvvSNnoAqt3ARrYZvUUKk3tqW+4ji0/anIeqlF0wPK/OZpMZC5cCEHHBj+4rIinH5YNiYu
3h4NAuGXv6AYXk8xhm2Itf7/WUrB2xerizgAn7dLPycPLV4H8y6CKuzP/4PbG3pwPC49+HfE3jyo
L0nXwAMwm+r4E9Kh2HeQ2+Zcc4ZOZZKMeRCraOZlt5JyfLxOwoqiR0sQpL6qjBPl0zc0d8NwsvXA
E+Fg03Y2ijJK30GlKlOaIsIs3XJtyPCHufOptwFK3WbpUzF6gNDBZfJOX5E0angOhDAjKgOmGjCy
8YsIB9cySKcAGnNPADnEBMsOJFZaS6hfvL8A80eSbYcR5ftKx77L9EuPtHV8afH04wPVsO72A9Pq
RLTO/yhLNqBHDjWe1JpOqQxUblXZ0JNssjZJEjtGPSdecSHfvO/GKaOOY2VXkJcCcInKhA5oQUEU
jt13VopRmBJX6aVBBELGGrz+yf6e6Dsuc3ghnHoKAukaNH+alhm0Qrtqv644bs1kEuLaLiEwIXeV
/F8b67QXwpY5Vt6WH6sjkQa3nhpB5fs1jrqCckI+RZU0sP0r1dQ19ByS+3IHGWXESuXgDmc7g7Tj
fvW49K2ECYUW9+KmVDBHyiqNWaUcTKpJRBzIi31Mg7rHvbe6ohkCkFE4EU2A5mGYoc8YO1C5JFFf
7L6YYKZpo4nRLjz0b0NO06N85d3aQZAulU/5QU3mMyur+5qGkHBa96jiDynSYLVbPcw7lnXgSYip
vpMMKYXnUxX85LFQ/vzYejlR8Xr5uienPJOjMuBFG1b34lmbirsIi+PuJmFVOaJxUexGz1UQa3Vg
VVwKpcho1H+xz0EsrKKJ73lfMfZ6iAty7HdO/77Ki3qnDEGL4iDHLB8hUyuL3rMd2dNR3/iDbVTo
54kOzeHHypBCnjV1mDbnOgiB9LpXX/pzbrBiZgG8JWOiSSJzqgh9HjI09k2GAUVSrYk0048F9Vk/
a+7ob7vUNLcfdWCqtSIt1Tjf1NLM9yFF+FuV1aLtT1RhCWpcT5qNT1f/qrMWSOOShUWLXGffYAvT
/IyHQfk6LDZCCDuMLZZf+JJ252/EXwMwj4R+nbCmSi21TAWU2C78H4j99HOx6eSugWGyxYR/z949
KTf2WuVckgP2toJvStVPlMK9WXrCzx4VtHoQ9ehdxBgkt6YbGP3xZ4PK4ukyeo66SvJMZwyxnYjy
ZbgJ2wOOaqTbCTdQ6SAryFD2DLbLG9scx+VtsEdi8XTz8WyHbNnldgWfVKtUUGjWbmYyavhiKhq6
u6tV6QW7HFOBJZisGB1qLKiJfvHVr5AJnpFyJPp31OzfP2eK+oI0jxoyusc0057LvB0fa758PLsq
Wnt5L49YK7e+gajV+TmGmedRp05vv+4h+T7MZ600GYjZxzdFdwlvzD75ZzntfRZmIVLDQbdP6ie6
plSf0L9jSTdBaGeM7BzHPcIiQhqlXJdnJr4y4NL3X83okdgC1qm8qYKdMkaOM3RMu5VCF9JzNCoJ
Nfb6ICgGpDtL9NDa8Z7cw24yRd53Ro5FYjbtNmpcqMk8vSXzjcwnGLuVP4dn2VgqI8AJTG5GpY6E
/TjGetSehiOpPPOixVKiHrNBXLMgx866NKOT2AjNUc+khSDRuS9WnrYv2fvrMYGnHZ98JPmsihKg
atfqkkM2lk1oLxIDwMjhKs+ekm7iWyXy+WeGiokVhN+xTY2j//G6EMOq+V624OaVjtmMngLJXc1M
EHzcyGFgkgioXT+OdNRm311MNX895twdegqjv1G/t0WT7o9sp8zUGHXZEtrn3h5vHNUZM3jj6f1x
CihXixYVScSv3UeNWMWPprUxLhcrGZ9Ey6NpA7LaxSvLvXo1BO3PczzMlhbBPvDMdVKMI88bUX+t
Fxc76oyG0HWhVIhJBMuRPUUIG3JzmZw+TOa6S0MnYs76z+FYDt+vhwzO1IvZUErpRQiw7c6VOkwI
N55DjKDLm4fkPfbOJh8Gbd8r8Bh9P6Yyv5q7Bja8XZLFfcxyJCSbW9o/fUwJOZTRLjHAfalqbvkj
lpu3B8e6ELCElkbogX+o9DhFnN2IsE4Gxw1DMW69EclW93nvUXzbNEN3fYcoCn+0bnebxdLIfXQq
ZnvLfZPUbdI5GBRYR4uk6pdKFUsa6P1Cv1okxow59T/Q3XwKO7gD2AiUhKJdOz7CUR7e3/TI4ET+
pCkTaRlpgyaciSJdKeCAkUDgRZFPlKMhDuS9alKV5zDa/GIo31XwIsYNNIYFawav1SU59OanPsYS
83gj/wk32fYsKS6nfsF79br0TDnn9pRtlIodII5V0T5QbefZbl10lL2FkPr8a6BfW2tHHCp0KAi0
98secNdsrGTYALrtzK2dyrh+yoqXYqeC2yfKR+mphalOqpiGz/Gt/fXezb2NuSG3JoV4Pl11P5Ab
kd+ybUgzD/N1/Q3AeXUe1hXDThSfbG/R5ayJEHJBTD2oRqsTkhVCXSWjSMa/AO3etOrMqAn3TNHn
tH9HTKTRWWSk34CA3p8l95hK9c/PFLYzseTWb3ZZZ7li1dCKzc3B3SrIMTrTaE/VjAC9pBWsM6WF
mBPWTmaCwOde/1dnr3mmceZupYgVij1l0O5mIudb88OFdFEKWmrHoaHcmPjHVsCQMAmqbRJ5RegQ
0dqWBQZ4o102yu07MgGpCwHzzQn5/gAW0QpJCcJZKfy1MRJOXRdMxRDU9sIFs93Zys7p1+jTZQwV
poxeCh0rUlyi2rdF3PY/QBNGOu7W/lSU3Kyk7sJcs2ZkFszT4IO+M2OeHb3hPptlVLjQBU7HpqCj
sIV91P2U5ntzp6x+mco0KtBgVRXmTGJFgfol6EYDQFQ9/CbPRMxutJ3GeKEBPoWMXf3wcyl1j2KI
lUxe1GuHZGOquAC/+NMpS2g4i20QbLQxjbpi/WUVAw1rtt5xqkPjVVO/Fsnyx+1HxkBGA1R8E34e
jBVkR7xuuQx84XvFgJq8mLth0LWkDquLJ+lN/fBJGfwYwUfvkqN9ymHWWlwJDJU6Iidwnk51w0yr
mOgbMIsEJRhV+ac5zZvtNoBc4imXapYHkzIpw+xJhDo73E+hZHzt8xmY/CW8GFLrLfk3uoeBvIfN
Ys7uS00CoA/Mai1gwiUs1/T8HB6tpKVVkelw1z7EOsCe4HcXY8l7KJykg5TyWmOlDcjSi56go6NZ
5DYNQy5ik6xPvwosUxgRAjASHiGY8KaLISUnvgrgZC5hKSCjFjnh3j2IluiTq9ITxttsb6F/5W8s
PxCl4rXMFX4RX+i0GvschgROy+IXyj0RbZppt4QAvW4208VdBIKruPYaf5KFglAAzAswbVjN9SLS
rqgqD6lh5ZOd1eLRRSyl3bHfoe9GH+pK4J9xX7bBJRXC3pfKeKxNQA8GuhYp5TOFAacI83algqEf
1Wlxz8fJE1icl0TscWSN+KDoIyp6Fv8TXK3XkeQ8Iig+cFNMfkEHaFY3x9xtbZt8k/KkKOejvRS5
PIT8qwvO8AHIKREnsn5GJMnLvLKyk1oA/0hNMRt0eC0SW9VK29C8lqndcrxRkgP6FHzVYlwK5o5u
p1eS7J4a3THWpx+r0huvPCwfG68bGv+X5pdAMAhJXrLi9mCoIxkx5v6sXq4nxS5WUlKFpRxk0vEp
8RvWgCCJW0FQPL+jP1uUZHx31+IvPhcAjUbxsKOSHmL/rvLIm6hAWpiChbqWKfOAlwfodPqp1Qvn
Itj95llEsxMDpqIIXXbq6uEXUzO/cvJMKj3PrlSv9+AJSeln7srWZjjwGjP8ucqa6FqU+MULUsZa
4y/5syNLFZSpFNzqdwWJUK7oF3byulNMcowjlqeJku+DThhZuXAmL23XmwZXAVADLk9KqxObKvu/
5k2suFpHh0nfClHP3OZMKE0uFwdmoYsKqU0gF3kdEzDM3V/cQaIB1rsgeEcbt/pAhLdp9eaqJ3Aq
MXzG9wdYuxqTJD4OPDC7Jewx/P8PzkMNyIZW3dsbCUdmGjtLlEAlyTOTToC4VfazEeOSDtGmjNIZ
Cqd8+hWeeMdc03Oxs3AXRpMiQyMWV0jXhkb+C8hOLQjIltubYK5ODIVsNUoLP51NWoAszIordDTJ
OZdh7xvbn9MLj2cb2nednWnVcbVWtPM7njGhqOaE5ONuQfROHBtRsfdSf5nSJAgJpXmSZmw3EA5Z
FOZ9AAfY2HRUfg2L6dgG7nAW6BQBGBs2uoFKXYjSMsM9r2IRpT4caTah2vbm3EmX95dzyV3u5Nbn
twbKfrEJSYmwfQN/vhHwVWdzBDVRi4akKfY3OEQY6v+XftbK+rY95SlvcPAQTHZFlJPgPzNacvr9
9mrSVhVgivPXMgxucj1AmPo9zlUlRJTSekkZ+H+QzAeCD4rwlTh8yKr48DV3r3oeeRSMl/biQ/Os
Z8XaqXxWt6why8+4kaQJUuleehuYH8itf4vk5HZgmewEaql1UYynrwUCWjCi4l6IlomEHyunRbE+
mlQGMWwoS3mtgXeu28HEo4l5iOzLwES7Lmty+Tv4lxaqE5YzK/sBXKKhiZaaaMae9RFh/2LFahFw
CeJQCpl5lSEvlh7k0jwaSBShS7odZvT3GJHMIpOWxw8i8CUehVagZ0onR1eH7T2zm2FjwTN8TOwu
NepHtkMFKqBm+zBE/Ug0O0JBKtEeXQUhjS1p5S7arQr6r4zYpa9ModFuMZqyPgVby7q1PstTTXm8
L9CxUWOzhICaqYH1M7yn6WcRRN3veNVdap19DltvyrK4GNd6/cJ7Rptt8XhV84zlzEAbZqSCBlKY
a2bm+y6Qo16Amu6FHifRKrzDuciF0XA8tXcA6HwGaayocLu8/A5p7D2RbfC7Fo0EhD6OZwPT1HaG
YzkLL9bDjI87ipV9NDn2OUeEyLwcKt19Qw0Nj5zbgq5K4hgHdGNv+rZfrY3ZbLtdPMF6JEKOJtle
m/6xhMvKxYJDpwFr1oeqekL9il+/1nKPNpA3dpHJ5SlsWkVYOjMnzxxfSK7phButjqQHsnFNUcgZ
dg+oUpXXSRyPhEYRns7XQhaP8Dya3t6KyoEN/PL6Q8ijKaB6Holb/hfbLeTATXKbD4t68vc4Q/2y
ix5OgCr5BprduABQwO4layxtQQ4vNdoy14P331rZ1HYX7PXaxOspPkmmPDX7/VdW86FNLVt6jx+Z
Bh6v/7nUEmegKLRe+9meAiv2Oq6et8VU5pIEvXLO5MwYUMqghq7C3N/VOBfD8sMYiZgcIjSuWTxQ
KBVgWCRFK8SwmTvVriPwHdUAT5jDVLX22y/0kNET0tfa1PK6/xoL3jrbfpv68oZBHD1HpjlruBOC
OZqA7pBv+r+qTARkc34NHJunDoN3CrKRUnlM7FBIDhUeC52fvJGN/86Jf6kvbCxcicBcTOW8wV82
fddlaX49tH6cHrCCND1OaIRC4CP+5akLrCVV7EDqKJDTKk/SkTaayOHIrJ4aC09yk3bsRST0/z9L
bWvfwgeggfeejX6wLogPc90o2wziq4xhsM0/F0ArmduEVEQmf9oM/1SWsGGam6XZqFGEDpwxBt6M
DGwMqXWRNZ1w33ZvvgwTCwcf0S3tYa9N6RUOdqJUzxnnjtz3NVwX53ZruJ80itUHFJ6QRMLCIsAZ
uNKeZH0nLLzLH3cJcakleBOTUkjXpiD5eq52xFmvIndY8v/TCkpgpibM3FH5GCvAULmiMP1R8Nnw
rpUidk2RGnpu9rb7uQ+rRKF6X7v/DPv2TcnT45UnDJHubZVsRp2rKi76PTYZvBYPyWIw1bgia4Yk
C5u+OTbDhtS2dF7i1DCCZuHJUQu7rBj/4HkMQAsiHZ4GRE+Dkxy+U/R5ucvdWXUuFHks42PP/50u
sEEyKeionQ9J5DJ2Z/vQHkfX7wTnPnZpbCYRPAQAGNjD1mnjrtEMvlr14qGL96tlGRXZPyWOOCDF
5/Zk7tN4yiJX3zSonMIkdJ5QIfRyu8VlUJ2p03GY8nH6GcToWG2oVSND5X1WDdbstKRsuqvRQ9CP
f+yjt2g8O/zwFISqt4GLiFl4PXDzTyUGdqBYTtVd9pC7lKKOVsKUO8nIU+PjagU9NPisnmDiRl9V
lqK5hGQl/ypivsHWwqjxrOEBjgz2dC/MD8+s4Huc5EvRWHbR2AteLBJIG4Hj4MazGkG9wmEZbCfX
2d6xrZC/ZHdGUZOPzR++WexRP6mEQ9CGgwJBWSnYAUGLJrhBoY6jEA+RspCpdeUObp8NX48b/J5o
Hu6YRtqOl2PcqJGVUYPjyZ0PMegrnck1Z9EBmk5Fhpc9GKOALJven+JTNjlS4vhvT+b/0FeKGGHm
kcQxf4jZ3PIJO7O0D/IL/lvJ4Ut55XTDq7Q4tGCs6Xc3NVyqUJmf+yVVPWHhT+66EemcDh9q0v/x
OdZHPpl33k2V7FaD4GJUpVU7xIEnCpgS0v7ScObeOnnhFeA2vaWU8o8UqHpB1N/Lf1B9IgzhJy+q
n0/Pi7AhTpb2n10RXnL30+hl96o05qMjYWm17E5gIEH2RAFF0GFzxieCp2a1/WkqReQ3Nborhmq1
ZIZhnn1xcXVoMCkZKC7Zn19C9pwhWR0jBSu/u9tHmp8Uc4bOvK5NBauuYpkmtILGM7w/TUjVLNs4
gP0lDX8eqpFxdsdj8szRh8a5yYk64eRBc2mAjVxu0QDG9Aj0bDwx6ZtzqWeOVqPeoAccQXkSnJA+
ZNJ4oOlwmmdBzhHvgtxLtTQ5aPCUk4ChtWu62lv03LDjeWsAxFvZd81Ki1auuW+wockMZeukFSmY
8M/H2urtj0+kfc25QGY/oyPOHB7PRG+CZ5/oxXDV7D7dysaNYWWVBqKOaS7jUWYg2QBRum00JFyP
WRAeLDBAIBzpZs54rLLZ+vN2Urjisv4pLSFEdq7RhTkaUeVpVBqlBX+oes8mxHV2ZlEjIwkI/Wtf
+XcNpEHOwksJQNmvqXebQxKiDw7SMeJ/Uj1uJuSzcboDxF2k0WKSPgu/NcF+TXLSjuxOIxaE5Me0
JSzGzbWBxZ8xwqsM0dF60urVNkr+fCA8UZPzd62kUOw9vEvGOwcK3Rnj8V5zS366GVdT0GONXYOE
Mr0IEf6slNvScWvFHrYCzWc5I51AxQJ93VdQPuj1xYiEIvo51ba9gZioR43z8csz2E4T6/MrSjmv
LDTwTdObElcoRZGzaJ+eE6qL+iZT5bFHq2dYYmzKBI1tO/6EOrY4mbcNxsTAL8Z2HzV4TR3nEj2f
UYHxHOzuN8IyEV8F1hcL5Tox0jA1SJx1zr+DjbTw6hJ5VvYBeznG1nf44YUee4QNrJ3Iir99TARk
qaKVa2If9CfNhFTVclsJNcXA6Wrbk2W7Qvqjt88XYFnaJXoW5rUOjM36w5W4bfJuTpQKbse344hE
N8w2IF8gpZfTrKMccVUDB17BVwSxDwL/uATCvNM4F2ROWP885e89886uGs3uagHC5kMc6evJvJK9
m2koCDgnFIkMm2MAHDROvOq0MdFfcE6Mv1Q6pW8xoWQKY9UQoLVNS6e3uoqBy4GCGPQnpsJuJdbl
JMKu4eQzlOxI2DU72G0ztAiHvMWt4tcpf6q3Fr+rKWU/upPu5S4bSvI7oMMLU2QZ6v+1TLoyoDO1
oCao1ffhGP9hwB6cP0AcfeaciN8OQUfhqRWfDEwLsAn+B6VEFACOxMEqKTsMu9rrERcSjdN95Bj4
groZnkbj94B3gCAsyhrglw0Ce/fkP38nTQvFsyp0GbJLgKosGcoZgPoQfDsSZkY9TUok9fuLA72m
1l8MN+jMlCpATPDqarOMxzcEqxBugmG1QF7c55Siwt4rcfXzagfvdNlQRyDm/9x5MWDlFvzHSJGw
SQglBd2Lrfef11uPoT6FZq6nX27EH0VPgassogf6hG2RygzvRYGbqtfy8bhoiyfRds/CoHoEuSRP
rbHE8ylo42e9bNJAiy4POG9xJmdJDGEvLBEy+4YIEWwcQXxfQlOqeVTNiymJU58/c1rSl1nQBnvr
EOCpnIyGKUgy+0jROTKY9+TrnNSwTe0DEDGuqRzZDbyD5u7mbIfUKl/9Fj9Ytifp1/4LOV2WUcUP
zG5qkfYUUGRl79v8RVARnLWjzse2wf8zJK3fl5yLTTKZAxAvQDG4fFo8crsDWld51OZVEegclEb1
8I6A+9nosigfLAS3P/3TkyFVgXsp7qufTXbgCMnxjCsfIs0jPjDXGx5aT3BsgqqYqhhJD3oTdSsg
jwa/Hkt6MbqYMyZrW5HXfqgztfFNz+MHQn8GQ+BESkmxFUFRIEUZq0sKeWXcWHFrh0P+u04Drnlx
jZuk+qf9tbOc/ejetAVVJ+8I+F/wBgCAQX/mEv8Nf20FPbs1nGKWBt+UagB8nVwE+4RJDYfCKrEE
7oUlQMyQTV3ysKdHKBS7hMVySLDJxHqfT5wZ9SnvKIbDtq6UTbhP/p45CcTHBTc17+TL9NZoNLYH
f9dtcgT/5dYU14F/Zf1l88AISmNa9eaYIlat8YeV4L7worjWf6Odlyfxetrxtbv7KhSjDycPuJcT
av968jtNt/5gvJg2pkQRW4yxlTX64ihwPB1ee5VpQ/DUjEizfXOymVNEgupmYq15Qy1nbFNGtoh9
nm/VxpkTdt7WYjg/6fY2SOfIv8Y7CImbsTtbVe8d2zJHL7QdBC8ZR04SXZnZrABXkMQ3ppKAonud
z5yEqGXxz7hG7bMWn+R5OqA8M32DUkt+ElnjF9Oi7e3ig0yVgFdIzMKP9UZXx3BY9eDxr25HiakX
b2Tytlqp4IEvZzxEJjnIpde9L/Kx7Ym+8/mYEy2ZrP0naRvOs6i5+1FLoZ1gYYtI6Ml69hCxdyUB
PEyZ39C4Hmzp3LJdqlgX3kqHPSEQ/oyqMxhjw9Tw9o+0FmOTpR08Gy8hGvtVl0wxrXyVk7srijms
YHEtyJi2j0lU5j/keCd86uL5nnH7dyFQzVpdyhuO2/+UbbC8y5akBWrQNZitlSH0MvhvLr1SwvXz
f0eHcF/K3xph2u2esl2LRbxSga95wBLuM90cGF8Dk0JmAjW5dALhKl/2iNz8AlWM2Q2/UQftLzcO
PP/bb3TXlEvzCYyjzpSvTBG6FRdyx/mrFWXfBahAoiYItKdo/oA0uy/hmTwW3nq2NpZza4f6+hGl
cuGTFgpf1TtPWsXTaI6zWC+e0URfiLCNxMlaK8gSSJ/0e0lvKfn6dJoBLOBn4uypGYs/jQJRn7AQ
CG18diZ+R4kf4Ix7Hk9lnNFG39+eib5WyesSoEL4ZHN8EXaTcBKM0ZTNXK3C9qsXFvNoBB8T90xg
754Kfe9YxnQy8agnMmvib2RXWFKrKCBXWpJcChZF06lxs8viMeRBfiAPyZHDnhe+003urcNN7iR/
DHEb5PtrE1i2IN1N2rorH0DEyXy9qbVBz5XbJnsN26YyYCYCxV2Mi6IA/cgOFw+bRAn2cPIEVipi
KBJIPIDIgz5IYRgkZ8s2ZnGgxzC2P61zxWZmWEU7r1s58l/5Ap0SHkcMpWRjNlt0e/TCnNWfxFrb
A1GajoXfUXI0LJsiHp9dDLW0zkW4TZpZEO3EAeJSdvfnqegJHpIsslQ9u5j1FvNiHSgXJa/5QfOO
oZ898FSUrW2GEkx2rhK5MNHbipP9errv3eAp9QCTgoFzEIrLvQsHA7SDMiRpYwjAcTBgnO8T+Iu5
945QkVm3NwGcAK+lT6cizV6ebV37ZLQQvkourVoYQy83WaF9QQu0XuL9VxrcgX8pISHNjO3O3ang
URr6Y+KCSSvK1L1XpctgaPKgtEgPl4gLPTkhhMSbUtZJECTEFWdF9e19a9bp09AvFKBABahf0VT7
e7lulSBnHCOnZGhd9x1UFbae5GQ/TFFQgSs/dj9icDl6genfCxFcbEE+e0ljKtsxrQCKYGJudIDC
Cx81OjzReIIxEPeL3SDq02YvJIQVOs3WIyC4ny6MU02pKq9IOI/q6MCy1X+j4ZWI/K2JO5XZJyoP
N4NX6znBnNTDQx2sWter/h+9c3nPlT3aOznH+lOeApOf2aslDMgwWxHB+wUEgSPAfL8QfrMyZWKR
Qxw15dFPZRkMZBN3fDBBYtEGBCNcjNpn0pfhypKW2I7l8hCWfjjaYKNZPucDx2Mtn9mfGqUeV431
7ip597FShUCCGqs2kwMvNwu1ruIZQkW13DXu5BMczfl0y4aMeKu9gDZz6/P1nIdmFGP0tuUTShU9
ltd9QXqmBX/WksBm+GRLbQGMq1p/Q/k7Iw3jDD1wN8qqP0gdepsYRi5XG8XmAp6oFLdK38Q7A4Vq
wnjXvQqej96HASbwAZiPTGsNv8RJBiAaUW28OsTJ2ikWsvC6vGweH6ynwzkkqJchOOT5mL9qXQiw
GHw3lrCYNgnWOPX0LbdSFJLmGGHTizOLC2WNwe5BoReqdQsDrhMGBi5NLMcqLPl0ZK+ouX6+HI9q
uCtj4PiOurBF0aOHLcfZKpTR2Je5ZsyEk6iys0vV3w8Hn3VJK2oDF+EXfd2EbV/c8o4LdLBvSZzO
eEDo0kSkZ5KoqSLrqw1bzH4ZTv/RnSZf6XBCN7ppMBSuLyU4gxDtAwFAp1y9ep3lSeEPixwG/doL
WSf588UuP7sZqkL46F8GkRLPygxKvhGPmZ7IvdlUA7Xp/vB+SEQ3XKxFxhEArffWWrHP/Cqo9AIS
AyS/lNjTgKu9hDMRtXYDUaRgj31+/ZGR1mUj8ANGMYcCw8eV8joZlgfMnUChhRy7F0LdpeI9/zwR
1xDz2SfPpdgIWJfbrP4pJAh2PZ/88ouxlLRmxfpXYEbdCpmhlFWA86LGoJp3cyA19fb1lNaRJc0T
cN+DKqGmxdnZ/SH2705hxqLHNScmZ5CMvkHhT5Md8GrW54sF2raGzvAaolgKTx7YmJUA67J3cf8y
pB9Zt+Qk2q4rBR8tXwxFyUHSKRMzn1Y5TC2r5VtYKaPhemeD4PXTYcbnHGjjFscMsmGC/S/uHVEW
WH2oR7o0M9BZyyHp4kpCzmddhRjnd0hLCQmrtNivVVlN1XIFsQRELvUZW9MlzSCuAlVqMoFrq08O
Ne3smJ98F1a+KdfpUoAqBorc4yuljLttAkRAYfLxvKQRVc9aBK23PuOMOE5h8NtEVDj6f5WI5wxr
lUXm826LVIlufpmm7ntE22v9GPqlPCPAR9nCpMeU2jbf0bOvKnEmce687pnzCTiSD9gew/fiTDw2
93TL4YCFbjWyJNQ1vg7hikE4+sSEiSGYfAhwe9jewoWe5WfKUP9IOuID9uu/+ofeKgY9ClWTtJYe
9rqNvxXNLOupeRCV0tQfxaIRux2oV3UUDPGLlb9pFM3PHrw/Dv0RFs1HsogM/s5+8V5AJOBjeSdS
bGFvEVZzC9yvuIg15h7pBzfsCNwXb+fWy40jftg39YbjgyQn6fSz/AKLbHh83COhCzW5CyEyrstk
gIP+crhQfBhkviFYD7kv6kovJehxYk84Jy0fkwlx6jsu87TvH9InRwCLAIiY8Dgtv89kt1vVrIKx
6G5VANm85wVjgX/eiee23D4A8eSn5E4eIPV0qKxqSdqZV1HxJriIMM8MxnymIdkz+oY/t9cpxXB4
YGV0lHUhlHp/iy5tbyYdSpcUYHMDjwWqLozOfTorsZDS35hUHkfnj/l1+Qp0JuRuQ0I5ZjVUV6if
u8MKHom3vTlzIL+x4iAaC2Jy6+Ynt/NydA3iCCMAEJ1hfhG+0Mw7gekgnEKAVETuSd+UoEWQlzUj
i+GlYR1tSzqfy5RdCI2OEyTISWvcQxfXxJSO/9t4/DRf/OkASeRAYyXvP6Ml4PKyX0j7Oi2wFC9b
3NaKMm0yiJN3KMSajsFOIHO3C1Xdsku2CiHzImr4D2sMQgQJi8tjT5FwupAbYWtZX8HBEMuP6j1n
qmYLYst6dN6v4w4B7TP9jlzyS5/CwovpOVaO6zPxPewAQuenPXYm/J9bKAKS5zz24I6n+GxpmrTw
r6NzxEEMPFUo4711fPUKALsrsk4Ie0PJVj9EQPcM0OBvJOGWvAtvwDdW+vAUhIxU18HfnQHNKPk1
oXUWlsKpAs/CMqz/HtQIhpAxxb8jDUkZ1NSayhh12a/bZ1YlsFP3NSXEHTVZft7fooYqOS1UONkz
Xn5nd8ukgvROKwRgwMBl2eS1fJhvGPS+r9FRUj3y0mJ4Cbi/qsMIqPOxcM7rVjU7WB96TzWcF7MG
Ocm1jXm8yOEBPjMs9FBA3nvAqBFDfA7+EYb+XdkUHJyP25/fYWZ4eWCXxW8ibzKxElqtZHkGrxE6
xDP3wAumyg1lAbt9XZAcUk+9kJS0zSSSLca1IB1cNzqUl1OemfRj07UqSGSp5H/bt2Nso5CuKFGl
J1N3fj47n2gGhVj6utitBVgv2j4MS4evEjrRqSAjNHWAvkynBg2/c6lZ7uO7/Z4KJ+U34c5esOoT
FSmg0DTakuH/DJTJN+lT0nh1ki7KOLURi8KU+Ww4PjM6GJGHnIVJoh973WWZ8FEjYbCH9RuYcp2D
qbc1U5K19QqBRjfpRPi8Ul4XDlKZVm4avzLJWZFNZCHyrkFmRRgT4PrOZIq4oKLemnPFzYrt0f8v
Iy9W24bk7kJ1TArQOfBkE0FmSu5UYMwvyhCgXXr8O/76yZQFzOsgVBbnPwxs35yVZiHd7xxN9SNc
EtqTTLEvHlDThL3AsUoYvvroDpBGZC597dq9Ia4IktJwwwu7EJrjVbBMbJiahJDp1s/P/k2wHK/L
5YMl99XV2kbxsUBK2u/DUexFHRQz3X9fLEi+7WVu6HtnN6H/L9tuN9YIirVD+ztEnRW/DN6tDKcz
9i4Ei9Agl4kN3LhX/BtrkhZ2eTQiwTjP5fIxiTipPG4V8ruM+lW2aC2E3ooEetu7MN1dQTEJMid7
ATwIcBL6o+pG+6XDyFFGgNcBxLLYNk681B1dwmOrV2FeT+52OtQ3Jm/FULLkbBXr4XM+VoRv+j44
2dQQogSJEqZYAM2EYAEmY3YyeufOVIVsXB/N99qEmlZrsK9MFf9NKtrQ3KdOk7e+jOM4uvN83ugH
hVOsb/lCqzQten051cMGmteTFhOF+FSqpzysVe78e3eVTCIZPqxf7oSbVcZrFzLxrGG0pnu+6hT/
rb1jmPjHxP9utpch+J/oqchPvNBah5vG01k8rjgArarZmRBWmfELzw9nDBR57Gbl2uXLr2WdYdrB
oR3CnXZ7qKrGJ4ayem10HxoEiLxLPc1IX8W0tA12x4nWjjGzQWPAIrlS5wqbDbqSyXGaTjyeJez2
Q8sD6OXVwy+gZhuZYFTi4a31oap/CPdYlDwfMIT3g93DrgE2OnLGUi1JjmCTOwysYk1hy58u5iIL
CLfY/MsHp5fCmIAEWnlC8yYVY4pLqFO7VOCxy/CfglzhU5urmAVWNgL5YgxA4bhDigsAwIRc/SQQ
vno/Zdosn/jeYToAdqovpsH1kCrQ6G5BIfeibrx7lWDGINiKktGKcNVlRIn/EJqb/fFYkfQtmpZm
MtmLdUVNsyuLwJ3Vpm314KturB6bbVLqdnCKI/g5nRYShDg149A+kU6EZYHjD0EHgOfySuc8Y4pT
SJL12PyLBrjStZqCaSLGVoFEdXOw2/+YEk1zIZKqilecOLVnabd47VKrZics3YYO3GnhlraA9eNj
/lOp3buQRUbeVg+SzKJtEtOJ2dwTvC0VpBXQQqW334Y2FFQIS9DnPn8GxxnX4XUGvaRPwwcvO010
WLiJlHQ7WgFb2ANKmenF/TKOFIdAWQEyvo03T7pteLOCqK5ZEF6GxIE9cAxSKUF40B+JgvPoWpOX
XwbyDr7Ii/HIZMB7jKDyVwuyjts1R+4h107qiODScgOIv6n+fga7q0FZ1ipQ1TQHQKDGdE4XcbpG
RRo43kqRf2NXeimjWu7Hf3vw5AOCpoWshseOxEguOGm7WtsCrl7nCewZHKew2oovRvOgDlhqvMQA
FWnGfyNGzbDa7JZw6rez10vc/pKCBbTABrX6Nk94VxeRzZse6iNAp6aCyhTluUgT8lXXUc331PHL
nZGGs4YB8yFlADggeYGkAvvFqvuDlxg5QYyWGyrF/LQA+JJXxISq9pVHAL/waGSzuSBYo2d7W+Xc
4fjUBvu0LArxtq8SeQEmxyrp8XZPol8h9SRpp6MlTDHerF/rjFhNJumY3WJyKKWrx9vPDT6FbzZo
u8L/gODV3VketlGjWKHsujghz91/emafasnKaBu1nD/mOx/1cTVR68vRWpB+rbETgGnb9CDP1e5E
tRSMVCTwYwWW6NWcATnfkD/5Awd4cc7NwxIG0CYpW4qdRBPspWXI1zEjK9iJxt4Me0CnCNpfbj9a
YV+dMezJTIDVSHNv1SgkvwNPT3EKrG7zq7KeB+zitgyjcuRxMAEIeB45DRPPU2kKAPH9wqDoyE+/
t0HsqNQeWUewBtadWIylPyLmbYZqTDHh2edFTwHRMi+MoIKl8joqFXR0ss/Ue1dOgE8arC+8KQ1M
gg3+zxW8arcO+wR4RhTZ89JWpeDBFiGRa4cAPTNFkubXrngpf3KZiwKe6K3rvWkabvXsq/7bC7xR
Zo0Y7pSqb4oy/CtGqfQ6OmQbqMcmQOocw3oqvfl0O51/uzD08lN2K6uJIWZCecuvWcLkjuNZMYqm
ZuHyrEnCPya6T4tIMyBq+sRlYyBk/S6PxyD9Gq+JRJgiQfw6cJGoMGnbzWn0rSvyuGf5ybd1Gw/e
kEjafQqYFaCOrBmjY5hd1RpBE8T15j+Rw4ka+2ZBihP8kJMAROfBxYwKl/fR6Z8+jWk+AAtb7W26
K/sHpzq9vTrkccR66dXk+TbZtNQTsEYbteLJDnhhWZTIpagMu1FT5Hgmepv6pj8jjUhTsAXfSj9p
uIZ/dWVJJh/DQqsSD2ogQ7Qxyx8DSnWVZ+6j7laSEdPkgi3omqcw72sO28bMpv/EX4tBgY3aNgDj
RJ4MYD8bSHlvzmg6L+MqaOMtV4Ro8TSzdrvVKGV0n+vGOALp22Lu19ZKXHTH5T5zRMWLfCU9VPCc
M9zB5Ua+8RZ4XZdZErSKpzAzUR7yXQygUPB8rhODznBddF+S/VPD/49Lvn2pqrmUFjO4ZwfwiOiD
ukJaQBwyo+fD0jCSu10CnM5znORZd2EYzraaHXcfUKKk8L2dPyE73sI1BwjnKH4vXJ8tG9viPido
G23MtXT3lTmYGeo9Zqr8+VThBADnWwDIvunG0FfCzxBS9LG0u6gbxemmmWvNN02e2BLK1F+82VWJ
snwZ8wQxRSxhYIWZLPQpdFE9qzuu+Ui/fxmXVJ8Mapej/aVmoi+VNfXFQMYycLnla+yMijvsOzlh
GvhuK+E2dgvh3OqRsTVFMsWTEkKjMI8dP4/defI/f0zYKViOIiskKzgSOXFNwBQr4hcynL0jrFst
MMyJb2jO/HZv2O8qEyLCNv0t5mS0CtySyH2Lx4POeL3xKsdlI/5FN+fbmT8N4tbASWF9sKXM01Dx
jhyiaMeRP+1JCySFSVp67kdb2tl9et0YSE21PwkXj0vai1xKiArPcZD9GtK6rRqWfpXCx5usuPeV
3vek5Ox8aFQP4UNFpRtCgaZD6gNJ1rxCiWJEPyeqw+f7wNezmQDVqDQ1zMfHTLXuCASyjoimbP9c
HSRI39YSzJuERXfrLtFBkc3uZS/Rdg17JtSUepqJ0lHhpm14i99jXrp1RQRMAzJzAWePWUJMPsO+
trVjevTCajPyB0MLCNXxvBezDlVcXM3hk3Zm/vjdTdl55Osnll7gbItgU3DXByAPX+uDn+UG1odb
Y0Vpl/zJUutDCMbKU9mUpb2aB1vpgU3nKPJsodQ/hy7FcJPQe714mx1ERsQK8pCo1P/zxFQvQLZy
piByD5vK/6iQF3g3wKaxVCwP1rnWu0zJ1rbFz+dW7zdHaW0kQzzMXFrwbfaGCnkwyoG+ON1ZnS5N
2lGqPZQ/QYkXUEAVQw1AzBNVDnXwBTS/jLkrmPLWHJjpUQxVS24o4FjjvxhxSJgrehn933VQVQM/
Y+Fvj3s/0o96VXVibpttyuvDZSHlgwwAv0LGfgxxqaZ+qdsjmqC1xmgBV6IMWE9O2QFvd9zi3tX+
m1IUzhFIYKdQ6+UHgQg90y4SN5bbYkUAp6jdioiKZHD9vrGUzSfcnEtNHE9NY7J600FacJTAyij8
kSa8haXufoWt2GmwyeRJVlIFl+gTzIGhn3Mc2kbWMtPrGY3EFdWFczyPeAIZ61UoDh5T6slZIQoQ
u7HKeyVgSOpYngwz0gkOjG2NmPk0mvFSoI6tjIxiBH0iB5SEVm8GBy6F6WOYhvmU27Mq7GICss9e
HEfwbc3J6xu/X9fnermBCYnxbQC7ieVJ2wDP53vpiUFJ2juKlEsdZhqbTbB9HQPTRVmE4ZPK25N1
co9XOAPrc6exGzL9F7plgopEO5Hyj7V/wnoL8UXtN+x7t5XePNbn0kq2+i5j051u6Th3ULUYBl4R
ykeCsUMIqclz52PB0ycdxmv7C50Iv11rCMKy5m9G1TTrgIZkhPZ5N0ci50FQUpMN6DT7viP4KyIj
mceX/Da0cs83rroc1YN0vJdlEXkDDkDFLJo0C8biulJagtqj8A74JqD1pH9p69T8AeebUPl7a9VJ
v6kP317IMQk/lZTL2dulVN5lPQz8QDP+6TuH48hMyaxR997mdU556q0Es0tQUYJDsJEBH/QWqv+/
+W2JmTUX2oWRx5FHY7O6Jtp4AyEUjn5sGKFvfwSSm6ol7l0caKN5NCO+k9xeA22F+yqwoTQk/qcK
r5UaUJd5MAwTfz9xNK6Nvtwh1IZcG6+YiVxtMxRTv4Wg68CDUqmd2BjWSqLRsYx5V+flOWyvVWfe
6bSDVFvnVrP3N3jdzQNYSDtOINw0idjd4pzigqC06pxMXTMuOY6w3rF7rf3Wz5fcn/q65Dwn3c5I
/Ps+sCtkVYfbx7UQxDPTnuPLjB619hSgvwMnGiYBM7CmIG/d8qQ+ooKQSGdtqq3su0mKzTMgw2VQ
x+CLhbTW621qWRnFP8I3uKHfzIU+JCgFMCIJjTFLaWZpqLHVT7Ro7sKl5xEe74wXF+KVeh21JLNw
wKEnPga8TK7oIjOEFGYOvYLUSYxmAVF+BGXuoyxKBqruAFzE1ppFBuTFkDDGGBg616HOoMIdM5ek
PHe0tBVRiNqbJarMfivqAwDlHr8aXKy+bRH37xyS9saheeFhAFNxbGayieLt8lGojE9xT/ZwrC18
cC9LMAvzGScWyujDcqviLT0wkkOjPIAo4Ns1s7HiVpdZJkc14hnGQhmbeH27rBj3EDwZxjtR+Aif
sR0hOPUiD0U/5McoYqaQOderblexCpMmJOVLTzWRjnMDbn8Gb6RT7psD1hTilzZAGfQE9QAxu4Ko
xCBK8SdCAi3+ErdGdc7Xf5mMPghSQvDjhDQVA+Hw1Yt31suLo3Ln3siuXUh/mbdJodvoVPnqoerm
m2yg01sBkpqgkyeC3GS2f1rHBDX5Ft8UIjFULlPeXrF+8HNdYV/Uz0xSkNktIblweJ471GX1BWIx
g1JMMAoeO+laQL1YWkkbaA+oNSz2lonjFXg+epFXvUh+GVwsT5Uj+8Trra3EjCnpmVX6/bjlm6Lh
cEjUTtfqHTKawPfFw8i+VqQYW8b016jGJinnvrKeJEPoRZTDZVI4/2ErbdsH+95U/xqF04Vh+OTP
DN5xSR90Y4u71VK3S9AZQaNZ4oiDDRMTdwNMEy3L+Be6ZbRgw35V+dQaUBcw720lnh5nJLQR+q6Y
x3xlfZ8Rl+nC4lI6QFr1iDDYhHzc2VaJ0vOjzv6oHwM5AmEgM4ytWCoNvikskukfVUerqtlynCWd
fmX8aGJOlhyUG3fDIs8Lgdjz0iHKggfoJacOKBvUUaV0SZlrvMlXa+hNuOocAhz4T3P4MRsgyqSu
KzmvgZjYt3XCZlhXtFepaARZdJ5KM0dcAASrXcbiQYa2KVEc8m4yjYiaXX0Le2XjhPc7RPYeRfqe
crUnJeKOw8WNEt4jNzXDe2pbb5gLChML3TUbpvPv1/qTFv2wXdbxMNOLOmdMcTsWXamO3SBQ28Bn
2ihcTeB6V09HUICiuYsYDLGAj7mYWJdTrgoLAcfBMuDJcpu46zXllJbXMSMt3akOdJabjC6g3Tti
G/qg3UZm/3i6L+nFjLytbG6sYUpT8pxCYpYCPmLOLpuH99eJhnxDR4WWZxCg9fRS8pCNFuqnCZ4a
duSk9D5gxck3MXrsTkB/r6ZySZnKS18dagSWn2+E2VR+zbxCDD/pL4ZF0XX50BKagj3V0IPs/eGy
LEey//eHRLHmTB+hcW0ock76HboectLc/XMDj+kbgQsxFyW/Dkrwjc7WPqEiewFA2EulaSXCfZrx
jKRqQHyMtacGlMlIR5+ZqkeZ1iEjSHQL5NnZXpEzzLbpLISTHzZ4xFenGelG0E+3zcE4woSiiKB+
2A7KEKoz51Ai6yydRGmB0CXicdfyjbDqP7e5Go7caA2FrkFLPvdbu7sB0pQm4R30GveUwYRJPRjT
89Byotux9fRmVZo1Egt8JSBGH8O33KxxC9cJQXlR1W7Bo+BwStb7xO3nGV29VbCt97dTFixU0kw3
lRk3pPrVRV1270BC3zSsnSorsrKDM8YKB2cfPffOcbwE3n65V0NQjgByUNpcjg43OZ/pulGya/ia
x4OsaJ+ooTDYyfepxeV3fH+Iq0Qg84kzDdLEmoeQ/uIR04DXUqWjZCfOmBsHLFkufUAc65km0wex
hyZ3XUccTsMO6qvb3vsbPPlbN8SCjdsjZ8pNwU8N8un/8/+X+pH8gOlwHcagPPTSOaD1Lb92GBbh
x4mMjseJE2HiMIOnd9X+jMoPqLh0B5eXkKUz9s3yrV6jMS+5RXbLGn0taUCFT87WCJFqJDSjwOkq
zIMT/6p7/bF9W5X+L8Ln9dzu7OE+zPSCmK3fw0dV3PKR4Tkny1IetX/QshU8Q5/lluXyx11xqZAI
VAGyWfhH7hNN0iXbFPEWcPTMuzmPyoCXQF/AtjRPIPorlGA+49FA97U/iKDvHxKlTKhdA5EHPjYx
Lr+TMQMQrTV1xthqLObpbhxXWKGeY7yooUv4fAcpi/7OzgOxhAy9SJIaHpWPkoGO3v1uPE+Pod67
TevpyCzDhv7dlgtw0RBFiOUtNOejgk+K37W9tsyAUVZz/bRP+s8orAdxRUUyC6JEEoODWDRarfRe
xA+hh7x/Lm6Mvllj/DyIi/9KprTu1J40oGOAL69KowubKq4X52B2ZOcC42qsdNQa05pYG1sJF7oE
dohd0Uqwi/gn3tuxqlNZQoBKO42BeM0OynNwrWCsBaoYv4ZANf3I8YK+bDblosJhRxB/V5/AO3wO
DHObjD+cC8FL0lvcM4BD+u3abMXW84qtdqjaUgglh0RQB6yamXN0PTYQX7vgcsUZLtVLzdJHq67T
60IGERHdV8Kmegs9Nbqpu8PGD0gbH00LhX6d3KIGXK0o3HdTT57pHdf+jWHkOYiRTBkyG50uowvx
aU/tpKRT2CqZjScQ8mh2VgFMVTvvG4VB01IYPH1UWwflB6gY9LSwB9b9RstGEn6bSLw0qKB/0Yi+
o0Q/7QxaYK4NKzPFb3mxGkQqmqy3q6LYdxzc+gIBlpi5jxhvEbeS5CsRINo6Me9PwF8tZ9MGzMCP
DMcu/WMGLrjRjzTxmL05uWXN0dhX35TTs0LT6N6yDLvxSP2JIB0cVQkridTnFLLHL5RnEBl/kt8P
Js3w6LQgYh5Y8+i7RhzjuzukwqmSHzfkdDSCxYsE4cimJVpg3d32EVR4W8bK4U/AnyH9iVb42hiP
FnM0v4H3HP/iZ6KGSkO6TQLNByCqWLWyYoQ3DW3aDMPDJpdFmlZO00p/ePNo7w8nXSPRhfvXFyno
dQV/jAOJcPOH7ZlwY5/i1oBE8/vJTwGGc1BOAm4HzEJdgrvkKnqrAf0ArveDmRfe1bGQvtV+KpUH
lvdfgpm4b67PNNP6bdTtnRG7IP3Mz07ifVdHwwUTindX6+4vzKiRHBrQOaCga+41Y2boTXVwY2M+
NB+ukwcON4NuCHCvYaODFxJCjeuBLEcMJKtfRQIyF8ZlT86gfiFWAR4n/nQSUyCWr1r6zJxQJQZB
S6ZInDWsKMJZAvz5WsECYc5fCcwoI/u+dOzCqMIXDdr+MfzUgoOi19AuD2hcj5DNBEfPcySB9X5s
dUazJP4Uaerq8jEgMmLff8Cuu22e68dyZlQJSvVLXgQnxqGj6Cd0KiurK/cdSU9k7RLm3WNpftiA
EmnSHTwtYYyY4knP9tV7P9d9gE5JPvDUOhskGtPOTNgfOaWbHQq9DH6VR48DMUNNzUKYzC5NSTyF
LU/z7FgvewZBNqTdW+NZMBd9QgND4XfIgEW8r7pCn6TvUe3uRp+qSNtMZDKCmeuyOejyaoFAmhs9
ExaMsGZtwv2O7uk5RDvp9B2DVHTm91opstasNIiecZ4XOXOx2GvqAMCRvdM0Ad1VhNNcbVamxX02
Y9gR3iFEq7t9q7hMe5NVcruHMc2atORSPHCwriZu2BUXZfPSPF2ndYo6/VFadNAgjdUFvlxbvvmg
fC5d7SlYKj+elAdXbqbSNgCpS3xulDFQtUSdiL0oVkquMNLUDXZPyfxGVOr9O9TjQ/SIJdMtzMCZ
cmpKkCSBhmCVH16fKCt327aDAO/7ggikL5N5h/SfhcMvSy16R634kn/ckoUf/H0RSzQJjehAbPcI
V0GQrhtvZwt36Sa2knLYFEJsdP1ukzaSqYy/rIQv/UUHYpYUof6qGUs2U7ufZGRQB/r2ZM14wkPi
kAw+1YhuB3/qIVciym3Kq68v3DNk4ikVbRc+zE202zFhhtpOrbpYvg0JmaOiCThPYLRpEXfRY4nq
vM6nRPlJQZqKs6lu0zT57HJ35FqHLhre4HFZ8fezoatafUi9Dq9u7PKCekB06fb6Tio+R6qELo+j
0gg/MF+MFLKNTonpp/1I1vDABaRbwV0vkq++aqnlGaU8GzEUpytVNAHCWR/qRyndHNfQ7rIx6D3Z
m6B/J7Suc5JgT1k35iVoeKqujcUwtlFCMYbuEOMW0VLDM9sA3de5ZiZZjD7ajgvL6RzZTFKwQedd
cePDmeDoBzX7kBWofrt6vZzdmTIyjjVipd2dZtcrBwlMJMzvh72+ooHAjYzjfqkAstPggXRXIWXR
S75Vwp//0Jy6TM5viKWQHlY9yS5bw3JemHDdkRmqudRmimCy/L31qTNWz9bY79MrPqZUvlfzBxgt
/r9tbAjkQg+HMnflzw8UQXnMKtOyvHlqt3A9WhUvM8wFd2V6GCVMYMGnlDx8wMA+KV0DQtQhnHTb
ekv+a2+fS7RDASg+JFnYdG1vbDANO1g3LL8i019TdixoYQLxrlzZAyqfBSzyg09aszV0o18d66YH
EI8gMOX8c8O859Dc3KiZeMvJMDLWKzklMgoykdfdkxUh4sOsOHez1rCS15oI+hlA3c7Aqoc0t8da
NiH+/naeKa/M5XeC2t5OQ5+fbppmgluxv5+CV+mQ4KJ7/NLeIz9e2Dq41y4+4lM59CWcZuvVWp8z
GzwrK7AoIcxnkiK0iduTzS+N3JBFRwi8GeDkFMQj4Y2hk4HdXCEG7lFFEwVy8/hkyMP+2a2tIbbv
TrJZlZEA4TWv7R7TbT0LkWkeAkarkv42hEz60scSRuPROl2b+b+ugJXB2X5s91Gm6n0zyvDv1yYG
TP/CqRywzfgkXonYFbA8oXwBY+H5UBJzCYMzERTh6sD4CG57m/mjJzcmaRgAt1EFs3eTVKChUSlv
wjFUFZYxs0T7yxgphRXO/keHLbiEoDikEpUhff2mRnzMEEe/6tM6kuoLGcgJCWACimVaf+dlGMwf
hPmMDnj+uDm0VotuthxBGv4r9RqAYIy0b4GYBuAnA1MHTC8zDHrJSKHMKgCs1p6ffdimRiKSkBp+
9gS1SRuquoCJFtt0z0uF4KiIUz9sQYypTpiY3ZYEvl0dUwcHZkfeTrKfObYCCcBsLAMhmrv8vr7b
h9lwwa4H2jGrtPMSE7D7Y13WPhgqz/+76miQLofc/6RL8LKHR2ciSw4gjAyGnPDXoy0jwGCFagJA
LPNVWQ9Skvir63oZTlofEQAa7rX4aL70gat8eoyTGHySQuPQbPmWsQ7P6/PtrCwn2DUis5MNCNRv
XgHXub5IBGpp6YLpFgtwiKe16dSAO248DRShzZPSzUtNIzt/Nri+0ck5v9JAgEsfQhcIhBs+flPB
1Ni3ihSLf5IQ7JsUDcXYJ9kRHy28NwFrLW3JQ/WOyL6hxGZFAle9VX3KqHFKTIX2pvai+2g73hlC
FaWJgKxDlqruXK6+HgbMS3yQ1fQ7aiKWyJWkN8AMXCaGL7sI5cuvVRDAvvzvLk/QzwtzsuEqb/+7
vkdzbCJxnq4bNcxYtlGhQ86CVuxGohlBeCp2nAioigQokUUmVVVaGEarnjQi4TUjFXczF+e70Jxo
gBB4DOB3t0ZbN+4Wzn3/VFzQ8ahAzDKIvkugFqeiVnu7/803zhU0V/ISC4xuvCJKrxVJeNEQ+CuX
4Pm9CafenYtxpmBn1RUlo9YMTBmpPYfWI4fEZ6M4QNKEp+4X2IcozaCvfvDOExTdOYbf3zxd3vVd
nn56azeGBhqPet27iu2AXX/DO5pgO4IyZ7Ezk1ALgIybCY87oyCPXuxKclLkO0S+eYtvFJ+XomSo
mhyisURbgHvQHzhzpd6biAoY1cz+YRykgf1K/y4ydtwdXC15gtfuVDMF4hl2RFToSaMrDvJgof4Z
pa9x/VxdkavSFvp6AOGzQo78y0F0pguuPV1qx7K+fP6zRGnptO5QVrlCUMpbaIZeWfUc4XMWGS5h
12msVfFrbBOKpZo21paiEDIp4BCVM99FXXKX8ACDG4XVSX04jv94HbliDH97jlkXzxr8osX7S4W9
mUxgop0ITTimEKNoSH7WGOh7nxvwa09H3L1USKNdE0JlNJwxKsff20+yIkncHjDPgpQQvMKjW9RA
/wT9f7usg41QRbuTeXGvubsC/8fpF1wzCThNHTYrCc8xwfyVtcaGGdSokr9+zxTUAX+oxsygbhYb
+1yhhuq3t67hhYcNNJHEB6sKlM6jlwnKMaJXZ7K0RaqaOvQVfRlK8qwCuEGIAVmcVsncQ+KNeMU2
lMgTeIURUX5PTskB8TRTb/eRD54a8HJk8M4mk2ZTaQdTVVsO7G3wcsPw7HoB43OxZ/lhdGKyLAOC
EhCwOVD4GHWv0TsrRiQRPs5AYLTM9+aqR4PZAV0ANUjVKqDCEgsNCBQQ6PvGBOedDvJxZ/kGzuVQ
IzVWjG1ftZJBu5gAdOCVqoSS1Lp2mA2adlmh6PZyv8fyAMEQuRvH8XC3quUHrFnorApnI+vmMIHz
fDV03WZC7iwm/NSnxx+B6fgRLCXGjQk/rWa/MCEaz/rTDhmq1VKgvOX/5UwPS2z8qVfiCRTC4Wwd
7JiOs6ERfYkd7IzVh/eGsjiwi/QywWykrpIT/45QIjLuHDKqfBo6kdSqaTirFTheSZB6WSbcA+Hg
RqdmWp+MAdKEkdsd3HeXgtOyNaqBjutofLioFImd8g21p12BAzJoBF+wrbSSBWrLTbeZkA5PL/gD
l5SOljyMua407vAoLNHMkDK3wIO1C1CzQ9Lg0uQwGFtO6q3JRHWCR38S6bGbewdPJu6edyegmD5V
kiTOWJN/zc2/GRFNzieQz4ZDDWF/ntCHiluzBfHI4IxN9lOj6vHaPxqxTH5GAVgzwBQXu4LvUDpX
1IBiUqC4+ObGAgR1SCa4UDKPdKmpLm8DkuNZjE7r5ktaiLQQENNLfRIYt0iXv4wNBYY9ZKvxTjK+
TouT5Uy2pxGGjEV/h1etlsLyIXbgKWClhJrwTwIDuZdQOiBEDMa5Y539rPbHUTzxOce1fUNsnxTC
r0JQrYhl7TXoUmOMI9p15Wb1fkVwqwlfgBPoqIQj34Nq+b7p900oLENdmptAgMBx0lSKm7h1WXUw
3Z+wO5p+RV4tO+LQuF3oiFsPS5vbP5oYEbmv/BcGjwksIN0bpa1RaUD/uBrwOqvf0KFjwEv6e3VD
B+mQqr4/VP77vqSTjZ4uE+YVyPN0L+FbbpmT7wlLuRElkOGv4r3XXDpK/2yfvuU+4UoL0hxu/bN/
/mLY6tOLDlrHdyyhy64+OOKM8qdITYKcGHY2pAJGlkYaM2Ct8xBfB+U75K/iJY7NBV0p3WcfH3L1
JXXbuV531RgpDkFZmmpKB7dAolfpsYcB5YkVNvvSMTihiYzyDTs0yn4RX+zzjL3NUG62/SCJCz6t
SiuqRbl4kPi0l1OvuPbA/ipzt4tPhhoQ6icFj+5mEbixuioVsPA0lcDdbbScupzINaXNuEIhF45V
+vieJleoy89j4o28AI+o1WYgweX4dVoflb2LuwCO23MmiCa/S1NxoMQDzrSZ6kCymooNqbpdNwLj
7Iumc0/pnW/RY6N5wNNorDa2nNRB9IYj8Dp3Xh/x+UbwwV01ZY/DLnjE0F0dwtaSwqTIEZuyG+rr
PoqWCMRrgLfITp6UI5v7kOHON6Jg3hVjgJ4mg7vo2SsXmQ3PJ3UsGkqdijJS0pX3hr6+Ws88zCq9
TyFfUVrdFTqNObaEruRh6pUXfitwf32C4OSimBHwR/8/hwvtUkraTHE6euoZ2PGb4bqebbOmQ8N1
xvJppV6TL3CPuzJokjBfAdZSZ0xlolJmcjcB7ip6KGUQmm3nex3+XDSnw/l0YkRRyl7T2Ghv6vFa
P24IFzU1Falqg1pHFiFFefWuOT+xadlkswpmZMe0RpfPnSIzSZ0qCAQrP8Rm22eT8wcdHFr4TNMt
3J1Nh4WfBu8nlCaXoCGU4QDqmd3ObNfyE7UywR/r6Y+qF5a8Dd4l3PycW+emEmCmclN8VsvyV8a9
PUaMMyocqXeT6QIIWRR0Ft+7jrYtl1idItqQic2U8NyfpFX0S3WYFCFNd2SY0bsocJgd+4y25Bdr
98mWCmO+4TTGvfUi3BclcPHZOYPM3bfUY0DSPzGWZi2y/ngLZgb9b1js+MKc3RqS/A9m/xjRfKnl
M5U6QvwmVbh1sHt7n9AEnRjcqE1Hi0KRYcvMIs3ubEtOAS9iCeEnfwt8AS1AgHAAENRUICVoSPjR
AjhROn77ENGG4TaWbXSSFY+3L4Sf7yuZxvsvSSHp+ff+xWorAOuHLH3t8Q3k7IpTlR9e2ZrFEjp5
UBCC3UQSU9qwD6EB+6AiqAC1vkWzwzGcX9J6P4k0827iCTU2EEulPlGhIjKBX1E+6d1jh7vto7ol
wsTEAkZLAiVUx0ey1l6/VQed1y2qVf8rjp6fZyuA06GHf2GZcT149yilt3fJMU6Mkpv+rUqE1UxR
IkqxhEQ+Q/CEhQ6tvIcYhPv0wVcmeKbEAkPAWnCr6Sa/0K8jr5Zw4WBcWPeVfSlTiOXev7oSIC1c
kFmUo28Zr40+ssE94QXlHKHKF3ib1COs8D5ACmVLvmSpbcMAZytVMm61Kcin1G+Qjae/lEhfiZNO
e+MdpG8xEj2yGetxrUVK6zzTy0vOt4kx+J+g0NvRxZMZeacXSn8WV1UXH5/fa7J/5c1zTEcYZuHP
kE3iEHWAFTs5WraXWrHzKgukGkZHhdZaeG6f4dfplvBxUrTdUGTR43KNn72tKXCBtLSfLJTz26LN
NpNpcV559JPSYrkCE4CfP49CL/wzwfPkH0PULv2cIuC/RKgbTe/O+X+EzgvS0opUXf2V9fJsD+ik
QRDFscxxqM9zRAX+Hr77c+wlmakuAmM6wGi/1yzEVkgHspmTMoA9Uj0u6VdRSM5R+aCoNudC/cbh
kNDPfTr8/9AttixxpOhxPxAoOJ9eQ7RxTMXDy+S6QXqLttL3Ks0zAO6TrdiByCZAgxXqD6V3EaBB
U/YP4zmFIJWuKv5zXeHf0vLkrNApDaP0h2isyQQFQe8FZFvRvFYOy6rvKco/wJWElYPY3R7QGrj0
vEn4oUvZcGyce54mpK5IbpWigSrMA7ns9ebhiyIuOp9TT4N5sEnmCchg2NlAAmoX4ax0Ro83ShtG
zc0DasQR3s5ugTsWdiuSXZ9TuX1ckdi3ak6OJ2d/j94M7R6xU3X4ZoxTvWK7qlrD/hhyKXScuVe9
Ay+anEUfpo6W1zIjzoXLOv4WGcqIAvzH6jH/XSZNLQnijG5UPPGfqrKxX4V8h8neVw5WpeSSJYGt
m3/T1egKgvYWjHlhFTzps0WANn5Xj20uaVunmEWLfs29Uvh0tPICMUmN5gaN4YpgmZz7ZJSSJQzY
glf8tz4zmCipZohy89sL72dd/ROFixxzmw/NgVEQEEC7qrzmdmu4skCRGxq7T7hT+DiUh09WqPLs
U+vORM3PCZY7vAcjouE0kuKg5Z8rl2jXVZX0bxWq5Jjy9lSHVn9YgyJXkgEmFV6QCdvC/omQo8md
kX7V0HWa0dL7+Gsq8x2sKUT/KP7BN7+Rx4zITUyTeA7233TwNV1y5anqRZsXVtme84Y00/wTi0me
k2Te8/C7fLFpUsGDiCgKttms9qI1k2SjhQh+mxVUEFq8St+8bfv0rJcOYRfOvKJCe0UaKWpUvw9L
qxUQK4yA3VDDFci+T4ED08uGeImbRrfaRsyjn+68KND8LZkTTzgiXPxYDEaM+uiMS9lk8QW2ZKaQ
6CcrlPe94GXJ76Hr4OKY15zzt0ZWRzEx7E93L1mphvi0zWa+TbDRHfrs4HlqQJ0sIj2ZQIsv7riW
Yza7ihCTdahKIvoMIgXeP/stwmazi23UhB4r93FLXPLN8UJvKh3G2DCh0MiHpBmSHMNR7s6IpVou
1jUuDUkhOGDL/EnemQavAA5HHgfvWKSK0cO45VVVvqL+4CaI3c5QaGXjW86E5uqrMEpwpR7/ryAZ
GwWURxvKHfAR/bJbMIst1n1egRTZVcNTr/dFykYEI4DNTyjmx62BBNg9Xq0sVL5y4Sb0/BzJciM6
iHtR2uxsEyRFmbN2be2iN4KMu3R+5/KplX+lYLyXx6eGUxtV5Hx61upMErWuAUcMFLmz4ovlbpyT
F5tmgNxrwI9Kie1fHtI2hhQeWm/bYxyYHPTIT3s2WcqK4hXOGaQ7BKJjKFFN/57gqETKAnhiJUkB
9WngUY3I9HY5P8nR47vTT8gQ68ZYoxXlZrWtqWG1lMQ8kvyKX8/Jm5r8uPET5Z0N9ubWtG1w3iIe
RqFkIehVk7J67Omyi3Of/TtrD7+PTsIibXJ9RYDb3GqTDKSRam4WGWoMUMU5yPKvtsR8ipc4UP9c
vF0VoXIWNzWMFEbksZywjW9Py3Aoa3qeE4tKuUnIEaOb1igYWpj9arbhAtubefYRYKbbhnpaim4z
BqAledlti8vaeJ26HF1tJiet22IS7J7ZziO90Z2sWdhsjcAnDeyc9efHDsPeYB8gofQWbEhTTNsd
3NwC/74Owaw2PsaNgLSyux4llg0tTAiOmdlwpRD4dv6ttI026daJF/CKZqSXeqmn63YJo3SpH2bJ
hB5TqsOzYMZjWPjdPXIiKZ+S+p0FBvqO3C/1CdE2TMnKCkjGWzY/6ezMkP5zgYeiLgcvetfCBNBU
UgUBZlH942oqcZyAtks4s1RHMWN4pArO9h690ZegZRtbV1yQRpaRsjzM9vbd4BuYHZxEd8CyAN/E
Ng3iAB9Q3V8yY29z6/N5cYoKvdSBFn66ajchQ4rOKZb1CM6oYX0vB04I4h8mT78MMscJXk2Jyx18
oIsgXlehOy9i35DII69hFE2MENMeyd3JJoRt63ZY2AL91hBRu29CoyYWvKOmGttPZixNfkt1k4QC
BDAzsgiV8QigojDd0qea/qf86d5Wuoi4t0JCqTwN/YklRt/IAdIK1cxTw6dbKg48rnviE7qvLxfo
rZAsDrF/C4JYA5vOx5beNQEmkDsgvfckArdw9Ua8a465jXGkOJOEHogDFbRwmF+IbmrueiGPNnPG
6idrXCNchIQip6uAgqxHuKRCgVBEZ4Pff69ng2mLEjQh/Pd50L7xtiZ952VYlEUzKt7h9836M6So
56RINKcjRCevz4/3n/9rEFEXcnaWealLdTacWLesGyC6EPgp6OkhFJyt2LNFXklLfjf41xDYXIfh
MggmlByjmXFOinCEzBhSRTLOafzZWaeI4vw9eMAxKAEt4zqLT/FcqcLB9x/I3AHIjbrTvgxKIEvc
UJgfRwE4sohdp8IOzsTOIcLjbZSIPRFnzgad88aUWqZjqzrvNLvoOBsFttgh0WDRec83NvAl7BB2
I8L/2Q6S09hIsThDOfIQXlHRVoZdtx0mtHYrbvyH/cVZUJLTygKEcbtshItcG0YlcZPl2czAzkKP
nQZs2YAxhs2iaaJ55ksx4c757mKafMzJ5Ngsqkyi/kdYkk/h50Lap/3pra3ay307de21jl4rJjPz
dvOYC0L+FujQdMCwmgvSnLCWDl5sGYqEslxiSwi8IER0QNvaTa4mxVoD68mD9zJqRee6l6rUWmX3
9ugdXmsooYNWJ24CMy8LHwMuz2DS/aOZgB1DChiCGIQu5JANA+UU5kPdMvLH6r8oCbN9yNH4RWzq
bhq4JpS2KcA2UaEGd16DzhvsWurlg9E4qvE9nuIDqmTB3oBdEJmSY/Qvjn92C0fFrxLlKtHX876C
mmQ7RkSzCFqSga/r7qcPTJsm5/zbEVHoneubTsbM7sdFeD3xFRAKxw1/INs+c898ydva0DyabiBT
r1V2aAcqFopjXAjFGhHvJrZBC4hT7AjwUFVoaNet1dD3miZfNgLHJeG5g76kVXGOhRgE6XS7Yl0B
0z7ZImWumw7epFli4hZCNs2M3vBw4hDDLZ58HfzBmy/QKN9qTedM/al/P+nwB0BxY7TWd9TuMJis
69BToxsgG2DgBPYPi2M3JJYFN4YhCXS65PxdqSxpFu2X6OOcRXb19Y4JV2R4rlikRvR1jsefwwXF
OWSIXsGZ90C4KE2RFxzUTmnGHjcnjttwHCLcWpvqT87f5cyXPTHeJH8ax6dqVPnZ5OUjRCqBbINd
7mrn2KbKpX1EZWTQN1GXThfRopcmOgUcRiWq/IYrd2L37QHhRFUPj1vqUDfIYWDIXoEm9yBjxMGn
lc/6vh7voEDYtMSar/qAksteM0vMcNfc8b3e8sDnYxKl/BFAYkrN+zyEPNr9kHhty1FIwSlmpf0s
AKAYDYbyh4RDUP0jMtWQVz0JYeOC+gkzPbtmyVoiqirq3OUX0wgDjq5yi8QRBtMiZqY9ashsdQyU
0ap1g6i6RzcWWgvBO98H60EDJCcVF+cHfVJgpcHjW35s/5C2s3QgNZvqJiBvHJheKvyBwcKskiTY
OAFpbar8+52lFpfiy4DZVEAORLuK5vFTJD1kcq2KrZKDglxQquPCPnJjlGkE+CnKsoDBX762iiFf
F8ucp4cfdysqHQO4ZZQeFlX3RP+DOC/iV//YAUNUbDcBZBdd3XyF1B7+1fivsumpjKYA2SB33KRN
05Z98ZBnUiXjS6gkZW5rnJGuGcDKLsnbNpNRg0KqQOAcyI28hawAFryhBF5tjEqDT8Isgx9BYy1g
N1/QHVDtJVe7KyE97rpmuVt/xZ1wvxwyfj9ERV/VKrlSE9lRjs0681HnlbvFRijVBq+j7Xs+ZzyA
EQDBsdhyLD/WCjg3n/tB/K7gSYfUg0Oq7mn7eDSk4WTY7f4/2agl5C7gUQMkTFbNlQVAPIdUqlbV
xky7Bb3MUGrgPNXIY7txuUJ5kwGbemY4AN98k6JrNUknvSWTaN4ydhuYDPv1DvQdl2+ighrzPwfE
ktBw4cV3JdZecundTRX5DQcfMlRnfalMBH3UAzGVF9Z7pcXru1vq7YkvrTurfZX1GXR9GqAapHW+
94pHtpTTCt5hOR+pn0BoaarHbULebp93XMg9WCropiJoED66T3TATtibdbV3t7fwJWc7ZF2pfFV1
Y+W7RXYLyDg8oVp31cxmdNotZptV3Ui/P7RLRXR74FCIKb8Cu3mglO5J7u9UNvaCIBzYXyZ0vyVt
CSgmt5aBtlbtrN/K5bD3r6UBEvnDmZwpsJhImDZTv8R3yzjbot+fMsAM3qV4RP+FK9wYSLclFn5D
qvjwmaDSEXhFc2NlfWk2IhAWHMc4HhrGExGXE/lmdIVC51mCTyq7aod+hx2MIgK7nezMm/a97miD
5AL3yAKtjLg3bFKzcbrMRio6UdgTS/yrHRDuFKns7iIOvLVK69ppEsfI72DDOBG5XhEbXPpCvAey
+TB2ArbRzxo1bW6eJXSTHo7Bw/B0q79wgKdJkRIGkDNhuBLrwgvaQzJxh33hlQVvvcbiLQ3LMFz6
scSQ9RiifGO7bQZD1jFm0jSgvOKP2W0byvx5AIIyedHNgAKAXAL5duWdQmLHSI7rD1yfuetr01eX
zqunPuJjSm3Jx1F+kTsETxgLWeBaD3c8YxlqpRo50a5h/em7bapfY/xHKGGWje7ykJQitu+fECIK
juzkC3PWcu/1NhHZJswOva0G3wfLol+3qjELHv2ZR+6bpBuL1ytekdTAgZ0XgkG2ilyju15K6ST2
7xLxDxRhzRmbPxrHLyiZWicfpNj1xhWJe4SomLmqwmIcz31FpY526mnU9o3ylv5X9TtOgHRbOen8
szlvX+U6gpuiz0TXjxmj+HboI3i74Bb1BptARyeYQjXtK4lXLU/Fu0MA3A3lYXvS/sGVgPPmO5HX
HnZMIi3KffvCtqoEm4pLjgUlzyDAWNSzb3sEbKURK384dz11WMtmnhg/BK0ErIwWPBb7+hZUcv9n
wM7LBbgzCjqxO8u1SOFa7fgk7/wzgo31X84jx8BGVjgv/Wh/Pb5QB/dSG5X7CwzhTCygNcqvqpLy
TAMATfsrw8CEwWwFoxYHOKvkdVD6WkMBFRo4wbaoiXsnQReS5bGYgQ5k7LUQO4zHcStlAfL6qlJh
2WVJocHup5uUUod5Cf1HwnKAh2CEP+SlmYP39u/9S7hDSpU+P/odtYRUf8fvImRsvA4WMevuGfM8
1j+rthldyd0I/ZDueK5yVflP/ABTV1TwGDw2SqTBeSdRzfG4tLWjZ2XL+h510cPhoxSV5F2XcF8R
xVC9ctn8aEUCo0exFDkao6txiuQqH4eRngD0y2NzEvuc0tJ9AiOa4H8QUNXFy4G5jfpD+sax6jIN
gQVDyIycnPck4stdOM0C94r1bsfXywtzHe2ahzDWxSBzhXhernGQzGjLd8ZUwnO10iydjveWDT7P
FkpAtSxXbjIV/jI+P9ySjETdKCJjGzzpyhI0tfSSNt15CSOYFkSy6l5hiOvpk89icn+UxgeZpfjF
2zeLkTnNwzmb9/yV2f8SKGAGWN7QM4e97o/LmLFrct1AO3Lg4UtP+tBCldGvs7g53e0pUZ5rDM+G
/d9ZAVLeo6hYcgNBfTxlkfzg1UdVkxlyicIhj4yhDaBtVhhHGE1XrtWzIoTXQ9BTjvALK3XNO1ix
NpttzbuHGrX6gpwtXFDx941mUcy+hY1Zm9JRjbxhC6hEXXtR/Sljo+tk9WDagyyZYbqMQLWt0DHo
gU2M+IFf3BhEc76uQ6tiVavxySSZU1e+qhbWn9XHnaulv633Pf4P7cZEF+PsSYr1LiiQVuONJrkB
U2vM4T+xGbX7X/f+DjITexW7FyLciX+mpY4HNOWPTW6xgyyF4ig1AifXe02ptwIPUqDxzFAQUFs/
u2Bpsww/f1RM5dvLeJQPDQKE3Vx5kYTtroIq1bEHkbRxT66Tw3ALkj+vl3DN+eNGOQNzowPZP6A9
7FJRdbRzmuKlItsg/IAM8FhEwdijRJ7TC0Mcl9hueFb+o1u28mn0idTFLnQW1YxM/6VxjkD+WJhP
rn/cWUIi0fPnuWHkxb2LC5Yrj99j/Ezgj+6OmYEyHqbzsGgEE5uj1/qu6xI9Y3LIIwPDvmx7RL22
EuGzDaGeDZ9L7QOfiKlnYBli4jDTGuW2LyzDWqo7vo+dNmYwmCp6ZTuTAjMWyxWd9c/4qErpRrha
Styeqegs1i4PR8NAFj7zXNpBoXFQsVT5QYgjvo+M8TF2emvl2zFEtXAuwZfeJF2DUKyWiz5qK+Mq
FfCVdhPmqzOu1wXqFzHKv+iXPeueGCG+nNl6ZlzgjI+3ddEokxpZplIevuHNv/ofSEtOTqz4Ji8P
NyZz8C+PagBoK+UjJkeUV4ziSIvM+0OHah+xMOYlJEHNYuod3IupPVtJ6xAs2ge+uXVGloeJLKs5
11UVfRSNpTaqnNXXXGBLXjdzFLBX9YlXyVEAy8EJPc4eTWFpAygMInTow6LvBWGBILQbhreS881U
Kib8YE2OpeOqelzb6HBSv/3FdOLwgCRn7lOzD5nZX6wKOb3Puv7nIjXmLKITbYk2QP3xJcu+TUks
0J4Erm7WlwdnxzPx5sr0tj1sxt4NPC20gQI21Znx4LoHgBtIXGihGTzdd48W+8zdT3UueV07F/vA
Vitc4xeVeeZuYTSvXecZa5LSn5XLJFkTjCZ6BGG7I/YJw7yMHDXDr0/c2KYxMucrakxUbbQQiUac
YXT0udud5DnhFAskR/U8DaERgcIKZ7yd7zs08cpAMwH1usRkBmLuPMPyLqVS5Mh1I+1q+qW0rJtC
n2E6JjR6e3a1SxYWOuDQmB3RcTYksdTSCLxqdvjJ/zIIK5CiXFN9EJYtzCz+4A1/7Uch76tb4OnX
Y0+b/oaDDK9KqC7yXBUZzzzK/nnau/x0VQhCRjpVKQ/yWCe9jXYF5yF5rKj9BfvFafvF07/CTW68
/g8ukayxF+xIkTcOmOvulJ8SHbzylSzUPQpko8XS04Cw1lcNygQM6/5/nglnbElDDgs4rXXFds23
5y+ZOuFAZzArUYp+G7YUrO0wwPb+xcx0qrl2bwHGwgD0TB4MkxRnxotacodWeOQy/50O3CyUEwW5
TqBN5rlsMffsiFdlx7gKiO+mKgHzlOtDq7eZIruHBjp4ok3rU86SOF4rIREeYQG35Yue4UGRhOWb
0DOvhY0anlUS9qD/C+t9GgfPH4tennMQiAPPgI9JBlqQRZitL1rjZUYt5TbJEq7KRSDlq5qO1ABj
WHkqalqOF87ldbGiFd3EOS+L/dku6R8GgNQOnkn2Q8oML4przAPWlskUlC6Xd7fxKs7tgOQLi75L
NC6ZmURz98cWZXJkYXmA4HiY9ynDhjgf78/G3dEsHKQ56zgzMFf5cFAKjUxVIWVBvg1q+V2LDYvq
aQ0LxjUfagN7Ghq2CQApqv+2XLkYCoqN1dxnRXNaQaIaM9ZdKA59WxCnNQNnGHFcAdF+nvrlS4TS
lexmjRzCX2Cti05UNYEt5jPJ22CuPAmX676F+jnKaFTzGrnESKNVu7z+heIY9T4pLnMjWjC/fu84
0/CaWZ7KxZgrhuWOecU1uLPhisBVlVmS1jgAB8nMDOM/b9063NW+elyGTHmmy3LcBq2Y46breRuo
gOlfcyrMlL7B0r6NFstpoH2qREonbQI0F1OvXREzUt2bDewk+wzkJiTJG2CjYheWko5KX79qbz95
ZYvzHEvD/rT6IwHiruaMoaNSSNoZqHpeeRdFEXhHUkTubtloR5hxpw6jtqJuc0OdZfBOBVd3+Xwz
MzlOmPKug1J+yxZu2i5YfTr/2DkwUA3A9TGkV6AZBayJVCLL9TTfdo76i8GzBie/NBiaKQTQz3aW
mT+R1tw9ooSKku9lecvs9S9afJercAwO1nGnz8zgFTPnbl8bDOY1W7uTU6cbwpGuSCwwtIKFQkLj
8Oq/xzK904Mwr1f/q9BTwvWEA6XLMG5sO6m7gCD+tM3muBanTB/QG1slpPc0ThaiGHjXVEkUYVFn
CJb3+hHLSKrodzhYbi63kvD7bQJtLi1yLZcBVYkkitbwVVGhYbvsJ5EMahiX8jf2338UJK9/59It
8Ns/6EEIxvXzVqRTeCkhmQTULHSSaV9l69tFMoqcHCJbkVVKzrtRRSvvNkyNLXkeNroAB/RIdacc
f3Ij9Tc87NB8Gg6zs8YhIcaJp/UJ9eKLV/kmgaTu0mO+AQSF0YTDaWbeoCi1cTSM7qogSEf4cxeL
pZOBhAu/27QYFi/g2TEVZOOFRD/CqSjcjgdlQddd6UkUpmIn35TvL2/oDSVs8/KqKRuM0UJcob1/
XdF/i8+VR0A8wRMqzbumXiYl1cHErxDDlYTXtROjmRTjWeA+DQYUNQyiJ1bqJkPpmejWJ6NGktOZ
g7tVTB1SNlvt3VXybWH+mMpEhD8LS3+Fa90zp0CwUaqyWcICyjtV2OKuMy4Lq8Qlxr7RSCppeEfD
vUXYnU+j4BGvbp64jQ1BYYEY2unT4WVMqRKpx5t63yT9514CpPrDoqhmYyHsbSAf62mcnnnwpXqr
1JKxuSi3hg0yfoFku31zBk1QT6Ce2iQ5I9mPkVc69mllrWeWpD72dw8EUECFCVe9vxpxtP7tskSJ
ZGKITepBa9TG1MLXtMSnG69YGmKGe9ZEQ9OVu9AKT62SBgNDAfMqHGkCvZHulxjgLFE4wnV1+Zv5
dGY+FH0i2Pb8bTG0KTn0GS2VfnKju00bv0JVKSP65Q3idTTVryfA3tzz+eJqnwoRLCiwgMqLZ7xW
zrm414RDPCzSuQbuggnrMsKaXmBzEEnAUbawczir4fCNEoi8JhPakLhdoebvHnfrYrinbzOWN/Uw
wSlgymJnoNGMaSJLGlr+8NkNepp0tC7AinTvg6t8OYrduxbY6QI2pvhl8+DXzoZYXUnVEIEop0Zd
5kHn9onBoWIU80fZeBQ1v9Kldlf9KpkOO8k34KhpRDxFA0wBqs63KRj56b3XV/NQojQdSETHBrNj
lysM0nErahXAqzcl4VitnmfXzOcs43XJs6CreOGSh6GKneNE3uVR4kRIsOcEnknmDSHOg354vPnM
8EqC9czcqiR9jCDYLzCX36zHVBw/uepboo1bl6XzgIyVG744Xa7lfxdv7IF9CYFLyXEWUZ1f/6db
/bCpJBCIq4RFU/i0/f9v7x2FRmtxzQeO6zn2K2KV1YTbORIn1KdR0ddiZkNwmqAPg+AkZuVk7B9Y
xTlpup4/D4C6IWsi8T1TVZuvDkmyVARjys9Kr6/jvP1/8lDtx5MEmOASsBK3SW5agChqZUYdXAo9
8xOx9N6IIxCY2K1Y4iJ2yumPlXxoNI1QfAZ1S4m8t6na6V8fnlMvxSEGGxEBUShT0wwqegdMiPLp
BX/WuWGZAZ9Bmk1j+NFDUCqWwGPaOAr5iwGyxi7Kv99sTSa7f+Rouh+pRXybMdpbqOK0NV/yNc7V
NUtkfewhEa6tNtexXEwUPMGp6dlJqMIhPPtEBccg+Loi4k3V4NDJg0LlutfmBOZTBkJZ2CqTC+Qe
Igg5CNrayxuDhXWCFgz0xZNyf9PnQ+6QqCm1jv3mMqSVUAjmH4RD3ype7D5FDfBNUvEF1Xjk7AkP
NCDygusCqusL+huUI8NJ5YERVfgWBEkILjEL8uWUhOIBuyrLW33ZrBT2X0fZBjTEHp99UYtaHKqE
RGVMKOaRlgXEXoeXw30cNZHwujG8q3QbmpCSjtkjA1OhsaLztizGHqjWzV1PDFOpwfNAKqa2qdGT
v4IwJaz8x4zUpMW7sgqhRoOFmL23wHMMUG2Ovvgj+/My9LvKtcTbO+BIxKxJzSuhqpXpRnYSPEwC
hTfMwd6a32orbblDdjs2nc72n8UqOlduCONa1a0uEq7qMCeAL6j2kkF+K4fq0x3MFdYwLttHdw4W
IkWzMaI+4oenOVYhd4NEfm0nTvQBH5Eilx0tpXGBAXZ//TrdUVNFpXsnMSFdWGS/kxg0RFaVfOtC
AACcb64kiXoIyvdNU8v7bLg0NERz7uhq8mcIsQSlIyz4HqaQ0ah2LpHn/v7pnU7je/r4lLMP/1EQ
uvB2Uf9+LekQtIEaSWI5tve5VkrIur2u1AwbHuM8J2qb2dwgI+EoG1gli0TS+5dDPSsIOTvE3iEN
juuxXE0JO9W/vFN2hf776wgf3Ra7RwIZbTpMNrpu1/1d3bds3zqPiGmPsfXUmooCo4ZaDuVi14Z7
lgg851/BkPyuXel5+Fyk3sOk8cAIn5/ntiy2jmasGQGrlQW7LTcmG6EsqhZfxFwjtDmOreABwhF5
Dz38xR1JM5PI38WKFjo0ZUkXdcCdaI8viwR+w/HHaUvdyTIJSI+XWpjQ+AXjgmO3uzK+6HlIWzsg
181KSA94zd0wsy+ZjQYDthSIR6aCL03S4t7JbU5QpvJHJr44zK/p2CngElSVWuSSmGjEZrTuS5fU
x6WKiC+zL/qnkFkBEcVxtfyK5jeBqnEHzATCpvblnwv+ltYwgcQqrxLQJojNXcRiswD/WBGj0qyg
IRYihwZEtQ/EpEQKQ8k0c2vqAkJAYVnr6C6VkHfepKvT/amglT77mNTicK1yEG7HR37Rgd1qIHo3
VG4A7moafhIiNH6I+ZvigsLpiJSgXpRYmfIbCP3uWkydDq8dKd6cWu4mX0hWDlZW5op/DD8o+uGz
iIm8T9LVwVSKtroMUXiu332TkfFwl/ydh2HkMZiMRMpcI9TSythFu/U/bubRyvgQsfIHZF51Z9Ai
pzR940GrX/zFeKkq4zdvRkRpxbZXB7HdTCTmJ5WxSw7sJbU/ciVfmBT0a96+NIJHJDsWj400PLU6
Jv2tY9j19laCy6rQYzxTCkndnYRo0Drmdx65rpvG5lnd/b28dmFerOS5T0REwF5tcZ1YuN/hOneW
3u0bIz14xVQZbVUrv+p60CZKNkmUHIwE1Qpb0357S1RKjUNwIRhNXU7ZxL1z3JLoXFd3sPF+OWRK
6VFM07aVxdVj1QH03I+ZNCxeaVVIWVkpbNgkEMY1cGqLtNVVyl0Suc1hnfdlme2Ahyv3grjQk3BR
ORWWeKLEB07TSAYVxUarodJAqZUPKEPuCugh/z3hVw4kTct1BKCg8HMY4Mxu26pcJm1epJoDVN4Y
nBb8MAr2YTTXRTqvpEG1VF+NzV5E3+Q5jVN4R157sqeQMrvAmHRe1t1XiG3llb917BoYnkc6Tt4Q
XIY1dRzfevGBTj6Xoxc7xfMAt1075FcKwL0XSGssPbf44/7o+RrVGx74KhHV1BD9gGqckXPIIE+L
NZ4aJJ2W0mSz+lEWknFyTCLjb7Jq+MeKkxg+cXPvDH8QwLdaxUUthp8Uhmc6NwRSTpm4mmdEHgrE
ffD1s5tArYCWfkAUvdUXQda1jQKcX9rpD1gr8dKFkDrgHUHZhcEddCJIxvYnt25dYDOZN64bjnaf
wTvnAwKy+rADc5hdD8wLZKFbWNjwAW62S4R5BsoqLXhx7Yc+5L3m+D3rdTd51wgu/cXP9wA5qCRd
Nc/bQRXNBwR3MLghzGsiqTo4atxIVEWSUMSvGd+jFsYC1GGZq8jxDFmbWuy986kYoPXesa1yJvxp
aUSkQUkTvtVXLlFnmjMJHdk6ucBBmT5kaQerEKJm9RAXmxYQ6bkFGDoW423iLtuZA71ssBGIm+u1
jTALCapPvDQpMjcJYv/rkAmWN1bef+8Bscwq5LiO1/zu8mCjy4nIZmdmoUaeC0jVikJwzE/5xSBt
igzji9BUWK9VzsWCJcjAo7BV02nxzGHESxL3/qYWnmeBCSw2KxxDjFmdwm9KXH/hObkLHEEfZPii
aDx46nq1VdalIPkJujzys2rQu31mSl2H++/3UFMlJQHRu/lGhCXRL9k7z7bKDHasT4Oflq8BBc8D
cNRKI3lAF9yRWlHUECpKhCi7dYkQ4SXldZYkon4wM38Jcm5NQC9A2d2CGfoGr8y0cw57en0B3wi4
573spqMcUCbcw+KgHGupibhLZ26wF3hd21XYx3s3Q0wT2LEuOIW8b9aif7O2Vpf8W0wBbrQvep2Q
1u/l2Q+E/xrwFGYLsXpV1bXGgdRI/7Cc03dJ4DSdyFLgmZ0mkVeJOPh0bLysQU9Jmr2W6Fml/HjT
7BpToZbsJUudwI8ulQqSZ7tRRdCNmq4SElc2iyDfgMsXHkn1gVNmU/RUTCjprV82ZRa6SpLZer1c
3lbODfFwYvGbqC0F5XWcQCI2uUxg7x5RzyfHq1aEIYe0F7rM5lV6oPpwO0b7Z6ADivVKeKx4bENC
dsnxjLzkDADf0f+kaw3lHdajpBinZNngfTGifMRCvMA86j8jmnE4/ioTrs0JytuMbYEzknQMKa8w
rUkjsPSQv1QpKuxLfZxgCiP61d77ynlx8QSDL+TplaRjNWOCYbuaquGGCrPeXlgtU5VluTmAcG5g
72H0tzYHsS6pPuBzceuyoDxO4I2DohmQZeS7YqWnd+qIN+S0z9MT480pz9dVfVnnpgYEUV/iSna6
G9o9Gsxp0UMQhGqm8pT2ubuTeNtga7/Cof36znrRsVzcpurGp0YE2VB6/dAot9a90IluuQ/Fsv+W
bGnjGPrGpU4HkadSd86v4glL8c2fZdO23e1bui+zIilzGt9M7aYC5SjRXJJCSbymKX3/KEvEloMI
JNygPHDBU2rHo4E5ZcF3rEw//JwukXkkeGK0cDqw/FEP51mqufGRVvSBEWTtPUDvvsdDjshU4kEA
4rCa5w3HRJ3gG3D6embIY7q5musLQW7hCvLKipEubPfSl6aFhRV7pqLMqBRtuxW7wIdj9f1BCkk7
5Nd6XtUMayV88Xn2BG4yKf7olHGR+i9fvX8Sn1VKd0dr4AU5oK0/YbirBY6Iw8k+jqweZ+y2Y0/c
Rci326YpgPj4435/cfVtbvN2jqNvxsr6mucbW9jEKWJVuCqliuqBFW+YdtJR9BI5I+1iqqoeK25b
gaXa5DrbYEm0xidQJf6oqROmm6aafh1IwsgpGiEe5Pksnip43ugyWuO+gIdj9rmM6xGqmT6bDj6f
/QqZpeaLwhLcQmOP2dzPo0kg3lS1cjYcLLiIPMbmjufwGQ/AXLGBFtSKvLe5xQRRmodDnmGpIBQ6
KJgEniK+C6yAccwLaPdYr8wkEgdHWQWpyIUj15ctUWa0/r0DIcUdagvl6BLDSiuG0OT52E2F27yX
dWhXEDjL51/GQJJD3HDbzCoUe1+ZH9kNxbvHgy9cF6FpcIM6OxcCkfOc9WtRl7WV7r6DhxibohXs
qwoPG4LPSWotS49YdzAf0nmz/RtybXPO4XB4dQt7cBGyFisZto9YEehTTlD0MEUp0W7BQXwAjYwW
/7rjaq9GmGwoduSortolNE/Nd6MKReLdaibFFmOHdR6aI6b835m5EXg+p2kSALQP1ssdB9UYXoCG
BeVlCDqfk6WBa10/rir9qwbnHab7UTKA7y2iW9sEApHL4cEIq6ZXvqa6dKwbbIJCXS9MGcB6QSsJ
S1WxdOwJvjmXL2CcC6KoL9ZrieYK1Wk3kXMMMm2a5FHm5fhsAWNO6xLHLfWFYJgwmDXmG2O2ns1G
/ezUuoc9ELymkfBPbx8PozkvAoI4nkD4dR33bXpS8cY1Z6yYY0U5zmQ/8SlqyW+LPU010mWMdhsy
uF1yR1RQnu8wsM7H1ivpOTOprTSS7gmnXoWI3dcTXbguCdcUwAwHIbjWQAd+f3t3nL2QAkSS0FFv
5JoGZ80m6nPuIWa/FC7GkhY7TBfXzAkSGlfumELypKgFLD9tXpggXsBtutCT+CJKz0EskhP4vt5V
HELB7hp3CCiv7CP+qO1mc+z4OjemMLNEFkIcgnclRaRjCiqJvpfOGYM8soSo+DFINPli+/gKSfIF
uKeg6/t6bcKu9jsgOc72WZ7IILZYoJpLBP+sCHYpri/Gf+/uBFt0AgS6kDTId6pYF+3hcZioMjhr
rG7DLTQeRc/0cCXCEdLug2eusGrFH1b+CzUq/tUKsOQfMFueXI+0xP1XoF5hD8OsTG1w/COrwArB
mFE6+b39KOAcAci9q3MbLp70hr+n6NLBNaAHBrJqY3uHgx14JMSq15WggzdAzDE0PARWIJZZs2TV
tNQq0nw3sm+UnaF6FmFxsTRAIfz2IZuqo89kSg41SbDVQMWW56soo7PNomSjDPeVn5mFSytxMmLg
Rd7cHt9Zao5x/0sqP0k2ufcGl4VKsocdbrnIJ0iPFzRDprslntAGeZM2iWd0Uwip0bXcLsoRhr+y
njunL3GR0/toLEwsHFTIxlTLOqUi4l0fvpwaCd6F8UJBx2RCJlJMLAo3oNWX3cATTG627h5ZtaYV
KgMLjkUxCo+DCFay08VJTUX786VEv95uJZJZ0ckRymYhUfK+MR06KdqNg3TVA4LqF9Z/y4GeEere
txzvSF/utEqEa6ZG8s93MOmk3Xl/M8h4oXXF/ioRybHRwQPtBJBbDnVjbVOBV0FXCSYXlhItBIcj
HfNmIruHINXbQN7CJqqzHX4LmWrkwQE6d/zjulKKH4IWp/rWWVx58p9Zb0dvCvskGZZgVMl+x7QV
vu2hhSXCTZJC0axTmYxxoiE+/EWiqsSx2DFjj5/oZHJX0p90HaPP58S0Yr15YsNMoepCIbXDpsGo
o3gb+tu1Ib1nIWfr0KR3nR6cMNd8JmKrDM3BDYzg54lrXZhap38lFBK+A92+wUNiA/Y+XT85U2rV
8aJ3bgv85GniV1sexePRMW7r2h3DKE9V0dg+PH9EbYntpI4+ZVAmUm9HRfwKJsXusK8LsOwUKbUq
cA81jKLhzU8POVpDWB/jx4LCdGWXq6a2Z/BNmXh14QXyQ/QsoATNKjUNrl4t6mXzjZFBiN7WIcdO
tOCx/kvfoyDs7Z0HU0uMPxUM3/y1+64+a6lfNW8WosM03S+/1HPrQ632p/n5Wb7KCHBO/u6IQz2E
EAjbB/raw+C17DV+VwhXgB5TmNq+Qid6YOWEfFr+XZIFIY9oWwz9HWDLepPYCaN8z0m1Y0LCH0oZ
i+mONKgLojuVyyJkO/6jhmgcZlz7oWaP99kNdveRCmg3nteQEFkqlUyzaG0vfEZRTcpMKVYE1X2D
EPLmQgu4EN9jZblLgE7ipvC5cS7uE+GmxGHb9bBn36cWsV0q+1tolvLShLa2Iyc39+4bPP13z1yH
Auim7ale8JpqRQzBIx6FO+gsqM+Yd3EerKy08iHfWYvTfstFbb2wamBrX59cdam0KRpyS/eCfU8V
5H+zjD8heqduqURwMAEL1I2m6LSjDpYAsmFeJaL1rtkKs//9nQPPWbr9lXdgLZH5LoRLFTnd/JOe
Z4wioXN3vGXN6EcCF5a7i2VSoIERU0Tm0+ZDaEN/y/BCj7zNTeRvLtm5UOFE2v7rdF92tb1+gViZ
MHfPsce8mpjOHUuomBQF6EJB4dFq72v3ev4cuh2fvUEWXYR6pmttuYV6fdc2CDn7c9OPUTof6jJn
Qu4PlOY8iAdAMaI5Dvq66yZ+HmSD8wJHpPAf8lBz5u/yIzLokhDevkr3gEBjQimalKI2QDzc8brJ
o8sdC2lEu0GDAg/OedJZ+wAN+BUzFTlwmODJ3/7kcpE2GoroGPZkaWANKgw5aaLPkOzTo/GCs5rK
J3zgkNdyDuid7LiTvBVSyDLqB3LDQTfROEW+F9+HcvzMZGOluh/v+J+vLsJCLcZL96VQ7ZBN3aNQ
5Ayl6ndtdvk1rLPzcRSY4c8qSn1eSY9AhCRU2fN8rnJ2xJo0yT1NnmSULC7cW2+2UGdhAdBz/mvn
qiiqoMo8EnJnKlxI5pg6giF4lNYLTaTMVRqcjlBt6xIa49Suq/agb7XpylKfxvXbWNyicwOZx47T
SRmOvi6L/uPZc7Ic6S0MnzcW12xFEAxuk53glqOZobDHpwZL1ZquUjMofqKEElBmu9Wq5CkEGAyg
iKV6r1MfAOkKnPrPtYzkRcGjXd10g9qI4W8muit/+IiyPebNPdrUg1JmoRoNWD/uiijYkbbbzkAn
q+65YjDQT0aqe9zaK548Kpy0kIxHWmCBTxdsDvwiX3ILPAQ7yohVBGj9UPPrpQnivuXgKZr+twl6
ou5YxEVPJyEmWuyKVj1hk4j02M8EQUlV4smp1zT8n4SKlXX8peSbfkZ1SxGjdT9VnBv4yPuA3SoB
59QnOmCFu7td+b9Kqmkh0cgwlm0VC6Vjyj6V0N7kDTTJvjGP9DCF95+iw1R9UjkvIQFErJXJCUOJ
QZhtE0QSGyFHDSxGi+uH2otOFY93BG0tpRQmkWsGXchGHSTTYdVvnl7U02jW9LUoBhLxQOAh0tbL
b34zJ5JZPXmvBh061lJIvfjV5plJTYt7gzOKN2/OoWseXXJieM5ukKbu1Q5lYKn6MwzQ9uSinG/0
1FW7AjDLYMeOs8kyMZmg0MKTLhWmEDm0XehXzf1TXNqbFUpFL7Ryl+ardmIE5hv6NCgGmt4V6d/I
P60bAn0FdaOJq9uki4Sul5fA/ma+0Loy2/LEhRIeEZ9cgxsz+qi3jxf+6CLiSmdnAej64hYMlG0E
WIt5+cbOWtULc9MiRF50A2V9M1ynYu+4OZzTEBtLMj7EeUsNcd+HCh1+JOXKsjZq0Vpe53juCRuk
xVgTFIE27uQKQCq5cm6IBNx5LLcA5Ku3UAXmqisQ132JsWWst2VI3FpFKcbG/jbi+q/xUe6em5n7
eRtfKR92YLqSULy/K7DSAchfSeO52j25ghrM4686ga7T/GFnNGGjjplN1S6LwGhMStiMUpzSGi+V
7cvZbZd9rn6jzfCy77mUFdQZv70QC0pKCKPROWiCnZFFvVhgrlRrOUbcwGXMis2hlj2d7DQ444f/
ik2UjO/dHr+GhHS7oDAEkL4VVaBMy5Gy5NjcIYJcUvB1EqkQZyoIAlfuiyLtzkdmX6B7WdIabcAi
jr2rLfSRGQ9/BTaaXUC2RQgorKVQwdxwaKv1mKinmkBtCPMXV5NtgxTrGfjJ20SHj9Hrhxtg+ql+
6ZzeDG45mpY2Vwp2Szt8Dy2AXPeMs4gk2pgYl9a10Y7gjd+G89RKJ3NqlGfD+lwW5ZIUvk09TztH
xQA665Mv7+JkHBtrG8svGjH1em1TOAIQfNkzpo8blVrdFmIUoooguFZXi+WGl3/1g2L8HzxtnBpz
KfWqYuMTr4s42WsCV/qyERdQHnBdUq6UbF9JiAn1flu1xrWSeJql0b7Exbu9i40lprzN3YnTDP9M
KkcIrD4k1U4aNsYfiSwp76hRv5dutTFK8ZdzThSWAE2+aYFyVMCOS1w/S7rNeWBpxa1fvmBHT+TG
GWqlFJFNSw8ElhVYGgkogcPf1Q6CQDPVOVgwnP3iD77Kdzrplg/NLo4LHo95Cnm3wiltMBTwcn7B
WEtGAxL1JxQsPWS2atFo7quMaKc5fjnEMcCqigKFYq5wzw3Y5E68wmqKIzXn1XePHy3eC9S7tqnS
o+KerpOHWWgcL/JSu8nbyVm6wNA1icBcQfh3xi/iNjNmTdbi1yNb3qMVIs3LV2Q+XTmMKZKoCEsS
xCP5skplzrvJERoDkNO0qnnGoRVdS2lCaN42VuKUOERmuNKtDz2Es2peOLp6p6oXgd2EA0IMv4mF
CYl65kTbbK1vaUyxUjvmsCt5tL7lLInDb5QZpOR29PZ+A7EWBkLFTIkhzl2XZe6mksKfgbW1ngyg
6WdGQ57XALVkMC6OL4SH/ObvhEKC4plNdYZd0nyltALZMVR0i+rKzNsrZZ8SBKJCUbOV1+DSuqG2
dzSmqlGn/hEBWy29kV4/CANyGuqC9gfPsxlHR/CSLTsbrJUapK4TYPCuG6+khjdxnRDL0YB1MUFr
7UuUt+qXEz+lml4yPyNgReCrglUhmYDdx7IJ41C7KlPFyoQUFdADuyaAmMeSQuzQcOisYngFdSwD
KDVdXGNxSdInHXY8ehn2TpfGIbDXYqN92tbav8EMNokpy4Lwc9PHSAYagfSVQ3W15uymudxGI57m
RSjAn9xzfV41DHl2/5l3ccfnrn3g0Bx1z7JMOVjpUYY9wCdmLMXMpCrKT6lsSYtt4NGuMjy7b1zD
VTCAzQjZRuBZBNgT9aEffYQfmq0sZkjzcBEhQ5mio7FIMe7MdqigDy0f9fintKn97AC2NhWEBVwM
0HIZPwWV56B071k3LSo2WPEWcyOCLchfEB3lvzSCsY7PsgA3YoGRcyYESAAVqSM1Fpq8kIviVLcx
ykHrddO3APxJJq0Is8DrYqu/F7hS2FepDDs8nKoxrK0n5i6u4Rh6VFMsm4HyooL4rTGFf3OCj4ud
ZvykqWuN22x5CUQujiAQQkgmH9VWeIACqWMKThBlkPcVMxjLXjv10UmUCzpMZScKjG9JWLdaGYmE
4k+kj3MNS5xPeLV7GIKaBf3pOTo3ox+e+bZiTscjGCn9SqV3/h125QVaL5FWt/vFVU9bTgdEo1z2
vWQU6X1lFoUt8ty3u/r6wnhtQxOyaYUofPI59/WhH3lJJ/14G5k3BNNdvQKjoB0q0qmU7AIBYruK
4qeT3dhVkBH6q02u+8qUtKcycuBIphltZ0o9ltCYgdZ/z3wUprum4XH2pOCErRUd4j2Udy9POZby
CSnw89+gDo6kt8xwUqPreUiYOQMduRAnNgTtXFZV+ihnpEDXipdOyctRi1FuK5dszP13LSrbCEEN
i0K2y4Nf+kXSIvbRbUfjRx/u6ZMLY4FJlbPfEu0YsfJnVoBM+1EJ+SFoiuw5stlJxD2yHq4X1YCM
vlcouf28LiXyTAmLOVgfVV9aYfSuc5WIsxKLWFMi6u9xLrPkgoYkZEB7KCjaHjoIGxzDluRod2FP
sCfQLEVgPxOs3KYT51OQybdT9pbXFT2ON7ru9yyiGU+8MenGZp7UIMyQB53nNZkvj2yTEDFIZA4/
AUg/ysHS+E1lizyX4tg88QBl74Tm2I1Q20dVAZWEocf3ie5MXEQGOw6EaKt6SAdstYIANZ2lBTAw
EXQuE/sqwtYkaw2m39E4nGuHDhCheQAQMEiIlcYUgpDRUJ0Vm+NhmewSuM0JsgZPwJv0sA+DLT8Z
+HgK2XDOGB0b/BQpz4/omknOQXA+nDhL23Qw+jfdZRUPjNagvwAoSxLdEnZArYTVqBEcuAMfFhT3
KCQs4/6BfKGl01MYhHKZ8ILBy8x4/Jh39dBzrpZLzaH7izXuPstLmDYcBOPVQufvOGzZVPssAIOm
x0566fWRUQi/OrspeaAFWu2MMjpvAS+Y0kanVz8qbdBYIK+JBbv1NrvM50ypAZugBjz7EwbrJ+5u
A4llPHbzkKrlnzzpnshvQ7kqiyS1caCMuSIoqCQWejPWGZriL7k/sg4/zOibYqU5cE3fUczwbYyA
kw4KOYavOox9MlI8DNa7XRXlUvMKwiIGMxurxkxqUjNRt54C70DS1uaU46w7O/vSuEc9ENRunA5G
9GbgUKg+EpUCcYEfpKb6XhQ2U98HwxcPudMUoTnySpeRQwIjEpav90yKhBx5QasfFoYd57wk5MQv
ZhdzW+XYFQxBRpahCRivULCzwgtvtsXm4uVWy9KiPkG41/O/X853Rilx6dDm8LdXtkTa/27+bFcj
BZM1bzhHA6A4BDK4wLHp7PT7vSgouKARP09Ua9VswVEtccQ2Ey/smt6DIw4wxhUGSooa2c7GTDlG
UjSUXg2qPeyE638eOXfOOEMWwYMpMwzAQGMGlVN7o3ypWqHnvOrDBNE6mO0f6eJQ6MCP3crOwMoq
9Ch+uQPq+YvN5Fv9w5+EdFeNnPux57lWyZwe52M16vg4Yh7ZvamotnKWW7glX/Txax5V7Shhvzfn
Yn1G2xnibWCN1cL/J4/eCiqBVviJUvBQVsVusVknijW1K7x/LVDtPDW6sZiCtd+sJJafq7FJkBrV
lWzmCPDZC+WV1AIU/kb6EGFT+4QmDToSD05VaVlt8SondJLNyfW5ITlCOumwTsSOeElqQ+EJvfDO
wuK4DDQ3iuh8imOqPfQAixtoZ8Gf1DXAfCtD7oYlQXslC+/pZ5pDQ3zebuT07c2vt0mR+fM02kpX
f6YrHn+cJRq99FmRUxrzYZypdsT6VvszeiP7eOtj5qWfJXAWIvLZ+ckUdvBP3q3I/GuQXCpRenKC
7pQAgbIfxmY/rcJJ+mV3vijv5GAQrhMu/0R5gummqBfI3HuOAH04AgFqCKgw0TU5KmQjmVw6OvdB
0uXBq7qpNojfLTaL2gH7eOCvTSOl+wgPIrw3NDubgRigxjwNd2eZQwOOafbKXrUbDwfrd/NdDosb
IL5d178F1wUNgsQn2d4aCtns6RD3CgYEV1vZtTBYqws9mqoboSRIK4KKskSN2eF5uTPvhC0nORlB
n5gNVcexcocznq0P9zc1l5t929aqsI+8C99Rwq+u0MbOSWzsxwGAIfoBxj+2s7g/hCliN+I/llOY
W69EgRYTuk8dLXJrYMNd2fxJ2JEzGB38iQdcNTav0QIOF5auKV1VSx5B5x/QK1i69wFQnAUU1g8b
HFVffSqDDCce+FoDfOf7V5ptLamCAuO/23PIdvclb0MyfSHXXzMmtPSeXk9ypnq3sQLNhB0KZUow
nll61bxHmOCZuWwaRtu+zHKnQwPMP3UuReQE1SZ/nsIDYzmspQzjc1e/oQ46Q98NaP37FtLe0GUY
lt5EQUd3JFxMdH4aZ/L7gDnHK5wzfiDMd5xqeB71nMzyPuasUxJvUNHmO9oSd712qoLZFBWqbAdV
a396nQSyR5+TXFTuM36LgwjCqGH8aSoVGZh6ld0+eczlK9FRpCD59yCyfk0U4qcbZWVYV98WNsOb
TqwsCyEHaMG5063zm3yELkQCq3BLCfCevFHAECjiWVja2xvMFp/CeKFG+PDEVt/8qvEk+qM+w8G0
DKWUSlKaAtUPYcKKJcZFh9PmbzJHh3XIlU8TWB6XpSazvg9jOz7+VghD4k0dEK+ptoG0gFw/kRjs
aZmRDznuGffMCmausjds/HzIYAKTBmkGzDBRu0RvrsNrz5nEFWLkLKS4jk04klITPhPVKWugTfT4
IwsppCnTPgp9j/Of4P3/+ZvH4lxHdCNQBS3I6Vw1kY7BE3mb2MVt10rmzjnCtxXBljVHsA7wZ1f1
A7gjsxkkHbTh66P447D0WfAKTa/nr7b99gjrK2dKYt1xija6WtDyTyWGG+vE4eWFWQgff3PyDS+5
vQG1MrSKDeMKgidbwXqkrHuYIlChmZLJqpoRoCXdXdWXrUQbsaroXsjI83UoqVo/lvVs0jkXEeia
0OKHbcBU0u1jiA9prfTmDFLHpN18pRPymNJZma4DUhWzIfNZURJrhPzzR9e5Ax1JtUakuBXmSS54
gzqqh8KT9j/THHss2JTV1CsBF7qt6G9EC72w9WBEIrBrFe9XN5ooIJ+32Ur3qySPC6+Wp/HAxVNu
v4afjw15lieCYDb2/4mLdYfW5u4hIZdTYKwxcI6c0HBlt3TWsg0T+7ZMj35EtFDlcftUWAXKeLPR
z3Wq2mgxnLOQIJJ3MZC10OZVel3/9M2UvqTMQtwn9oafsdZZeIMjLpL0bem0Y40E76/dtwKA3TfD
cx4yY11jp6PKvlt8sehaSoBRuL8Yfag+PEJkF8XKs+ZyCcnsUjoN6tGHfXRkn4FB8ywaQTGVVZxG
vp6LS4Y+C/VgwiooFnsbRk0aiENWQdKgC3v7iVpBP26rHtr71GGSmSFjNrWlSqMC5MX12c93RGEa
62fDegBPSAHhH+CcyE4Q4MDrwkXnZe+pHo/4rrlCafbYi5gLm+mGoDOlqWuUt0NLQ3LFyoI0jwp9
KkQ4ZXsxUglOJR8mM9IrGEBV3cL04H77X2oEU2Sao6nWOV+kYzjS2g0Ri3NWzgoCI+ldEjhz2Zqw
CgZaXuSAsyff0OcqQTFGNmQfC+oF/k2wyKoPdLMzRfsvQ2W/fW4f1wRVSMBtYZijcPVkdUXcN/qX
gl2cm2pdOpkEPDimhCZrZkmPxFsOizpD4zJFokQknVIubI8PdRbcuSXik6u1YZYdSP+FmaJ5uDOt
fyP1UuYloZS3XFlEv5CgpOETqUDBeE4zKPTxfKwigFa7gm9IdLqTLgk3YEVx4TNqt+m6/S23+Aok
zxEqcjQ1X5h7yeqBBw62Uo+jhGq8ZGQmiwQ7m/KjBLW1m6EccHfGHPkFbHyP92m+prqkXrEPpoBq
SH9Ccx3NfnbNjrBzaRmnRvLryhQ7Ks3MvsS8OSpbqDJXCKueW2u5hI797mc9qsv82BgwncjUAhzq
TGvFBbX8VeZ1GnA9Rzuef7EHw5hO1XUGAv7XBbtSdghONAT9MTwf9R/wS1erLFZX+g5C50EP3aYZ
FOdmXIX4CqW55C2+HavWUFpKmOYK07PoadNUnbPrIdbxg3Au2gEwNkZoqMWLGWtj7H40aDF3xNo5
a+3yrg47W8RzdBiJjreLd6/MEGsz0AZ96jFiuSPlbi+QV155TpRK8Y9SsP78tE8hMIton6LQ5KmA
330ynxCnUXxIBAC82M69Aezvjd9xyCOV7KyjlknVPkJgVvTzHptZRWYB9gaGJ5XLglE1G/vuj/rW
aP3Ee+ODXwkvskToof4FWKMMxerKs9iU8k8xGWzFWLyjopZwCLXlG7VgSvTF93IVjtBpHJ8BwDyf
REOl2ZJGEWXK+tqOGcDBAIBccji6WT1suWRj9Q81fxVlMWMgDEjHXnKnyM3kvCqqDTMp4C5PYMRd
1WNefRk4U+jAg54H1iSiYHwBDeXkkD5XAc/0qWCWVMidIiKaPitRLDaG8SPAmGCNZLJbJoLwkSz6
1LfINSciVWHD3nVw1YxrAK38hOnRXS8lZ0M05m6siMoKyltoiKyW0Mv3lKRWUd7HGUpquFzxbRsR
VXuyjhxXhiKQAUREiHfQC+nPVRPBI3yFzPgWxQCuorL/NKp6Z2BXkUaT3BqNfqrxT57hK94tocBD
pM4ygl/tovDt2ikJl9DmBfiDZy0hpgTvQW7CaTsepIYq+pwKUrDWOs+qNdnjFpNQEu0RLUuir74T
6WMjgd1FxewwFHpHh8n3aFyHca6suYxE5LSaJHivmORcoLwbgI2JyHlpjEOUFFTJc0mInGM+IXXc
k8OdU0z0/wdpWPDNVslARmKogZm/Z0IK0D/1OcNYf1u04igQ5s0VxNVPfUJ11jVMCJ/DF3h8V2LE
MtZdcIboERDt9SvBNYsBia8VgHmZJd/8SQhu796CQoe4r0/QJ3AOnwwhbRq82yjCdze7NHCpyRU4
4YfEtXSU5Wrd+5E5qHPHT3tBRb0OfBataiJj29L6/3OcXtOWxx8j4SzGPmzITUJ8DRJ91ZkI5XeL
g9boWMWlSnwVDZEOZFjk7Nkdq2pt/837F1EovuJl1FrsNElGbVGUexHXOqimZaTIUcP3Bo9ulQIR
4460P3qmn3J1rZJS4hnjt4UkwFHph5hFEaDmJsG3wUeYmSjJWKYfwUZPJvCkJ5AOstyErWgX1dcZ
4yyEQMplX+gadpyb9wDNTIF0DtXWRGYUnv4HNsG5iVE1zJ+H8wgEak6mYkfZ5dIwv5E0IltUd8Op
e9Rfn1W45ZRRfT8UU0xfBf7l4+GOzbgCqMId1M+IUcIMnH+7NdK7iguPo4dm8Z69ykpAWQ2MBAuL
gtkBx9Igo7A8fE9dK5JL6Y1BNGB072Fvg+anljbPK6qLttVuzz8Oz4rhDUK80BSK1QzO4oNJeTQ6
wAr+ECptSKqHO03/WF6IA/VITVMLUkyyeF+yDndQ9eBD2cNgiLCxt7vyI8L2hHj6R18fzDXHowlM
IfmqZUGfZhQg3sTyFlAi6oYRNHqFjqjvP6NM9Po5MaO3dXIM8kK18r44j+qF1qzrMj9/zvA68JVn
wKC3TenL2seqWnS3nDbaV/rn6z+9GpXk0Rt2AFzB0ASAkD0Z0hs07pqhR1JjN6QxRhjhujWCM/Tw
UV6shHpRUf8dMTk1wUpk9THhmCFvNpYA5BFF04dNG0NiWVzO/2QBuOAnNih5mgaObUYMNwaZmmkg
4zezIU+Onll+LTXhDLWZI82KuOXCOTQBS/fwk7JRKJapztcfOPUdIVSEi1eUHOhRiyokEwQGshvz
eVdBm7OeXI01DxICNu2GRAhAHIqtDkx/QEKBYSfBe5SHBn84uHGw9nhuhvNfA+Qgkimo9sFWCIIJ
+BMkbkL9d93BRNvq7hyFbrBb8of6S6/ioUYgoc5tSxLapbyr0NejXfuyPVJUfhfGV0ai3AA50a/s
hxDjwWZ/gpge7ik9uBivECMf+1NHlBqmqoETHfGV3YVFof1gzv5DB2jV3HieRV2rVzh1uFSnHnuL
GfUe4ICrPqE9lE6r+4CMXBHEMUTkzhK634w+A3x56CVHE04Ck1XMmb9u3whR1zxDp2v6LwSnJ4IW
t3jQCpENSlb8pAEuBSR4IJj8GjJ+Sll2Y3CvjKaUT90v8RJyGiovgl3WzezF9wdEEwVZK223Iaod
5UhVglCjF+YuJQxOqdj2x69N1vbtgnxVxi6wAaSaXAF0kLroeKX44p+qtMEPFZwjAXBnwpbjDYwk
XstIPEgBXqmNhbohIFcAIwXgkl+AQG+stVjp3mIZvIhIHp7+zU9vfG5k+I+RSjIXPJMzHjGMezpB
VgWfCLYt7K74N7GBotQ5Wegc8Yxf6u2uCDg6QkR/RIe/EItt69J6/ECVPqLw5/cUE9Kotj0d2xFJ
AQjHRNsF4adP9MGDAdyp6rkuh5pm4NtYKpHGckGiMOyh0mlrM7abDgov/QUNOnT43N5LFCpHdCw7
2PE1Z6DKAhA9eFYY4UacdP/zwio9cEo5SgwLv+a4lc+SptnRI4PUQnn4zSwkPD2HJoG+oc8vECA7
YG2JA0KRkD0e1wvGYCFYnXILgfiiDUbaZebbCrTu08j8s8l9/tgk3/OH1BNdSurDG/qrE7btQeE+
d80C6pxxHzuC9I5fZef3vNXTQWugn34deUSPPhbOiGnqAs1VSj79lZrGhfAnIrdQpzGvwCD2eKE2
UGarKT2wfMfmyN50OJyu4S5KSk+CDJvl8+shNEBAgQ4I7KnQyErgn9qt+gcSY1VICwcR690a6KOE
pa9uT1H5eeDnCgSDq6OZdsE26DskZLXg7MktBvvtGz1MOOMJjKn+zeK0e9PhT5qDYTOUxD0meyQE
m/bZzDgzlp0+GYokk8rZjjlR2cL7RVWNLBY2/puQmyZ2zbmkB0cJ35bO0qpi7vYqS+DVgiGCAvYQ
VQGvkzaMRuC3sZ44tqkfZes7FYWlkit/0v/vL+szcSit8e+mGvs7Ndp+WCZsuvaquVGnncRjnDzZ
tscuE6xfZI7VuQzjkM8bm1O9zTSRwCCInI6jXKWUxwW/MTpKOGLURu4PB0SFLYunYhp0IY1xD+S2
Aw6WHyXJJBJ7aneia6RIgvC/6T8va6eF2yfvI03wrrO0XNBU9tpCm5BZHFW2opTk7IDP+f0cH7bY
2mWdzNp400MHuXEaeBqUIp3cB5QBPUZ5DglLqhxG8kxHGU3UNUxxyHSO4p35engrycHF90s6/BKs
xoZPanqBS2/drqL5pwtQW+DS2bpHM32V2APocpj7ud90QKk8d+ml1lrwvJkBk2Z9vPN021h/GML8
C8vLBoKi/VzXl3JCUC53mLgyna69ZTcBnAcOHN1nX7ODzCT2N2I0u6/+XZVl+PjpcAK+/yd9lxvo
406Txxy2mQ4h/uY1vQuUt1Z9An2jKhkDGCV6B4KOzLsVnqs7rzCc91/sKEdvs6Q+x/3JvdeI0WeK
59vWEWPiXwD8OtPHf0UVAiVGxAIZXgeL5FcjGFc9MmPHTMfmhrQUvgBYNYdPz0YaO+KhDuqwlUtm
H17dZm/o1cAv/415xOF8pNVaKOhiTIUoPGDWLQ/0idXWtdp56+Sm60S6t/xuu8ByDctHBtHWAZBo
5DeEd1BffWenikxefuUQoVSQAg7XMVyWGhWgfQTa235IXwc/G+hjEEv9I4lWP9JvyBgwqWzCjJij
BM/zWkkOC9L+zQMWV4AL+oi1u5CsTyUZ+FR+TzXEXSWTRyiOP8nudEjJnAjs6TxMDckCXW9+MGPt
p6Gigp02ohCk9MNnQPUZzEXGtLztXd6skpcClsiphJkakAq7tGA4XVZbtmPdaFkz3/TK7ZXrViwZ
aV72ojJE85c6ta7ug3CXRwve4KmKcnue2sP3nVcvHUaVWVEfIN7zwLQ17wCp8tvD++OVsNwcl/NH
SYJOf4eK73XnI3VFwSaDwW8E6e/j3sL3undwyvm8gRvw/fRarX8Yn0GIFz2Vt1q5xa0T+IG0TunG
FLPmTYrSebjP8S5AbBLrLDdaRUnrc0MVTMFf4FQQydTWlMTN0RXYRHcpuoAqaJ9oFHehpJyK8sq7
Zg5vY5lsXp0LudaHmWqlwZR5dT9QNRERAaoWuwlEXnUF1hSzq/m/wZ3xKSJxXbQK1Pf7Ftn7NhEV
PO/5hJCXwavo/ky5rzcEf1eShc3sJcpu1ch/P4Wc+Fvp024G3oI+ybh7AcB0DWKHDT44D3oitzdF
DArFZYUvQtcSam1PHPtGPIi7YYHaDogl6VMrJ6MYVlZde3czT2laB3kXKn+WHgrSr3AwmgYsVXTu
riTx5aek/pKjZlv9CWVO/n2GXuXV+gmyLgaR8JZHq2jEZ6x/KT0RTs46sRGN5mneTnmky6t1vj1i
BM2zGWe/qrz1DDwbID6w8YZMw8IbuNzdMKMqV4mJt/QPbV8qh7NX9uCZDK0YVUPH4HikeurJxV5D
MaurMEdIvxDh88TKFl33GYhYrhgUc/cNzZ0WbODZyFgqw6q05qFUDOKbdxZbTyTAscFUMH6sq9dp
TXrsI0J2DNXwb9Umw8WqAJ40hoaIaHwcu8mqZ/VZme/WJ5j/uGEqdwleDFBr8rBgl5QcUwdhaLfH
1C7iH7cNGgdJH4ky1ChTiCL6sCEyUtraovQjN7crOfYb4paJfQAO4Xt9kKuDIlgoyDUl4Kyjln3u
kwyh08I6Rvt0ONLWI+Hs5tXYcsJhxTExMv8ZfBVlKI0UklbOJZqzA2LbfpI7bhmw6P/E+yhuqc9W
EU5yJpu3shKMmchO5vsWen7KRc6kWVQJhu1jYcuqjLoY4MPtPEe8luB9C5wEOB22uSEQdSXzwn3H
zOyFZXGJWo5YdCRgRlnWjYnmS1QnZd05OTuueoPcfQHUEYLQgYvPmhAvwXnjiWt5Uftmw2+gi7YY
qsV2eYqKR7295L9O0FiBz+BFPZS3T34vikwCfyAAj8k30TvCtxBwAItSiFpzz/27haUy3Nx1IrBs
sMhK0JIi5+0NiryLcohWUXQOHP9Tofa/uCqMsqQ9cIwh1GRLzXsb7s1oopjHyY5WKcC0Ct1/IUnr
r5tyxKmt79xsHempAQjk8KYRuek4QgU1XvyT5DsL1UgaIcqSCK3Pbwfh+fG1kedvzF6gr0tdMIKK
3UwphIDPbH70a7sOs28RrJqaaW0653RfRDBEiULiGT5vhsrm662KC1Xh56WE5XxpRl5uMJbdCZer
0BOhhzYPzU5xqSgfqIOKQ8EqHYvvNHcW+n/zzKMG788Tdg8v3P6GrtMGVxNH4awS9gLmf8ScntP+
TD+hUMuRhKClrPvPG1Hs/z6opPt8iw0JTeYpajunusGC02TS/TWzFAND+0eMdrBRKqSilLszYpjY
rsa4OhcXbK8m7Sa/Rb8J+a1JoJXyjt0lrltFQG9R7EyNrbNfCuet4A+1gHt5IUTOrZ8sdmL0FcJP
yM6+2oZECg1/Z3WGXI8bl0fSHfKhpJXdTJjjtM2gNxBMuXMULVMb1FqqpGx+IAws7+2a7iddMnpj
iYvUorERe+CogqF1JDCF+mYrM1EWevOxafkKnoQTMNp+GUIl6ijLBXPJHWwKFXsFilvGpCluE7GP
t/mo0lu/w2eRoZ0+iD7wEvxf1W/hovQ/Dyd0kgdR6NAhhIsxtgiBtEwM5TKIUAeXTspp/NUwtpJ8
dx/SojiQ0bSjZVo5kgtYrWvsl7jpSmoxnod3YFET/0fPsxpVDOOGDff+VPVqtAskho4VzkAK2aT8
TJiEb5sxVa6NQAfMg88bZgVcQagWoQgQHSLor9LK7FeKHtB5F2RbpULu+piu1wTuusfxHuY+eWoN
mwwalfKt14wZUb4YCJLlo0iFyiHLbZIkGdHr8Qz108rYo68yprGFYEP6iaoeWv31/olCAmR8IiL2
q+5RbiiXIDp95eIIIF/Mf3VQ4PzZrAzrtSYUVvRwB9tYTB7SomtVY7xPD6LWB9//ERB+mUXib1oE
d/uM2wt7tX2lxUT4o+LIla2RdH9ji0BlYaVVX5HOTEhydAzqBkkTp91ol2udh2j+sywcS05D19/G
z/1dIrmdfkuCu6hC9RyB9ACqgmwHpJnKqXNeD8Ia+vniHxvGgo3mX3f1ed8OGtkE7VtL60igWcuN
D0UbKQJO9JhC15VFpq5Md5rG1pr6iWVy5uL8ljZSMinn/Z4j5WrpjRuDXMfBJssHgHwyzihvjs+3
GrISe6duxwNEGbG5dOGdMfk1CIF0lTrhhA0ZUDE8y5vjsE1aIntO/nOxjRa4fD1QByQu+PaCxWD7
WIA6ggzJ12NnCk6DNLSFvK0378Xtq54uxHHRA7YVV4XuON6dbU4JNUpF9J94HzcdreNuwNmkCmGR
4WGQrF5wgqCWyYmQ1F6u3a4sXn6DnoCNO0gc3+eh+cAFALwTyEAYx9BNsaknBz+ihlNpEwViVJ50
1sQrAQU1oQKv1o3Ne6pZ4NxYsmu0UA4Xm4WkF3bYDeS68AS5vVnHjzqYImMJttMaZD/Crprv4+f7
keN5G724ylRZKvQaq5AM82yMxhTOd0xiobIy/lNzjnHDrZ9nEjQwqrYtZRY3ttIEAxbbwL3rJofb
FcMnlkqlcjyGy7TY/vRAzJPcgXIoMF1ev1RnRLedGjmE3TvDBcbh1uSxjEFk2J2nx7XVvehP3to4
UeMuesGFv6WTcZGqsUqKYVmUXXkFUI17xa26UXdNrvLwzELbpPYuTIH7+ENgCbopmw2B5QOz+V5k
5921UiCgtoWRrOPqt061WFWe2mc4deACgO4MeB+UIWbzcf/FpvN474mIwfN+V52QKK6QxC0vt+p5
RIcijEwazQ0zCQfZAyKhUFtWEO0HG6ReSo/k7ksEakAoAtWJfJERPn2jUb5F/gx9gBuGkeaQ6M5T
FoJgXeukPueynGnD9qO/HHgv/ESpFHb3csoIinAYvgQGMsSG51vqsEouFIHlTZ4zn7yq201UegE3
fAvkb0sC9fDPYPkWajKiiW07qXJkacBAi0TjPrjsW382CBADc5G/lzqq0D8w1l4dFcnCHDpXG7DB
7crUbigw0O8ulYTmcT1qeQw0qqdHy/LTh5pMtbRBGrOJ/tixtCTXV8dvTR1ShkmV068fv6KGs2Bt
EDVqBvF9FuAD2R5BPadqEVo817CpapXqFKqBvjbTA3kokPhbc8mYGmcmaHa5CxR/ctlxxdGhFFPu
djnYVCL/XvYBFQUBHnGdfoasaGnlCbpx1mpq594mQFvGupP2VNDQWM5x/2Kj5LVZWS7OMDq45sr7
mEhNuQNjds55eNPCbak58HD9HxYG5ce4hiyjXoRPMJiQ745rBLtr+F0u48l3r3COlGtKbyQ/MMkf
8oNRKxviAPsrBZ5dJ9IURkChwp//UqzOr/1ek76izYX307zNSnUSQH3HpJZcRUmKy2u355LQ8O9H
C64zMNEKtp+WVkph98c/5F9RfJEy+IVwPe7OUguS4A+vJnCBwZV7jEr1EaTnfq0WqeI6uMQA/eq2
Wpy7d9uF3kDpfOYlxMYHkcPBQcEQIFqhy8HcuH73FR/uOpXD7d27Pvi7X5F3NMwZmZW84KHFiC6a
U+TUWHb3TA4s9yCJ3lPKiSIQeW7QNkthzHVyEvZFOLea/Zj97R6PLYaRgixPrXnWg9PUJjxDFk5s
55cFUy/kfWJj89wF9CVgON1AB7M0tbKTNjFP8jXHOkM528mJQvgLAKwzL4iOt+407nJ2SlaKhz/H
/rDYPT9rf616eqynTa5olXnUD2NwiqFS9ukGOceOP0hEEw3mbOjbZ4xMUy4FzQcwW3IG5I+l547x
ggz0IcWIB3DfXWfJv5yrCyb3+tYpJBmhj6m0n+n9pQ0bZ5qFO5s5ThXTEda4DmHnxdEWeb89Zg8X
q+WmGjKqyvbu3QbJ6/WqvZMoZ8iOUC85sK5uLqyS+WKB5M2lPzAYWZDcVMsbPcXZYJ7OSD2FLGLh
BWfbR6v4tGBQ40MpzWIO+OAbj5eZaIqRoOGkcCr418O0Ei4HY0LxLx9gZuKo+jhJYk0tXWnhbSzx
IwbUpgAOonMTL5m8VdKwblxEVlSzISShfOJGzuSWMAqDfTGb0yEE4EYkskl4oNUUVR+4QWC2M4Y0
RwQbIaxZnBFepgV4EGeioUpcETv97pp69odr8Sy+OwCGl6u0ogOdqDiixOa4fjdssSPrweHsIZAe
gKDoNvDGLfyjfyvuaDCofpeDFqTOhDy0/fiYAhVb7VIwusPvau1SMsK2vH9+8JKr6vvcHapssR1R
Ah9nI7bQEq944tQP0b2gFX2eLZNPvGeUv3V47uOzePe6hvBPRBgNBUta9IERSMHZDW3Zgr3HUu9H
i3F6hcx4IRn3mED/bq1JxTc0cNlpX0aVO+3eZpNSF2NspdJLt/cvZMsD7Y2+R+EuawJDbuCb63h4
GF0fjZIbRg0Y7Jr9VzGwJK1H6d+MPDDRL/1AolTlSsPpOwvCe4h1sQd1oxdktctAk+REEORsQrU3
Uk5IEoqZL9aJRQHrCxuz1SJAvCtJe/apjZvv0E2KeCp4NZcxjSB3y0TfTa8/GzZXrxIkNsXzMvrc
TiZncMWI9z6/pCWpbhM3beDp/zwGDeU8hux96vqXAVxls6v2QC/rKBMorwawPVXOVHnAibw6Eu3/
kcqkL9YbCx671z1embUisk8EgOHYbcSSmOpE8lEeQnPPT+5PZN4zJTXUjoj5P3BmRyxrev+j0JBZ
qvt279JStW4/j5hvi2/GHmILOPxcAOKWiEUBtgjZSoi3SKAQj6Tu3JDD0UCYz/w8tHpnH/vslXDR
1rZIJ6yyxYvJ/m0DTXJnYevdqomDSJbX8IF5y1b/pdJ2bmGPSD7kE9xtEoI26DWAkeCfOETF6V0s
/2t5FqM213sgKC/Q50Ij5H23W6h2htgNQDqsgrNchyjNx98sl1A72KERdJecxBN2VUrieCwWlnPZ
zJA7c2nvwobNe/kQKv1Tsw7CZtMNciRwha38/rxHDN/zn/KQGsMK2J1qdcWUt295Q8GobILCx87o
lEg+HOCK0YZCz24t+qNIxcVl5BSyYbSeHCR9R+tMNo95xqqrL6JtwfFKefNwY/JAUWCzhAWp0hXn
7tvtIQSLcqHJIL3NPE0FY1HegPGcbQway7quFnLsxFCU3xWCjwKHL5YzrzLCJtX6rAHbpKe2vCO4
YwmUOys1wsEHzNRsxPuyuw5cWsi11ei4DZ9cfzif3I0cwxL9tedUvLIV2Eoddqf6EB7izsd713OH
tUVKzdMRQB5Q85DmyYKH9CI390UR9EC+tgOCON520arT5sGVYGSdeaY/psSo35xctiyujeDClykk
Y8P+Xf+9ngDs5rFZjeA/b8wNmYGrpAk3elcLjVOV+v4BSlriWymderh2fHEHhdupvizzXfTxw7fK
q3lRvBegqsWbKMsOuwg52dGWQM6nio9UxLnrA8lqO+PgzYyoOI+cXvD/1+pSB0XbelR0uP4/7Dry
D9xOp2UMUVaH6tk0JjMcnQGlLJf81qgW38uqQVDEDWFCqf/67G3wicQuQyJUb9UJRP0cWg66IITJ
cn6KD9TGn97Xg7AiEXKNCmHwlRjfJqmI6gSQFA2dEEB0ADHoT+Xhj0G1TCvsRjz40CVAyJ4mUkIa
3av7geOqscpLNzU3Xot/DfuEYQ0jS+YHCWiC5RmdYIcdzbOI3LyoT7YRdvhK4psoPlD7dLFHh3Ql
FLxyGqZEc0VrOghHRV3G4RPbIT+LxHVvMC2JKjfieNVMi/e/zYmp1vcS7sFgtq18eGnXyrfXzfiz
P40RlXL3DPyN4Brqyx6wbg/ayu7W3qLyK541ezHkx443kd9wmymf/kL4+OMccZ6IytBB55KdbUL0
OHIlskhNYYJZQSoRDys42Ge3xP4TDcd80MMu/gNC3utTLoVxVxfCH55nu7I5P+2zC4xMchOln/YO
A+bmC5hBLbKcMOdOYW+WGIm6S0U75Wr4/7Dtv2GubtOusyzdw1jaqMoWznpTg6FoOBVC0LVNCtHv
SlChT5cdpQiMbLMd/IaBMLzoAibnDLHHY3goNhIUA/iZXRzgUtjy4Pxam3quAwHq4srmNrrdqV5M
t7wuaGE1ByB6+XH3ex14V68OUkLIG4NNt/K/M7XNHndL/4qk+bpqrKLG0jBI1dOLdpjRz9ltHUH2
3O+W2QJ8pmTNX8AW8CY2ob5oeuvMNIOie+8Cwtf3G+WssDkPJQDfo8R/uhG9nhT75/mwvuULAAP6
tVrstsA2FoLx/2bJmOkrI8hzyT1pN+h1eRBUg9R2qA4ENWFzdH5s9shqIVs2XRRLZfGug+uUrvJR
9IAlj8rZZiHq4dEF3hSR5+Quf+C/w1b6EfFxocReZfb9nAEHYKFWQYgK7/FswQX5xqPokX3JW/nk
Ou2ORbUzVsw5EZyje1NFiWyC1aIqGfpipt7SonqwKTU2TnR2W7QD+ejhqOKdAFr6T9hQC0x/gWLY
eYstBslJiO7pSQnKlz6gWFFXu66Wcu5ge34nJHjz9ZL/19HqotgEgGufLQcCahgbbJcJSh/a92wj
emiDR4hoEN2kC6WYw12jbPfLjI+WMs72ECNhJRceBCisfk+K5bjPyvs620fmzyE6ytOGC/o4YkE+
/FYNAZHsz5UuiTj0PNDkDj21KWYRagcmCwXxOog/g9WlafgPuWLWKk1vcfm5nwDsnjTEe4f2KX6b
gdIwx4ahckWRhU5PziwhGK1f5kpUBDosR8EsuH5ovGTFU65QR2KgWV2ILnhtSKzvF3fSJ1qDCyTn
1dDBJoMg25ifLLYfJSIfcpLk6p0oG8Jfbonknv3k1nJX9alVjdr4XX806Vw/eLwvHMXMYeUAgQ1s
ei3GxuAP9iks+rrzfvZeGVBoCznUT8qVJ6hQ95oTvh7/wb8hXZchHVSNdh2aUxnPbnB5CWGX/J3b
+Ekg6j5DwQWeDJG1z4LMQeH4USnL4fhXNTb2XdJbaESTzYImYbpJZhKEIFi1OROHaz/cpMtLoJwO
NwvcnW9kA6euX8JnKWkAH1nnJNr7/lNgmH7ZCHqFdYOg37GppGhRov6ZovpeDNht79rwpvQSeFoB
eRpQoN0ygZ3Bvnc70uLARkJoDDcwFtAt/2Uj3q/EkC1XHEFuILfdSuVL2498oFBX0TlY4c9VwOas
6wWWXMi8paoYk8FumT9TwcBl0Pvn87mU/HfHNS3AhC8/pWtyOomqzbKR5yf+gafTUdqSNaK3Ez+c
vpnxAFOFcA0/ZBbQTNXcstYQgo4gaxpkoFv7MIcfj7dWbzgx7RYa1kT+IECKc5fUI7+tQFDnbXcd
xHnWxY5s0vqvTXAuMVdFDJXe/KK4R8cHrdmxJ2soP11gGIrf59OtSo5PlXB4i9Y57B79pRJSY2ll
4xClwk/rmqyLACccJSUlWPrHQBV/F6GB9vuhJepvVL5ljCFI/LdWPyZuBnxBE7xWkE4fGL6zBUtM
PAgDN3zGWYv7PPQspfnqhnb4lH0FOhEOIk7QwY0/EUrFlOtLdiFd/FdsE7gRhRUx7gTZf7j4bnyA
nzdRAbabFQZDT+a9s8dDV1jdvOv1CT9E7F/6dZpNFlFcfeMMAfywrW2grTMfBKr1QvVmetVyDUlP
SY4JOTiih90LIrEb/A53ONye4xff8D5KY99x+UsJWynppPYItYxyLHsXl6pSl8bjJArpmTp2MeQf
UpljcdPgx8giCt5a4y1QLDaS3c5N9JsyAmBHDk00SJdNEN5tG7d6xS7oT+PyqYii4FqWT+WaxX3S
Nav9hcKLs7fl8KeGtT7ln7ZBXsk5APgesZTbcNRO2vJUcetcRb6nKmIVC7nUOvU1zew99q2dVITy
7la6QtyjW0zO1NsSb+WnSO1HlDAF4Tl9xfnLz3fTojGNaxQdno1RJHNZZOLWn/QTJ0W2buRwHsrf
y+N0hKw1wznG02eJi1KhY69dNgTEAcVfWIc3ClU+dmdgLBKbtKUQSkIzcJwXFex4bacyHYEHFUvX
Kzp4KcbtYEwZ2S21+SpfWw4ceKMwSid7eC0nKG8cS0Nfx2L47I+va+/2b4wZMJUHE4De5i3Z2GS4
aKQ93ubuVfsFlIyfEakSnxVUOizjvVPXnFcfVNCeTlYG7nsQKKz/3qkX7IoRaKvzJldaB2h0oPgj
PLjtamfoUsLPu/YNGYfy1ALBKjGquxVTxsVhD8hvPumbTChwPvT9wo/UemSPLwU1y0QK/G8hTJMo
x/OtVKtac0O6RRthb3aPj4GbK2B+pvsS7ZOs64VL2cWySCXyF+3E0lmzNMbVjaqVzI1T7Da1gMS/
+cTmuBjwCDMnsc92UGXlZRXQm5OvgClXagSmHvIVpqG1HJ632ZOPIzLms1vJrj1JFXQ0DY4wnKzO
b8ikLG62he7lfd2j0hyFcU1/NyNNp31WWmdZLvCFoEyoKMofKINYu8xomgzTOaAIYBZNFsZ8njn5
aAJkXYTa9I2h0IjS16fgvN1k3L05oC2uE1C72uto2OvPDYTyomT+Ru02ZrF7Lz1fgk3k+dsHj+FQ
FdQtQ/erJpJW8ar092bmJRHpvC0NmNnNbedR27/QGGXsRLit5gI1moNdrAWFIhBufrlEURsle+Aw
vOc7OLJLbsRYodIPxPzA0MWbby4MsVet0wnFG9k8yI6ahQVhhK16IQZtHXMem2CAyJMqg/VqHFDN
OiOGs68YQDSsW7G8lm89w5W/zv+JxnTmQDRo+/RwyryFqG7hMFueLXX8j9S+v788cEMWDiBzrx95
tNXaed1ArgB/SIB5Zlx0F81Y33IdEM3UNPXPtThSTRJkSk61dAmS1O4SEXDUcuBzf/RZWWOC4bKM
Gz1ny6/WYeKu8CH4XhjIs6ViOTbhDVxYU5lJXhXg7QM1zGjz0rwvlgPSOgg7Zia6GIb1aF1degTu
EM/iXme604NLSo3Qb2644ZF4VZMNf3H43tkutzu5NVHQ0ETX2g7VFlNRqrK3H2mkJU5PnseKoiN5
xEE6WZaZ9CS7WH7tQfXV3brZlID9rhdDDwmJhuMclX7zodXiDbyGuOEHtbc1gABSUY003oZpICAn
UsPZJsyoyQ/x5zR+bsokViFw1XMcEiY3zlhCwXchOC/MlrvTjDd6Rc1FPrSTtR6mRYqKB7F4sWTY
mVg/UaSEzOJU9/v0S9+iVunZMs4sgsCGDS29oDezluGnk7g6dsDo3TuT9kTbnttrxyyfbNMhfN0D
twlBmhp8OQwRFJssOhI49owtXm6UFsMGTKSqWqNF/3fajZzL1ah+dQ0BqWHTfQ5IZtFUE/zjPTfe
V7F8kWBO08YEHQ8cmJaLN8hYlCwzUxW5Lq/+b1SYn2XyYlS7W6gHBJbSgxt2yxlapFl9ZysyOhWS
Uf3krZsdt3LasbFa0bzQHCArKviypvYPawZkUrlYJGWviflnlrb8zczGSgOPDjg5ABv/sPIYQjKE
wLgY6JJTtRZ+FMg9WaaFHIcDPtcQkqsmMmylvFm18+PXYpIYMRv2ZgNrdCkN3scySgmWTUCXDM8Y
tzSgn3F7XzmjInUdUUELXXOhJOR0tbA3kUEfiGlhRc3aIeKZxr9QV21ndWmBYoUkpKvrGjqtznDS
nYh4eUTKq+sZtCzbXklk694uHeQjgtGHzb0T3uzt3//pEY6mv3osuzOivLN+VTT0o/wYhM5e+YSN
3yNkiAAlgVM6dG1aI/1GmRuH4VawSyso385PMyuzYpMg42u9fj01CEvO1rIJayWEGBM2hvsN2iIA
Rg8GKBFwEzuQr4dS4htwM778gzFBCoved5RP1OV/2Idb3xerWYiZeq0oZc8B9AByPPvvZIA6urdb
oducqAsIuc1lN4SDhQomC5hy+pJXTpL3UeyP1kxo55ZZKzZNZDJr86VNVrf8wrL6wDA7Pm40tWci
dDt3UhF5VuNWwtKJn6Vl5KP0mKI6X3u4nHzfccuZWMS7261dk6OjdBdj1IePWEmiBOl7xdUS6POr
z1TG/1XNR04kVmxHBnL/CglxQI7OU5s1XMrIKhrhW+ebIE74R+AfeIzM6/v4+rYNYgEMFz5og6/K
iSOxn3kgaQk/hkg/GDGOVQjANW3HQf9bpaeOCxU9wFoiEoaxYbJO6zMsccNUGMp3k6wJT5sT1hmg
infl+NUEw/TruG0QN5wITT3t6i5Ec0MR8cVv3bRzbxgIRH2TBdOBaVJW6yHOBLpXt1jlKb4qHLn6
50ggkpeJac82ErwMGWrOzrJJmGyjN2BnUfC0U0iklv83olpOxJEQ/lWZYoTRau1CZjfh03TDIbZc
15MX7Lm/pv+ifGLxAVAwjv93e21OpYobBDNpyJ8ca3OqHHgtc/d4jKShCxzGWbxlTORpo6zvnTuk
Vxg1AACq/iF+CD4OqFcNpTsr0nGinzqEoieKg6bwgQJ8eg4zrPLyq40OjzAH3YAjWUIxyePVL6rG
nCk4F4oq/jLGNZsB2XvQhEzGkTLSHeGtrorehyvhq7eoDEaJavVN8HIt8CWY+wl+sewNJOp0UyNd
0lBohJ0lNG9zm1jDTNmMGpQKL3irg3psiX07GnHQ3kAHC3hNP+vyJm2Gb8TbrSU+kHfr+uSBoeZV
0M5HYdy/hAFElN3eXzN+RRp4oJQpBlXEhOsQNT5LqtOdn8cB7XRaUqZ844k7ztL5XZpg2uNdWPYn
XrlTpnL39dVe5TyB7irasSditSNJtPG9VvpaZqyxIf5EgwvltjXByNYTANTdaCB+/9QFdae/1TrX
aWWvI0CA7lSFVHaEFU7b+0Usi70Qy0TUrUUrtwqjcZHK1c63lkl7XAgbf5F4rztLBhx1WHgjGWLW
QHfxE1S9yN/rI1RDIVleyQOdFb+rMtuz7YA1YlodsQwAjCOQGZ8krZkYzjoQdb5/2kH4PrI9Yy6l
cQ2Jr/jmO8CsrB6ZCxH3aTgkQk24wyObuos6dV8LcEg3FuMXsVmqg0tXZ/xV3kC8Y2O4IcD3ztf6
clmLJPMKuIRiTe0ditgw77KuFNTYVY5FRzopDm4yzwAzWAZTkE7UOTjbX16HtYtfdKYrBPnm1/zd
cHbgii6oVFFEsRjI7qvU6MWn87mM6CFy7t2xDcJoup0tiW3wE4arwzL2h8i+Bgw+/ZjXeiC1caST
x6OGuAc9Rh25Kwj4FxjUaTOQOsB6XWSQzNYw+YeZk1QKEoLLdRcgd0bAfHDiHq+6fhkf0j5mTVr3
v8g+otWfi2bI+85HtteozQlb/MWwVkZvsxMa49uZbTEWOD1goOFgQqN/ByFm4acqmYOIIlIq4gl8
F1YAhmTMef7KC4bcz9sOGV3mCOn7y0eLL/A199eSbYmEddPhrM2tBrds0hm528UjbKpRZYhHP1Zy
317E3V43JFGuX9Y51UOgTrHV4dVFN09mJJlZPbr27umI4HCDJvbksRaMXDqNHYB5bpWEkggzBuJM
Lz93gqdJ0XpM5c1CIDuUhph9I0dvph8VcD9DbjZno60kOIWsPpojzPLnVgedxIPeUo8DE4wpn/+4
K05yGZWSzKoQQVZNxTdtFDsp05S397nDfrzT/axM9Y0wNAg0yaJhuma58PLj/efBK5f66LSL7Vli
Ye4bWDjX7ETIGuOHG5b3Bhbtrped+S4eKQpS6Lgz5egNNYCsANVmfXVd6/mmj4H34sHMTVrFdgiM
29Hoct1mmkQNaLDZHCMuvKMzbWqlSC3lyoQcxOEKcNM2h6voNjAjff90X8KZIGLn9erK5C87wW8L
hA7v3NdLTJTlkSNNXOYIp4Pv29RrVNxfKRbAAvlGAnTO8XSA6G24k1oKDw/XMG/0Uqu1Y/+c0qF1
IL3EUTMjeYzbGpuH2j/Gdvc5GmnJBG/opmuSgzyFM4tKtzrejma4X3WcRqtznFbrwkuNDEdpVn1R
xL1HDpXoOdNhu+3zEiu0Ol4yGJZu9KYBsWR896wr3VQ1i69W5uOLNjG6hYLn9gCSo36bRkmM+0MN
4ztB+LW3V0O6lBtB12OOcopX9B5fKkQhaVAspIGE4sgnlUNu3Ndotutf7Uq1vItww2ONYSJpjn2R
Md4ngmg51dO3Vb0Pg8oorjwQ8h1XVTgaJfDKTU2D8lNHZK7KHL67A/9Q07d0pRDh0l7BTzHfNoGt
hTCP47DrU581Lwh9qNRPng7Wpnk3dJfadGPVi02Hfq8+dKyJ/Oh8/Y1lgioljAt4LSU373Bz00ZF
dtc/C8bk/Hpyt+S89GJ/zOcsZqhne8z3Wq0cHuwk2n3wxxMZ50KGA7HHS0SspOO8Dm8GXN5pqlF9
eNFJvj0yIWzs0PqLZG4GQBuopNSCoRtgd4Cirn3FtK/xb7fHTYncWgQ8HcDqHjk0IciZpbBQsFcl
5NMcZ246e6KPBssZhcFQsUV6zpwuUHhhdeKZj6xgpe4s9jyECZ5SHUus128PrC3266I1ZuMsWkZz
xmtm8wKv7JdLIcnHW/1MsEtUSUTYUkf6kAaBwK2alUnj/OZ+jBVXR6taP6XJp1w90sW8fHMcaugS
S2wcXyedNPSjnWDZQ3kHK0lSGcA7OkSssDmQ5nLkWDqx4eNf907C4BXua3F8zAFlApFp5oxOy1mZ
BbGDGf8Y2a9q3pD5sARnmujqoDZj8ALnX6uwSkzFUEeW4bsJ3fSTizrZwErrul1TSBpAYvH+EB7X
rbRykA8JWFh7clj+wzbhvFxnkHvyr4aRGhpweBGnRDIqT4fT3gracWm0Qqq/jth1fw92ab30YhuQ
s01jJuU/rcONttm+EUJsKYBiRdW4tSAzmS32wqRQk5W8A7hJ40GuEL+3swgMXOpeE3clTl/5DWed
5RDMXfvlPJCMthzHmTAYXZ1q/6rve7kV5kPjYdos38diNrQ9pG4chRJdhD4MB1e9sTa39VGa1USK
iQS/lFSWT6cMET2Qphrn9q7srtqpkGuoc0sN+tebYI08SNUr1eVVbL3kM17QKF4h59ZTriWnKatx
rzeyc03wUjTpni/R/pXC07xJJ9DHZ3RRTvl4erdfR0qLKtgc+bhXgwrEqKS7fX4zVqFHnM7aSNZc
aVVgHiPR2sJJeDGrp61MagIKee0IBp7Vk1cTDNIAJ4z78Ns/LckUg4LBELvhpFnYdUnGemDVBmZ5
2qO48b8+FDw3RDKe1GTqu9C12GyxnJmtQGSNPkfi319Eoe95FjkNaqRXDNzFNVtr3T1jDRGDBTOF
4HA5DQjS6KTlfgpfMQqcr68+oTikf0sVGxhQ6psgx5nye33L1HUCUnvSQmlRLZZfznV2v0bKI2FQ
HutC+pd6aGjyjK+Dnirqg+VgVu0WHzwGWO7XFQLq5DWBboPH4S6/BiRhioepTBo1qMDAZly9VDTd
LH7xy1awZhEOgbVOZ5EVFyHjd5yWq+8NKcCPm7/KtleZiXw9KPJcy+7lWXMxB87Fd5nkFERQmlj3
t44cizwjLWjDqp8FxamGKe3eELbntwxUeDi39C+cmMpMCcU0NOi1lbahwYV7w4p+b9QvqnYv8BfR
zj4zeCIBopcXOp/aEZpxbKkwQWYh9/JfipbiZWESDShD9OJP8nY0csb0Jt8mtoCJ6Lr/0uWd4gIT
0/Yvm2I2AQRlK5jWtkfE/erLrD/taeh92OCZUxHdIpLWmmz5Qwtw9/8TapVmSsKb1dBVQAJwNs5R
a9NIXoSyVRgKnVIXJUk9Fxhroa3og2KJrnuLhrHVJkoT16dZrpdAECY8EFgXQ6QlGj6mi74uJeTT
C3FdYAeDMa0wnDWug9dqpNSB7fjQ+RhaMg+FXOXt92204kx7UgSesw2BHDuRnw3H0XU9cP7XJpAE
BYSNhoKUCPLJqMg7ossrszoy2wcn+dueHI9NhfkJ5ugTqIz6EJt3jVRE3mHZoGx6GpWsDOToEvYC
zjnbmeqm2DxOtfwZHrYBCsLe05tGJaY4YJei2Y0sMKL0t6ml980TzFMLLSBsn/pqpgCMs9N77dpP
kLfksIW/9+Bnh3Em/KGBF5DwtQLuUTghotD/tzY/anWidRWORkW2cRu9qbymXTQuiABxcBp8OOIK
gckMCc9cx+jquZ4U/1X6q9a8l5CZTwgBe/WC10OAo2/DhiCXNQ6hZBPCRBKyYFrXbMYvrwJrIiaX
2Am7gZebRaCTdZnt7nbRfbrOO8egYjZkfeNzQ7bXoOreg2za6sRkhrMxQsRlH0qilx5TZfjl+PCB
+rJYPTDpHfHX3KPHyzR+IcE2JNPRVu8JMNG/fPEnT93tO3pfqk3oUgRBweT+Nn3Q1Bxy0o0mQWDK
kmQb/91L4IZnqmVpI2ksSXml5mpwsJLbEU1rrJJmQ9G1zjTGCwOi9zgOm0M+qfdL3hr432zsmS8c
1v08uHbG5+dB/9WXjNsIgQthfE1pJcP7uyziJiZLPwkkuB8SwBW5310T9e+fsyktzHTH24OsnyxN
LDccdtUGGXz5QZ+NV5xRJ6vevI9aD2SUR5yM8xlbWEVbpuH9fSIWLLLLw5ynnYmt6eoqMKSNtRw4
Bcti4pKyAi+oa/GhYmhGKtURpeIPJvryFryX17q0tA5nZyNUJi9IbkY3gOM7lcfcJESMEE8nagcx
wsb4NSjgOQXq02MASsLcAbGXQBo17Pm7Rxu5qRBlKK8D2xJSSSKxlsrIHG68nJF4icVDgwpoIrDT
8T33kAj40pz0A5jtZCfnMz886RLfD/ynZ1cFdOZt9quGn3+D8NR4Sjh1kIpYmHTJIuA+p1UC4UD+
MGiHheeB9niL9gjQ1GIl6lvKY5VSIAMgTTBBFrjBKLNogSk6tohfd58BN9AaT2Xd1jgQutlpWTM3
PdO6DdWX3o+eX8DSuLpHpdy5LM5cpmX/6n61tGc6RiNQ9+WCWYvrdF/u52t1SQRblXWAJ8aRo0jJ
fFN1oxHTJGQ8JO8Pwqz8vdsUowq1EfRafrrHCznUz4NT0qp1lcHOYjicrsI/IOh97CKOh7TxCIvQ
QHtE7He+a3XG2XHpWSJux0Jrpd7MZHKDAvZ5Opw1cCvH8khzt2hzJQgWBNPGgMazh2XMzoZsw8G0
4siCtaQrTC9zzEy2yqZUN7vusfgPRztmrmeqyD83tcBUR3xxl245J0wpzHUoGRTQouDs3pICqDA4
B7dvATA+E6u98TrdYrWPDGp1Jscugo7mu5jbvwSYAh/GLKrW8hAl3B0LU4NAZN1/pwCu07B14hlo
cqGZq8mnwZqpPe3cD6bOuJzg2Y043ZeF/pOVFczMhAcNRMvd19hmgZNGx02FJMA5BVRlj8cxsGJt
hXyTYsZ5HU6TxRAfRIsx2F3wXuyHn5OGlusO2x+e0jPqdjnf5iSuwSsgUXYtr0WUANSgH4fQt/w5
FLIsieb7NgbR/Kfv3bjNcKIivNI5ezJ1K5qECyb7IfhOorRd1bfzGWn2ZQs5yR6uZgeSiOfvd4wF
azfYAs7bswVi7CEw98yeRFtARH8jWIF2nQx524X2W8iYIPD4rNJGXRuVZ+I0La+e4FvVhRQqXKTO
6NIYqVVPKKEnLsS9qlwgJavMUMNDmEEAdzt3ciojaBdkAppR0FTNCX6TA62m80WZDxASjpbr+4pu
ymFwy1uUuQ3IUGso8ChmGTgXmYPamx+Blpy5jErGyUHHxTI/lEtZVmLiBuhxfv/GA6O1iRu0NdBa
HZrrSrGp3QZTl1XNpwEO3lS3pCReqqHYt6Nkco7+RRSpDZMm/Fp2iegbQv2qPi6BCehY9kTEvWwh
FIQNE6rvQTGF8YNGgbJnV0jx9zQ8EJsJ+ka+Q/cBswFYpOaccUSE94lsHAT+b3MFKkwOC6luq+7F
TRZnV5IsmDTzyELZKUR2hYg70r2kVAGLruk+G0f7kaHrpw+CNiRiR1OGJtqBYc10qRUe2tocjp0d
q2VM3GxXBExrfwV0Tj3+RDfBwA16tUcQW1pZAxexpM0jMMwnWvMXHMGqe2o3747TzF6srswWBAAA
SkjT0Ui27zMf2f7x3PIHZw6rHXaJUxkCrtpWcpg/gfd4rdz3vpmq5g91I0FkzrC6jmdQIPzjUh8w
qIXzX7KmgSOULSga0z1/nFLRmIIigKjgvYimlgnvvh01F5YrDsWclXxtJRKT7YNxE5FoiKCXxA8d
sVgms+YcddzpFMkHgTB9SM0eR3jrnzjba17TgfUnnWXmUo9+5SMqJMX0rZsJTgvjxnwJxfU+ASAJ
0z9VdwhYIUpzFJpKgB/hGF8rQvUw9nD5fqlz66n6Pb+8R8a/chj4tfRFicVD8LaLjNrCItvlqFxr
6/8z6EpAA4Xv7oBB3giwunAFzTIi2DFoEVsg/0Vee4ZQe0lchAfVx65/xQinTLmpJ5mdV/UrpMFS
+6FhB/kzEEQH4BDC64RkCx2TcOSUoLmPZU+29p0jGVOU2GyzQS2NTv/vtc1T6j9iaEmrzV7YB0zO
xLo4VaSZxtDeYfZe/krlRU9PzzET2cs/Xmdsu71LsOhMJtQaD4Vta9jtFSRQhuSC+9fDFr9xTDV4
CQu/DJYM1XhgFiAl1aZHyWsg3x0ohpq8xjrOuckubDl//fP4oB8t98kaNFbYLmcyhzw7x7TDlr4E
XgMJPoA0YEnv1iQ2qpRfZUEUAfYHPChKWbWw40+3Pxw5qTh/oWX9WS6bS2owEQmh5Q+P3/w7zg0Z
0UQX5DZMw/nQ+zhihkkuHsu4bTnhTKAXOAWdwrOvZvixd1YaCljSUnuztzjRHFlR8KCNnngQHpsd
bAgNU1U4mVO3cMXxhmbTbX3p+Zm0mFDfQ5GLKnc+0gI89ogbvfnKZ4kn7Tp1SuXG+R+mhmDrCjzV
JzfNCEzjlutIk1R9N1VdIp0VAN4BTE8g3zjsTsFWH3wOC8RIEkMUSk1bU+pItuhAAH2ndSTmqB5T
yRG5oXZmi6r06WybeVOmezI71y0dLWtmJNNQRIOdsM9pJLePB9s2IASWY6G7Gv+Fr5TdHUuEA9XI
e68WrMuHI72Ljlgf6MBoO0m6E6PFdHG7Xh+XAtPkXMGeEWVBLmRngu7KZBA+faVnw0qeGZZBKdQ5
kqmlKA1vs+OHMypJbHV7BPb0cKM9kiavbapyUbPXH7/O/TpOi3JDs00r/NC3i/jOv4VBN8KL8zgt
WQNMgj4Zt/4khBvcbpJfCls5gpRwkMQN/SkowyOEv0Ow10e3343QtCoASCg8OTqxM3pxDNmqedYt
n3fNwOf33cmt35uC0sC4vshOMS9mB1nKfcvCqaQC4sTi7Ez/6S8H7vWTZayOtHs30kBvWRTTEiye
qouMU68sdk8nKkerzvHPFJSHah0QCI+YIZBPBCYdyqHydD855qfuVJXsbqMzzPQ8t4SB9MnZ/Qfy
uKah1fJ5MTjGRbOMGhnje4MHIKeFJR7HD2GBheJrUu88cm5gokhYvhYDk+Jzne/BrQSlFfyO58pH
33SaQlrLAX+f3OC02lSWb+ZbKdqjhjgMxD6183cHGvGRfMhTYcDLGod/3b1g0jlJQZ+WUCg3+6tj
HLnUVXrnrBpywIye7H4g4Q/bGi95RyE4WOQt8sBGJ+58xQh3YjjyccmLf/vM4lOJpGJ4iQpvqHMi
isvLeXS7Zmi8xOZ/VDFO1MFFrX3PwIu8Qm54jY+z1uyNkDekWbcroJ580r3J39/G77qSZRau5URv
aGHVLEuPMUy2dTqCyZmi3iVojVygoC9yDLX7C3l3wKExMm5AtE3iG49yD0qNH+AI9A7ojreAMZ+H
6b1tMQOyXuQcKOlGvnFmZ9x4jgILw4kD7M/xU+afiKC1XGEPBQQ0/Pxi+fuRYP8bs6SFDPD/qwEi
YQ2rpU4c0CkIkvaDBnPpkq/o21nEUfHCtDQF3VAC0ah/G21gkysvYD0dq1CgK+KYwfB6ZHYDC7Dc
3oLEfq8Pn+IeDAwEx7nNQ6ZLP+gKNVEV6vmmRxTWliaOrTdPuEQv28KxJfadxYX0ZmU1pMTF5UZw
WIqu2VlqTGVZ3DDleuKs0/R/+2a7N7shjzn0J2h5fJj99272JOQHW/Fp6gDkVfvFoChETPDovRWO
vu+/bCn0cRZGxUsmWbEuWxK9O5gsVT+z0006i7dj5JT6UM1qqyTBnZdIUZ2qU8qavky9jAwuZxXX
d90XVBo5tybcar2MVWLDLSmtbl8tMrpyYrunV+K54SYoQeFmRL0s7dGgwtxq+DKkp+wVoi0UjSzJ
zrpKoXISoOjUGxJTUidq8a/swcpHPEuJgz1A3FIcn4ugFHEiNan0kJGQXtmamZ8oORA014MVL5oI
uFifG8tlCd7FMyamXxzaPHmWn59qgHfpw4r8IaHXI5Kw+tcvQExCoyLPlLUHap2QXr7/DoxYyHxt
vWxXuMp2vJI3QRxe/YtHEyHugkuvx4wWItH63NvsHECo8yySKz8OQe+XeO002f7riPM4375EdE70
w/6qZkz+d6ECUYrsXyogh3NdlmYGplnm8mho84pgF3MrE/BR1KJY4dHvvXv1mgh5VVzl2ZXOXrbp
f4YSHwkY/2BXxTojWUlZaCquEvHYOtfR2/cfEiE8jaW7zKOoSDFP83B+QQGpSqtdsC47buasDgcc
8tH91ygg3BKXXjFEtjlLLpELmMZpJ+P240QWBBu9nnpLdlHwnWO+A7/mDPnHovy1SrCRTR639rMe
ZUjtxQec7UPBQMU5R9Yd6l4Sp6rUnDOXUMyM3Dj8/KFkNtIDPPIFglVPBf4KbTsLiaBIfsPmC91q
NEmOPWAyYQYGUcGYyK/LfsQECbnfpkOGW+iJ1fpv3mf0Z/CqXTR/+FeC5V1Mz9yRM6GhhFvYmaQO
hi0dlYmsKXjR5djxve+xYAtkvgIFsFuHI6w70HIPmIoPAemIdZQzur9YBJydKUO1g/xT0BZxchcS
Wq9VeeNxGrYbg2P1q5+QDBZP/QrytaKiwHXiJf7mOabbZiXtfyFhT698F5nu/COcvDi+Zjq+m892
9IDOk5tflyAD+pDf73AyCmsP0gTJe68wFKBaZYYZ062GxSWCYKqBG0dQiFksitOT4FMli3hWAbxL
64oSg+0um/qvAaleIkJzJGaEi2tnrRMeWtP2dz/WiVe36Uof2ZgoPJ1QES1+VjaAROeB0WK3z56Z
FeuccHnAe+8cSRDFf9h2cUyg4iOcvbaVjEu07K0RLPTCssYTQNSPfhS0P9fA3PW+BBnLXk/8MF00
P+rAmFQTnLOvNxUPHCp9FwsAyd/4/EsvPyPWuimGes2UFg+z611oc32dHQKpBUaUsbmlvkTr4F+C
yMuEy/mNRjyquQ6yYUayPd6C4JBUZ0d679EDt0VxkMtBdncHT1indE53kj34sLr/kkwpDqEJ09ua
W6sJjj/C2+v4ynKcatNc43ZEZLNFQAPVpfdgiNFJDGxd4WvANZ5QzGS2o+InKAxtCZvIt0ONx/2u
nvkuZ45rtD0seQgTXhv7TJObs8HFI4thY8YG2Dbdy3fVRkDro0Ah9VbWTZyJqEn0MkvhAYssW0wp
iYrDcLBx5RTvNYAUnCkEzKPqgQ5Efv1rjowONmY7Nab/VuvIUju0yfoZCb9+JwVquawx6atCqVd2
NyVANAFecfoe6LKWtOPSmmHeiqzhhaG1qyGrpDKmCbwldj/udnPqTeB8toIrmAji5+7b/dosiTCy
VOiiwTPek6oqBBJhvnK45qiY0+9hOQ+JSss5YFCD92JjqzC4lUElzf0m6YwC57meFPKNHLSkUK80
hb0evVVGFvKurmXali3CRTKsByvwnXvwUxkcYWRLl87Q8kffckH2Z+MwFQsIRs3Urxh963i0Tsjy
y98DkAAm1V5i16n8/ySNwLjOSs8ekgA3czKW0MJ4Sd30BQ6cpIzKBWMfSBVNSXioVcK7RL0rzo7Q
judd27N5H8OMQ/lBXiURhmpLr/KwoLkmnwfyABV2js8KoEo6KSZ4EENGqy88rO0ClmgjMArr2Z4W
2+v4kWUYssURggDILK/PYq+bvaKS8tuEFq9U9s0CUVTDB9m9Dq2/751hfqYx9Q0GTMlsltdBlTqy
8GQURKk9rS4wCGazEwHiQJtobpuG1aUZcFIFP6oa2InR2w6irX+YQGnOp8UUsMr3lgbxf9Ti2FUn
2DpRq5/4VSjMCctbMm76kQsqJcH4fHhcE3x6Q9qwnxntbdBcHpfnH8YYNX4XS+AutpfJQ+NprglE
OB8VZR4MnCDb7PGzC7jVBnyIVDVGnOVG1qM8ZY5zQoICy4dyos9ebI77/9+7SC6YsB5eKwjBAgiJ
jRih6ui+AlS3/sRyQSZGu35GSSZORxrU4cjPcNyYt3NXfXZfArbFDRyJGQoUBPHcmTtkQ1tYeJGK
+0NBwg6hXD7Pe0cIYVbz+O4Q1mKty453jCS9v6q7H97Z0xphcHjbqAw5NR+j6eCBP+Qk1B5CHIIl
8G+yDdaZyFqzwif6SOGTt85jPhNXvDRs38nM0U4RhsgZh4tmx+UArdfCTjCr97f7D7zMHtGJ2vRz
RAFe5RvOVDzo5Q3XflYkfaELUnzcmGEgaaNRcvlvhc12ilLxYXO6cTg42wZYGObRkLq8pqiHiJmA
dBQ5Jzn/zjOJPkEtnNCrcYLHBLQKKKgioOisfKljhZI+3SBJEr9taUtzx47fnnYRxCMUpUWPFsuT
LF3XdkZjXj/hXZThkpBBUftGCtJtDGfylyJlGQA3gtXqxyd1RuzBSEVpSjHqiZxGt7/aEnO6vVcP
km+kJb/TQd9yz67qYnlGraHL3fLCOjMOdtUR99eE2RrOMFI/61pmG5sr7E7PkNvXk3U4F3Mp7zNc
nsQi2OR6XzEY0VlPQNR9ns5bkyGJOjekS4jSbd1lJn4Jy0J2bfQ15LG9JRVU2ybvCkddn9jcDv43
1J4GEJ7VpsutIcMIp+R9wdJ/yL51imRfFMETaBu6IZwpzi2SuyUUUfN3RclG24piKhitaT3OOeqN
yvFPc7p6gTZPYw0xsTSMJobST3v5NtiMXAkFu3E7iYBuEX2JmVT84h+8cHNvGsETLmPVq5S6P4z5
us95KcI0mMeBDCoHC1BZTdSinlZGU5OB2jQlERsjrmR2z52cqp0w8+spuRf+lMdh9qVpXz9pl1iW
QjUDCaTNp7GI7XGQ2NZdbn+mNWDd+hdH8ukQFY8tlp7lmjN4qNrtYpaAegcU5aZ0ffJ15PxbJAuP
c7xh2tL02CdA2bNU7YZEp/ZK/j6PkPDlGn2RUobPSlmW95FbynICt+WfoyGveuIeWsxwVvuf0d+5
z8vZeFJJN/wHAsja8LNF0Qk1BbQL1+BSsUiwIaN2BnLbUBVE4/8lHzMWFSI3OSf2ZL9Bjz/JFU7N
4sLXEf0wMyf96gN1rGai0wytGiPzyIRX5JakXDd3xHez9gEmsxFiWf3gh6ebQLiL0J9rwbUaNJcV
8fO+dK2Am8nElDy0s05eA/uTHjvl8s8mL7pTl2SNvwHW2Gg7vJzPTwDwUT1p7RMQ14mjHH88w8ag
+qpuUuTSlI9x0OINaPX5T+XMa832XiIup+1LTVXqUvxQfD1F82OdnLghL/sRIt3cqPp0IyMF7zte
o22y8zTjGqc16qv/tv+wjHOzNTZnnCcpuPyfh9vOoMeEd8bmjec6kpdoPQcz80sYIGVLgY4RdSb0
ekUCHSKbH+539hNrggC+DevHY8c+8yt5794rMKJofcxBanD2Sct0atnBJsSa0Us4GIzWhTAzkLhI
q+qr5uk/hA7+DhcL8BO9JIk7uEGJPrv4ryolBuvsFmlgHVnlyVNMF1BDRifJZt+j9WMDLDqJeODv
4WcIKKDf2l43JTx8aZpEQS7A4DMz7TbxXFuiKHylbrvoUxQteRDAh8huEPiCy9eU8UZbVVAkyvmQ
cT2Hg1C4+OezOPJZk5dCGyF+w4cBaPLe4FVb+ID8eQ0fdHTMpp4Rsdw38NOy01NlqcT6GRB/oMug
8Uq9RlCzngKX53Rx1aTld9/XF8ZaQ4ShQO3s7+sT+ub6gWW7+3fEufXcRY0djMla2CQv/FnXmqrf
rUy6Pax8ezzZaFiI4cinRDLaqz285tBvR4u78ncyqykEbJiUnS4+DeAHe30kOwN1uwrEl2sq+94m
MOy0o+XfnljBI4uJ/CzYIu1xGTdEDZQ9LtSBaKOPhSAyNz73/79WmAn9+GQDzM3hjnR5Chtipa+a
+DfYMbeAu+jYxlolVdroaoeo6MihijPa9h0qTxpq5Sasb3v2nPoQQZLbIHrPV9b6iTZoKfkye5T9
O5S0uWe4oRhNSWIAh/rrvaOFr/iMvfwmEDkC6IhCBUHfn/+9KuDaCOCqcQkI/dWzZyeFPAvvF6kA
he7rj9PRId3fqJThLAREe4AuldmjjRTVvCjnXbCcoDRR0fJa00NHPN2bgCWTfrbudkJAxcgSgrnD
9NvQ4r0mMFDIZUB7ljUSEYCS38mgS4SGqOIC8jMZpVRTCmHhV4D29tKzwRzaik6HgkoaZuxaucme
u4R3IaFVRJeo8oO6ghkzNDogviMmdW21rx+f2B0n9nNQEebHm3lLTov0oeJGkUf7SdeJmIELbBPw
gD8TyI6zzhSRSACJmMPyc35PeQgfAkhPkoee4MJHNEXZwYNWyKkCL3xS4LzMkmMu4XxWGrIhZaZK
2qNyhgX8fuwCg189m8OXkKezCSkddIfG12U/57Q0yNO+8chldB7AcS+qxeK4eYxXYSxkTN9sj6mg
hYW7ivWCFKqxwDqpjSOZA8EXdrUGxCUTzS38xQtUUWFIKgW8co6+RSkBoeffVmr1ycz44It93vQD
BSvOYfVN1i3yB7r3bw/1HtjVErYM9DEiN9geIknJco3Sxbwyb7giHc3TTNBD4PastsImwv6OlPBQ
AevxagA+sOedqvmr/W9cszVO8uaetut7mr9C2IXZabMvUybnxjjTbJU8vRiWOUJUXqIVYDurUnMK
q4LUgNq/yZwu3eCuOO+aKCGnOyopBvv25A7WFMHfNGGCo5IrM6WrcZuVkJkqjWadYAqfrxl8ZI4A
MweytCT9E423swZrwSAV0XoETjFDI0NDHGdu+jPR9SiPeSe9GkfvRyM07xnIVAODnZSLsOrx4bCc
VkNruddb8kUc5dHpPKaTVwe5BXI9/T7cop4jCqVTYTP4F+SKme2dADQz9ov1clhgO7s7kF6YnzYZ
2xkY8A3aygwfPNjQNKrLZG0gDi19sMs4DMi0yl1qthrm2ZleU6yhRiK/KUoajLI5dBunB3SGqX51
XRec5acy2m49dLI0P+/YuQoQRyM1qnQCk4JzWiA1PWcF10bxbE3i/QTQpyKdZONFGD51biwOmPKM
r4sLWfkQzluVJv32diFKg0N4iQlfRPRPlii/990nv7ejhDrxaTuD/6uF5cxAlJLMn3akwUNWj3Em
Ms267KQq899/5e7T3k1684xNbppj33Pv6WF0BOprOQ93OftpiXNcp2PLj+dVSHW70W+rO7pZFcYP
mYMCnDhZ5+5g57q8C+0E/YSsghYbE+f0AkqT3rA7zHAC/KF3XQ7fqH8tl6yXcYX/3nO/kgUZTRau
h8Kf0upCK+B/iUTg00x3ZDCMfZL4Uc/Vo0fDhXkRA8rN6ZsYp5quFMmd4F4/ezU1tywA/2w+GhGx
ft8jWYiy0wEmZP7NKegkxQaa/mubGDpuidPNcs+cUqWKEReSi/jmzbuiXauGPdMECJzrWeCIZslw
fsvSVYHv01rUBaOpj4R7miEpsYYh9mI3Oew3wJ6tideutGz/w8p4KbVcDwuUw4caFlyGaJbPyrns
bQWb7CsuXRSgPJMBLe8+Ypvm20q8NgyWaqm58qTMZ0UK7TZhF6gc15hiREl+qqTIkNmt3+SUH1SH
X3eKJyIBDtLC+os1QMHO26wojIjFFN5w9CSiDqX0we9Ltd708Cae/2hOun9vyr3vrP/XVxcsdgg6
8rDS7jnWirClx6rXD4IsMl9JkHKuy4VO1vk6puhDKpcB8dU1Dm9wGydE1QR6847MbpMaqna/Yev+
f97aJoY0rDx9i46ql/gCmtZ+dxZRE0Lkh8QMFIPbcgNc9zEfEH34nhM0rJ9Zz9aSimsxLrNcKY4F
jFTBxxNINViyzbVKAjRiEBlTFbVQgA/sIDCtfP4/UH/RW04ocwmaOWdSXbC127mPtgvymH0bA4az
ufUdXa8zo/9RyoxNTVVjclwgGYbYFRZyKYotDpACn33tnXKIeYnpvpb8q/OgMbQ9pZqg3QO9Mv8D
S8GZhhh2XgsyfLjpfsyWKkEqMIyu2+C4mEfIUbzB481/8uWrikZbGFzCwnCYmUHWevxmXIzQRWay
9bCr7/Au6CdUT0XW5kvBp7pR+gcHg2RFxc7RMVUUczJjf0f3js+xL3KJT7uC3G5V4oIHFZA01rFw
1MKdms5UkG4P6Si/BtYA/O+yU3KzPOtutXOeGZkw2mhxGGDzeSAADPN2jZQtU9PsPL7HzmdGdbO/
8l5Z2F50KNBOVOb8CENxnAFWYktC+73X3UIAY4hJ8fl32fGzkHfEtxKqdv3cRT+gsnAOaPVX6ibr
YNXOzeFD5TH5ENhmtX6jIfLuKXkY90sGwDOiyNW35/RrAqyODJ1cmS3eMO+fPUjdhsOlZGQ4f9Sp
xuqnDd18wuNBdY830XWeozK58afj+jzeooqty5bT558hiCVRgslrNq8HN6SIsiXXV2bEw8aqiRvf
KL7uNCA5NKVXb5KZ+FvaHAHh31HNubdUyMD93i5RG+nZ6bcx9HRW6LfccqIUzD/Bp0ZvfDfiuGyI
rACQ+ayJUr3B/iW8jn0Z/pi11LluhssmDv2ig1oF1ECOGKf75/Y9ic2XtWqKyvZSzU0Ufnt7K4l0
+JKsnTjb0PUhPPTiOy2q3Vhm3VXMkBPQ+txScUtb86K7/v+eZbGtnp8dUPMak7ssLnB5DBimhZrN
ovNyGkVV6OadpVZFiyn0/cwv1tzWPPAxVrVhEVSU6rrcyPy3ugIzqc9MfEHlJiu+NMYN/XBfE7v9
vEt57mcmrMtWvb7G+c11VHT3EeJ1EU0IVXV5AyKrDlGNlMfXPmuNdR1AkH0XMOPxxBNWeR4DSp+P
IXIoLRBNfHli/ZU8WL52Z36UYp9paLzEZ7qBkn87RktuQXtlWYhMR83/LXKC1swUdY86aO3VdLKf
dITkeXGSdsA4bdXuML9cxLeQ0K5RbWoxBviXLK5Nq8OKc3okq9AegHusZzx6JBpKZ4BzLpdHLtlb
pzTNS22nKnfFB4CsYe6jTriekzX+styE2Oad9+1ObGGsSS0LthpymwsIWc4iSfAV9FaBm7WlucRk
/d5az4ZZOHrbNpr+SSAIeZBJoq5Lzs9xjntuZqk9rLPwN4xSzqAr+n6rZ4jnYG0V+Q8Ho2fmT1yV
mYkbfKsfzC2IXH4YiugvVmAo2ZP8Y0i/5rv8o2WzEoBKFXl32RTH/KXKBbSmcgmN+yggL0Qe8jex
6+06qlKclQJxvM60uvBcTsfNTSqxk9sHz5Bg0tT2tNcgoHZyPlm0HxlsaARpP2ZsNJNYhdCo8BFl
RfPEmJMzdtMxA3dsgAHgw3WFXGTtait9wpiRiUZzG6wHq1P05fKEnenpwIxSa1rw9VV5lvNnZ1LD
9+pR+jYdorZdFI55MPKbGBIRbKYsoAETD8UhYERo/GfzLppZS7yRtYKNGDkS4HUNduMImjuolahW
oPFDNLF3iyJPQfiszMy4DRBEOwyAgPhDdFwua8bewJHsXW5Y8w5+5JdFoK5Hk6ZyxrVrC9T2k4y2
XUqB6xrmHHY2jKe7S0UH2iaibX2PVvP9ex+gogv/WHiL4WNPUzne1baaxBTXMu7UO9oPdB9dQEB6
u1IMQXsRjpOwXGnqPJ1usnJeBEJYCRbq/AhARViC27/l1se3+bG8cFopt4MaicjzlX+iMxJe2TJ2
gaZE1Gsp+qYws2srToshSSvRKzjAnIP/q4T9oJIHzh4Ar73d6GetZQihFpPsY9ySznYSC8T1DS/s
IcTTTb+izFl2PekHMtXG8CVoEB+GqosVnMOECK/npZuBMzwIaBTcYKLUpteiWXTZIP7y5DyeD31M
GuTp4w2VS4JUVehr7pODuVsqhCRj1xOVgvHojslZ5u2VGnHbeJWo+B++HDuPTrXdk+rlstg17wWk
VryCIX3yXKr5Q4u77FPTJKOP+yio6rc2244jeVmuXl5I4eQJ5+GhmO2K+TvGwrUmXdXIZ+2yUJFO
KlY4QBGsiWbtPxUQOzPqKDzcis/8O557JPasq4mNyWbrqU8xl/f9gB2GlkoiOm4NvL36qTU1dhMq
0UEggIg5hkDRfa3PFIDSsL40/dJVPuDIrXTkzDAcUAe+0UHI8iQYJDh6UTniLolNI+upPMkomwSU
XL/X5bkPtDjjggRpCwFWC7nuIRKU65fye2/Fsj7y8rankDGIXrgrAt+ZfpglC/+YWDXyRh+yU2/U
kesBsa0GFb5Cvf2ZjEWbyjGlJ1V68+FIE236ZfOnOkBDv8AQSUBK77FTxH7tSQECp5HmB+xIOlv7
jCSS2jsz3wg4fxNksulWYzfc04Omenn+1LD590J79NGJkIgnH/MDL222zoQRwMxzj9//L7daS5U9
ZoxULYkMuZgM+hnNl+X+c36EegpzxxrXYoxlewFwtZsfzTvqJ2T+fL4lH6pgJXlP+J+Onb5OL9J0
0yVkG0UEMTKERRYDBXnonbKK9IzFLwdvJ1jQ1HWhds49y/pTBEsLmbOvqdfvd+S3cws/gYAmlZI/
G7cGHpRGkqUfxnsz5mKf1kcOyg+q6wqQqozvNbvtnupbb979SMqbxNAI8ksyN5LCDVvA5SL6YW9T
+sR6lnVfP3B2KN0TnQtlHY9gj1sPOazl8AkG0oqHV7DHY7efNEi5QmnUMiY9YglLlO7hQ0gEvdON
3aVsZwC78gJ1zA8JLNQz5SX7NvV9IQL1KQfOQsvCp59OyVx3pWvLqNbsNJ2mHpFxlg9d6pkEDx8g
JN0poCP09leul1lGc/x2zY7LMV+iB1SxklXXxAV4m17T6zRJ8DdneX4oeDg5+3yzAYHdNPdMR9QW
UyhcR9oHWRKhToThVi5k9WXDNE3BgI/qvkUm5uu6ChZugUL6NwBb/FAbpGQU/SvxhCHsTD8Ozqi/
BYRsbwrez9UbgBKY1xWawM8qHo/GzIOh0TYUtrUUHNhmb5qQPRBU4/vYP/ld6Xerz6P3EE1LNtCv
qnUWXIpPY2pmwqNSJnEzTm24/Eatw3c/+jvfgEY0J5YslnUZW/Q91uCtcuREXbwnmsg9VKGi8I9v
YVbdLOL/Y7IdZQ6TKjx3bpoKjaQeFrjX2cb8+glsS/lDgRv3ECLJb3IofPrV2frGVESvZzX5FMZ0
NvHv8IjbwE1CR0e7ZI0Hydu0+WuXNozrH3goacuz+rl0jckUT8EP54P8ruEhNvBpTvfffND98qc3
nEZyhCrpsRmVMR5qVdr5IDftWavOWvo8QexAvBJzpzb+weZCeNRET3ibOutmYqc6+uP9zSLZThnz
aXgddjNyAzs2hnUAx6FUPmy1YUVybG/wsbFVFavzHz7QUOYWkBNs60ANgDz/B4gxXXe6GE9df84b
dHJm2eKDBv+vhv3RxZTDr0B6EbpT5z/lo9LnOguXiEz5Z/+P4gcE61cfdIuyNNwwx0DiwgiBsZ8S
xu/2gL3fi5/Sw5QTje5aVJUBTSh8+J0MmalyMg8wXZwaz/U+FywCRrA7hZMSyX+7FdkWKezd7pMD
BzSdJBmI6I+sGiy+HEniTQROSl7251WOITVU5Dv9Oj0cXUGc1IjTF8F02fY8zELwtGh23sEuXKjR
wPv6vcG1zRXNwaekPZwCqPi0xO9LawkNUWzBVbgiSC/vYf7OdZMCJzD+RQHKJKvb8k/7p3mDv4LI
TYAGNwzTq6g/+gsydxwbyp9AGWWdOOC2Ddb8aNDtoS0kDEAoFqcIIRn9H3XQAyY87mvphgwtKI32
dm533KvuxyLJ2GkrKlNmoEKpcDx7wxp8y2CKfFmRZibSp/ZH/xtpsJMNILwzho0W08/9+ZNVgPvs
yu1t5i35oUgMDcqYG+vYQoYtkpUVmF4qDJEIdGns3OBpsK3QTCnXqwZ3MemGBi7oMdn0aghabtmL
2ZSuB3YAhPkrtTDDQBTRzOQ0ZV/NKXn3f0KMe2oWhUgycUK7Bm0XchA5bwyM+eHluoLr58qooKhA
VuG5d9x6mzb84h5GD0GM37hwp5Tp++2WIUrVlxRs2ux99XjlK4rJV4hbGiMY00L1GDTYtPQryS1n
Gyl6hX43UalYQJaWew2eM/gbq+3CzNQcqA8tWtJvafJU0cb34lwx1Qutm33276cjF0q0xEeFQDug
DMCo1DQGX8/wm+ZvTLYZ89TtdNoPTc0aonmlgl1w5W3NicFhjArmxxVr9bBYj53ALHTTdMo0qUjV
ZkzdQ5S+DpD7kfRSL1zYeRKXq+FoFu8i0493U90tZT9kMuFOO2apUzgzT3HhKdtbOqJ6/uR5uPuM
L9SrnscqfoQnkAGIMMHzMXKaqyXXObje95ax1wXiiqlVs0a17wLg16BbNc29m5aGLu/MyqxziV/V
MA4WygQKujmaQDt3CoMhjKOCijJabu/JCa/241smwR+L1UUaYci19WRAVYwidiIoh/SbBj3ooUpf
j7kWRqM8+bBfpQGAY2qi++U2H5EH7lls2FWsEHoVEUaA1uDNCfmixBBP1QuYUBwiEP5JgWrG4lWr
VYNqFZUOd2iQ6yy3lIiIIJdcRstVbjy4VR+d4fPORm4+TRmqU9UV4blDGs8O61YEjnaecHt/yPj7
L8yKGioTnOVhz3fkjHQUBs8PFiGggzh9iKH0CfvzEvavYRcjBwqIDqR4c5c9NEVx+hjznCypwrMH
W9vIqk0PbTOtYpBobMvmayIQ5mJiFWxHt6GI1Ls94TBnENheVtqdI81DlCq9IS3cZDva3juzuW61
IMwu58BitXhhl90MIKtfF+xa+f3RXQN6Dc8BwM2yIe6EWArGJyJKLy3jULqXhYnLvSmlbX6lkaUX
JNvfmXB74UkzLludTfWXnU+3Oh1GD13FwhO7zbTjplgA/6zcCt/Nbu3Xr8h6QBuc+9gQwNiSh+aX
AFigx4fyS7gHigkjn2teFUKkZ2ysrFlAG1FiHs6x/8t0BW8ovKMdgwRV1VC/hnM5sql3uSXpWwF7
sXjNIR5wx+b/Uh4p0rwLxVpjpH2kVTJdPn7823w0IVPTH7dm4PbHlN535B1+q5t3VqlCRiuWEKvv
xl+0hjlo1J+LQ1TWU21Obe2giey6x0a04O/aBn0JV7XZshamqkePqn/tkxGiEBA5m/Eu51n/pTIv
2aZgBgd+lMiOrUpQB+CdJSfo9SGgIjqfzD40xE47mA+aj41wqtu7z+jGBWcsOjyiARKcVMiz4c7A
azz1x+WrBS+EFvsjrGPswPOxUF7KjzW/ZLbXHdKuMvZcCzqPZ3IJgHYgyCwWZnkn1Jg1ItsuxlgJ
gkHHVqUNOVD1nkDOWmj2AxzdasoiFUut1iWrVuqZMGrYNFgrLz0hhTVwIdxiOjHBJnwTpxARb6nF
Sn1EidFPCSOlubxQL3Ne0NsMDkNklFMBtMEhOZLd+RUxHW4/Gu1BD4OTfX4kEYVwZQD7kX2U9RyA
Pyru/XUoSjZ7WgLnobmsagDp+0d/M8GxXUwEYhWk02am6W7mYi/f8Z50VEH76JrwQ6Hr/vdYL9y8
33n9LoCTaAnKy88k18VdPKRgLRm6ztGw/I012QhYoQL14mrI3SbsXxv18ehaUB7VYPAJ6xwNUhok
vvGziSgD4BRcS1cXjSqXWNL1tNUUoS+DyBwQ+g+Ys5J42wzubzts5ukX/VZSyL7Rl03jxn7WzRM/
h3xKe6tvJVAP+5hoJSyTeyykXlgndGTJJ/XOyI+yNpIVkcEXfn11UMb8wWGyi804SusEdGuSdDqW
jCiJSu28/jrRo8YL0gspi2UFrpO2evXkNz0aF7mclhMblF0P1NTrzgfPSD4GCGRt4a5QMm2BKed+
+57iMss9jn+FrPhPssfDBGoMZscw7xVxnngizfOJualkV99/UFr16Kp/YX4v5jM8U9ku4I31nIKb
esgQehuQ84jg/zS7DNylOLZ33N2UeeDW0nqJJR4Y1W0GCgmwhC/s4toWg4UihOf0gR6349ZdtFFN
O2urTCfuXXxNS5XdqcjOQHrERSp1L1ei2qnD/TuTyaqC8kUgVCq83+hZrdXrvOYyrxbP02KZ7nhK
rzpBgErnOd9E7s7plvV/IdlTDqlZHdCx0RgJBYiAfy/WwnwP6WXTl0hK2I+J6fs8T/2DfoDHa2Dt
orAPhzVCEECSzT8/ApaYqUI9xKOcejnEdB3Mg0cneoPvs+/Q1N3nUSmYyUAzVLJ3sfkejXmnVoam
lcbqkIxA7FJX/YEGdanG1UaISwFrPqUVLtTji5XC7/uq1J9aTNliWpcmqj2SOdoG+xHBFYbPpBkR
dYa+SHxIWrDYDtEf+4jQYrRdMIgJC81KEcXwrioTKdtl96lQhwLOjMqCLGf/beu3AeKww7lyjIoz
wcddfwQ3U5N6qwSQCVYbUiHoDKFFM0nrS/RB3coFRyAeS711QGerF3Qb14RcBRgQ61/U8FS17BqT
UpcFKxWUgYLaGlMLMg4bK2IBaw09CHjZbn1eTacePtiZAZ+ECTwBzM5UM+5lY/kacdSKCRiaJ46S
cEdkircG+29HWkjU3298nrhGxyuibfoN2k/lElpltMWSd1RuQXQnwIAQaj/sXCbg7icYsy8P5vCn
sYGMmyJV9g8Hv2e27hvSEmHBtgIo7BplkhNszUhStz1SuxaKmLoCBu8r43O81wy1FvUr7WcEREqg
7EF4o1sIymfekAwiUe4K1aLL3nBmRMRZUsYUoAgV9GJpfjLYPJJFmEtnar250zn8aa7g74ocG+Nd
GA2LPBXXsmEBdx0cm2ZOH0f5tJ+nYVYN1793iWtR2D4PNJPIJzTZdriSwxCjK3Ti3Z0vjp+QzHFO
JTH0tPulXxuRXVSPeMoNGBEWKDXAwgcJYAcxwsIoav36OcCs/jOFPHEGNUlJmTzT6VZDbFkkHvNE
fxIvugI3aCVLTM7y3upoIwqM7v8I17+YDLhYKv+TUKCHah+nCddlXqN1La7zBQ98w8S/zHysmCH1
NkmYIwcIRzx99kDcR3YhYZd8zD9Du20oP74A0MfSUMg63fpTv2j2ZbNI2afUx2AfrWLVHYsNNUqR
HC/QYwVt5FpY2m5dwkaH/+GWfg05QGWFKOIbiMlJrd2u/E3OXjNKLmbQ1Y4DY4T5c3O9LIhy2iD4
svA7LazIyc4dQtqn15CqE7Gq7M/WlEFcvpOfZsI0LXdgTIeBCWQ01Je/vMFRntmmrkBqbVdobcJo
cyFOJhRnMrxP8eB9DZNKYLEpJCV2sk3+C5XRzTQamBKuP+hLsfbLC5bSE0c7PFgbSraJT2OUAnZG
fBQqenwkYWpt0NfeZ/lTc6LmmVWi7IpVgGADx0jOtDfiA+21agoNhF3o0Im7yPlBl6GWIno3SAy/
F5w5hJqjVXmqlJUaWNftP4qHAZA2tSQjx+cOhOr1+/3Fiy+4DRupcrd8MnF+K/paATRNsjHbGVhQ
9Tc5NhyTCZujMjBZWRru0ZkchyZEP4usjQUlDswGIWryckwyxyHfSAcD2L28f53sDKA0ZgRkzmQl
vdpcP87YMGYP+gSfZZXt2Fvdapl9vBT2tC+HSXy/oIdiawhInd6e/35i7nxdPd18UFtDKPc0XNm4
/SWMHJiyaJ643Fx9ct683WnTl6CNHu+Vq/iXtEKSmDJ/1865/r2aixxfyVda73a+P3R0O1Gppe5Q
UkrGBXutmQXu7qLhrRj9I41+6D6JnhXPanc9m90gLBFYWeZ/1FUO/SkJrfY5tX4RHPaXj7x0NKd0
iR40WP6rGpA7nG2H1Y4hj7RlwPugusYtHbrSji1pNv9vP0vuJSKIKhgxNEMC5+7VSLaJGGnAZXeg
T049MCtlaHYMFZGVyJDZlah00xNw4Ao7WVjIBS2qm96TdgLuznQoWOebLwp97qb/xZ+4hk0ut2+h
qZfdC3Sr+El3SHwK414emb7nW+5ql5d1ABLVf+JqAfvIAJiHJ3e85UGc/8yR/C8OdfIbpQrWnZd1
zuHdWYs0CnFkmlY4rJ9JZ2U6gMOOLtV4xVHVRcpZ3ZTMMTO8+o4oaP5kdnBU+/lxP7+Xua+BPkfV
5qilbt+Y65YZwmCQhXXn+lFoYR86piMvKD7Evi+HelL28H9bZLrN+hixNU5ANGJ7lMJI1TfdTmX0
0naJQxeHcuWhPMTwsIIHVh3i9iMUME51PeLIDZprAzzbmPzBmJko4CHrm55fjYydA4h29E0cx1WQ
9X5UKr7wOcZ5aJ83NJlbJKJiyfl3oagzpd+X/kR6AEJob2/T1Ha6ToKb0kWW/bmxBjNNu0bMHzSC
ve1DVFlaL+2v++u1QLtoTufDY08kGaW1lW916WmpKK9oAfXk3ToJtmKMuQFfa/rDW8HeWbahjXGG
4tLrySHnxGZ9viXdU7ePRAaW7Im/Owypsb7Vo+N4s8muLCU8twaHFvOGNs+k1HAl8aN1/3zpxbSR
45ve1fUiaop3ZDyB0OT7b1hF1vIC11AwuGv2LisTTyPw/FkEnbq7BEW8lZKOnK33feeksT1w7FIB
vr0BXJIy3YFBMoUXPLXqhP9vHTaTfG+TFQGdjQ7yaUxGirCvWGd4rLt5M5qx0hKk6+KVb+xa9GlC
ZREF88wbhC/E7G1yOeFikRcGzaIQ3rk98aRorfxZMqMCEr/xv/I5TF6MAMFP0DTvTzA//F2GGU/Y
325QK/aXfOPZjYgULavLXl/ybvfjTjHL8QFB4CfcwtzjSvGUNCQrNoi2YqNczNXpgSajWsMPAgSX
Ct/H9DxvpJnf/ViogI0hh81ZFPfgCBmluDONZwrsmgBoU2qyg/P6NJoS5EsUqQPL/4/sO48RzYpN
7fJdIfCoAFDBo5XGjksB8Qrbiv2hMto5FiJuXu4kmIA/a0/urPrpPwSWtP5ZcGmgHfWWgBe09bdj
qATVV0kEgq3dvlrudZW179npaO1VZiN/dBH/ELLIvR/N0IDMScf21LlVI2+DEun/0rE32/cZm9do
Q+eFksUhNjWBa6kzAVSJ+tW7vApmeOng4K/sPyIxTC5R0pocNJw+4GNzkhZci27Lvkh3dk5k9h6i
STopDNc9zQzNhRA7pdGb5cTY8OqS92sDU4ST63zJvNSQ2qH7Xpdbf1dnJhEE4Fx+b0K1tSTW62RU
4Eqyvbd80H94Got1R96dei6tdbSg1LFlgVoVDGLjPn8z2oUQWvI5kdkiqcGT14v/Ib+DiE2vU0dV
2wYp1XVy7EgSdXexFIiudl26WwvoRs2OSLI7Te3wz4oYQe0Vr7ZG90/vFFu5LNwzTO7QWIsRh2XQ
iziLWcymakweGSywqOuGrmfGzvaZGDg0/4AB7IGICI9z/0vUXf+mWdbdDCj07cvB0LYcCvW/Eq+5
YDXqxuxsfizU5vaGSkVzISXzw9yaxE8d7brS+EZMGU5TEyKBDfOc6j8dYujVf49rDF2ZtoQL47Jr
tBuS1McxqUm8ux5ZQ/MgDXlRCLS3iAMDutLlmKPNOYD9c8VguktT2Ymdm0IGHmDcznvDtlPElJ89
LpgY3Z8sz91aWqyHoUOAyXNBrRgIXpaj92SJ3pBR9YpH6GPmBUEPjdm8+iS8o02aPPsvJS1u7Wie
cvo/EuObkN6ue8uWvMfU9tMQK9itAS5h+lVoRrW4aHNPEfE7AeXzKUoQXrUUNUZk8FiOS3Q0qiFz
LNFbrNBcBn1OzEM+DxEW4MvpQmP8ZzD1fPfB3HLCH7eN2s2Tw5rNc6vhZMQAcOa3MnZfgOD4LA/4
7k5o2H/XkBY5hl59EPi7N/ytwMYjs9ZKD5WPS7X7k9vqFselERMBf4KAQCX7edx9pSiwZCQg4kpt
ZBzJCdGRaEaIWKMcFgqPMBI48iNdfDfUa1rcw9VbxKqYIG77ZIotRk4MzONxnBv9XObgsCoOCh3j
/svSNbdPA/Xvmr9ZN1eeeu2PJIHOdsuzs7lq6DzmQUQyhzV0RPG4+/FJ1qLQfHFBH4TVK3VnFN7d
NkG4UncgNXPTTmCHuOdtcoHvCojkWI5W07xIoA77DTsSUPNZee++B7DamO6psQXhSGTZ2QL0SYad
aQ1MWnU8+2nHsds/7tmUMgbO96ckxmzynqREsnVQHZKyY8XgZ4qCKnBj2bI5TmBjyVIEB0qtWGq/
7Qks7jILIDhLfXjYj3FFr3NkTz5XEFenE13Dx6NEt5lNJqPKXs+7qDrnKp4epbMFIEb8BeTi2QXu
dh2DVHtZeXm/F0Y4C4mWNteYaAJy2eMu3H+VWFMRf/axSJld/s2qgsXCKQt3NpjOLTuCKCHADrFV
RUAAF+VtgrcyWn6JaKKfLr3miPCLrP6P7ocp0DBTAK07dv+FNguE0My1b7FaVmg0+Cy6KaHlCuCf
2iJUKnifgNIxDcmBVTfAdNA1h09NaEX6kFA3+I8sqhAxdQNisOyhkI7IYIgMpecTTo+3J9Q3DB4X
5l/QNaojvjvzwshNc3i9Nc/so+BbZtfYghO/dMENZNZzmr6kyueJNo91fRpg/4m/gf1PRrj93Zsp
lnXzYCA92Ru5XhJ/ALOU2I3ApwVzXhFiQhBXE5acJlH/lSJrc1C7648vlffsqwJq3qxqhhdB88Q/
0my+CbzN5ZUzl8RhaFDO/FPUxOEsDEcr+X/EUMH2uS988K+W6Sj8Dcs6Z8an1Klk+rTpjytCNJjK
+15olRqEbn7yZXmtMensa3LTAq+zwl2CoqIy/FXFos72u78+/PtU5raQINg3xGxH8Ieq0dLCc+9s
oqlF3HK3nmkOzS3ff3gnwAAXtlQuED6cFF+kjqiP3maOWCRsNutl6tu2QFJTdrWHMLtPM3Fyf2AH
joIKdbAm5UT0wIz+1r44Fu/uYogohH9h2GTeHBG5NcoCaYbdlha8LEAs3Ofs5d4rTSaEnS0WWpKE
7NDd+MWkC8UNAXtFDS35yb3VUwUDNtbZH2YPulW06sRjAvmKncTvzlPsqehmdcrpJL4asijkSc2J
OStYw+3yztg2njeR8lyXFphUOaSUJ3Ute1WK0pub/wuKyF8gMDrttes8BYU44ZA2W/+vrhTL1yzF
7IfvJuaI1lC1xw+vYIaq3IhPuZlzHTMYRI/kXxrzeyB2n7I9VdlHJvOtNNkHVFiLcY4x62riAIoP
HaBLifYXinUEsI3Ml/ctDS9hE0/t1YmFuMbwy6z3dzWSot7DvZ+uSJczvN9089UVQIVY2DwYUpj9
0x93Z5OXeMtaxocdFm/dZmbamOITwjPHpSZURnXrHSq+PUSVWTOTMjZf0JgSgmp5rMS8bPDD+6sG
P/ezikTRgdtYs90uyh64X0dXMvvi+qGiYrQMWLPF2AzuhPRUgy4QsQ4ENFvPaf7zqsk9xYJLRx/c
WlgJF1xO8VM3tEajexRSINqNbhOnx7Kv5qU+ODxdS9vIOY+GmfKukzAS207RacFNMUW9cPXMCcTK
AShTbenidOmUS6q2jm3jmXtayVhRy5L+GUjaaaplcSlEebtOUYJY2dxcqsDf053jaJi30rVgJWPC
zidLT/30qaW7VRq7++ntEAHEZ8f5Bg2gfXGXQy2wbbKjpRJ54cgNyGvsdUkp468fu5QzkmEQjbon
vwdt/yQoz/z7+N8G+EhbmZ5iqAf0Qo4INng96tk3steQiaGhPk29Nqxq0xkYTjz0PKfizYJ2FfDF
TJ2d4xWZh4y9Bytmkg2UVgFykaT10WHsrUwOB28OOp+2GeHyyQDny7SUknJVYE2N8DLHJrJjz88R
KPfNei3l2FTrgdp1ci4xUxH/165EmcubdrRwzcvFHS3vC+sKvwPi8FvqSayw+wh/VcT2JEVX/299
naBWswqHyfaFJdyJeUSjXc0cqt2i1R+imSQxsmp/zIMzErgfmIkl4iuQRZDrve/PUeYf3iP3nJE8
oT6wzcTER+oNxHlSkAkY8WfR1NzvuhNeOkMNu7rl9WSC99gWZv+nMbA2YdmDFjImvL+C8P5uEJQr
iu3jynBB6FVoRqJMzzaen383JN2tgCHYeLBKSK0+6HlO+7lKuyRTRIMJ+hs0GnBQQH2YhG+FxSa1
7w/Mc6/ymkbXUiaG9jmQGMoynE6cfNbf6a2tPuJaCCd5A9vaQmWUtvFopsBiH/wPJSV/7l7kDK3m
at0XNAdyzS3l08JwQkra1J4UcsBGz2hTlNZan1vsqhgHJj6gUuYYiaMWy9TPewG2Wmrs/VFxk352
7u4FSCrS0TGb/yJ5yVe/8GYkKVPE+sug3m4SK6f5yH3m7KvCzI5xgOGYdHJWJ/vU7bXXlB/zgpZk
IVRAiNsEbGgQdXKK1bFKd4nxh0DkzAgSawcMbTpXzMDcXuhSPCKcdqKQRu3o2qgbehWH8F6fAtjn
33indaKkRmJalDDhVC3BLy2PC9i6s6R4oLNFgGguEe+SbEXObzdXFu/nno6scuFQxKIyr7PO8Ef/
vBBRkwJuC+xMYhMKX/r44Px+Z/aF9bzlqfJwKXrwFlg5qDfGHJFdRe1ZIUsU50I0jRtvAoDkzspV
20tqzoAmtBuhbPxPRXwOKrA+2QMkPWEnH5YYlQDi/TefodFIWGU03VQV2e2x9x5WqPfFwZCuu8m+
6YL2nW/dHZi3fp4cS20PmepIEpEK2pqpzJ0+xWwUK4nUyYELz3xdn0+yF00TDmZeifL/KO/1NJvw
UqHfyPohnTnBDeUyg+NDSAAQgM5f4YaYcUNwC26OvGNbIUAcZTzyqjtJZaE53xP0L7bfl09nFiky
IlIMam9O+p5Zin1RuWJkkHq9mwTE+XD9fBJ/FwGCJYJMbg++DO1qonQALNJX1L4eKHWbkC630++z
0S+Bu6GyOdmS9obRuUSN/zhBSgV6sMXBq7Lz6Pm76pvaq/EHy2BJ9jKraJFM8uAxN5iinEHyO5rp
ElIWXNUe5BQHLcUnD+Fj+vLw44tTCygGWdbESYDy8FVvM6isUOl7mu664cTToCg4BWz6Nzr6cH6+
/hkGJx+L8LaIAMtLVz3I1MYzgUTlsN6GWi0Ik07TlzXVhIoWf9xthQ7m14SIAnnbL0MSWv5cmKwN
PHUwfaUoE9AZnkUDWosWCRhVvquQdpibzw/YTum5+httGd5uyIHpxmRc7M687LjLaGufUWSzobu1
4XKNieAfu/B6r1ZPiK/DP42z4aiOG3mDxQal8Y/67//ug8iHCB6VeUFrqb0IJ2QSse00p1bJWjIE
rtHAx3bSh8pOMjqOc0u5wDscUBi8KUgWwVkIUQ5a7KH01v5GlUPd4ndZyl4vvpk8mT3t3SLkAQnD
Lw/E+C3H9q/BMBmwzHPPADoCIb+oPNP5x2Y5oLJxLeuFKcpeKCUUkCMht0ItO425zTPvswL/bDWx
SiUyKonEfbnSnmowzQ+nD27LRYgzPyFddoQ7wHRzpTyNf9pGj6tOm0lJVed7Z4DHUcsTstq3VgX8
50b7IxSXeCBjE+I3aMSW/PV9HgrZ6qSxrgnsz1i2eGSXUN3AfNoMDESba77UdNvKZZWTstXLoPKJ
f9jzup/P+wG0SFr+9+AYqenBGtUAnv6LqlH6ufHCfYAXh46G+Dtdco78NnlLNSNmq12UIi4ROlta
2pRp3YcbHv7BAwbbmo2HibxOktaMKEpRcyNUoK+rSYuSU962JdYH3YV84qHOUPR4a+GpPQe5GTbj
D3T5JLw2G1i2Tbq+PtZh/ttG8tyo5QlLRMmmYbbpBMmpHkIy6peFflKgTtu4bpkQQ6AAObFVLqDv
N/Aecm9zCrJ07O+FCp8HL3ZQMDSgI5B/a1yTOZVs3NYjcfCH2Wv/PAssb/JVScME6Z5IxNxEj0ej
j/ChD+/3g2G4ECJsME2KQpMoQXFEy401clHP0DWtI5bnQde+CMgfJ1zCg0uzodFTeh/jNgn84V2Z
GBxtpjlFqpwZPJnTgH8b45jLm0lfRDCM2fOEbevvmeHUAiQjQDF+lrb5cCQZhEhoblvf6panZX1q
0AZ2Ou0zAHLzRNb4yEX8yG07tH3tt1koTSuh09KneOkblNWRdFlD8pVEl1m05gLIRNdEtms856GE
SYss1eKrXWHJk11u0BO7osXYhuvYSEnPEb/eK298Bqu1hPDNbVSloDq4mEEI5/+rTvLwJlfKheEi
d0bEmXNs7H50MEc0J0IFxBaRFdTJhQxn+uKSqsgOjlY6LiXCvMHIkea35bmIRMAmljMOGGb416hn
FpAnI8oCUVU2XRSi9bw8LMHtwxeIKnj8cqyfLh4ahhJt/8Sg3aV235o3PL5nJM96I+GJR9WMoPVB
fDTJ4bmhOTNCafpYP/QP1MXdMz0qwoNbfAR7lMbXpp4uWVIW/kHrymy7sSWu+ym/u2VP4gpvW1ps
8lgucFbbNQElest4aCzElaJefMasgqsG5+Q3NVujn5iJ/7Wdj9Xg8HHyAaKtmJBmg3YWVMAaLrJL
7/IFLMuentM/6ALTsZ+GHQPX6Uq/JAH+UkvgTfIO29HyHCrxYkPq46RyTDVMhM01pkQJjDGtJZar
y3DrqKZmiKSltnJ1k5m01Uw9HnBm2J7N4RqFUNEWEhLW9QHBpkU5EaGXG5Wpv9v2pgUK0H3nFJAT
bOjORQIbzbjG0rEB3wVGznuFRDplIA8MT8PxxTBhDprXy+/ZclPh5wV2Df/1vjGkIhhRSgGtdzLQ
0jqzErZ+/9uE4owh2Wnnfn1dHMO7h4EBiJiiJYPbvS1YHpPo8qLweE7HifMEQ1yfSok6fZE25Z0q
A/9KnQQeVobFcv+Ek0k8jGLf0dVllpCJpxBimVCbCSn3x4pDSzoT/7BhK0hwUrrNSozb7toCCTvq
YXPQXW2ugSN1HWp+0u7MYtP5rmYB7K4a4s23WREYQJSlhp2q5mrFbcj9iW/wmWnePfaYpRlJISJy
UqVgS5sJmW6hfO8yDH0CIq/Xn9QLb/I5h9wgP/2GfV2GOnxZiFsqTNTHFnFFXabKdjjuyxebJqkH
CKzcjDvof87VyQyJFdMsOBYrIyGrPgoRY94ggrTrGecvdZteXpH/kqp3ThmzZLgBrVA7twPDjrNB
VEyPwcbfTrF16iyDy+fAE48GmTdHx056edMh0x/AQmvoefUfslHwXNnJfH7gxqmlRXbxKb3FNmsf
Yo/Lwq4a/sDd27r2UNjSsgZYHPkOeFTF4ZNuqs1sDMbXTD9qUG1JPm0D+rW2KVED0M310f/kRCZy
Z8ITqLyGFts6pU0XS4nTH848dHFc/lz3tjkN2IR8CTqr6CmQR8iqM5R26fstj1t/pmx1DUOrYiRZ
bsLgsSBzOxFFfB3mzXAPySQbZ0vDBTLjSS+LPAwl+TGkCuR08XaJcLDkh3GQKHxaEiR0+aXvDtwy
hkBOqMPzuhXWQxpIKxBx6HURmjXO6VxwFuPws3GRMea+1wrXrwMw24gjbKcvzr9O+Jn88n+xQ2iD
fUC1eh5fYn/hL8n1Lfd2peTi43zDvNspPJihJ0QuV0zqZuuDJdO3wt8atbOgfvJe9wNzI1ieY3+W
HtuipBA36ba20BM9jpeKlzkzVNADbJlvjKDG7n72MfFFF+u4lDJfppoR0FfmuE5A9icZt0yjrhXI
JiVFSHawUuEfcNYukx/LcrQrgaLYgja7kW+ZGPxnfgE/UqPOvrQZWq+q8hmXO0QKXNdsxBJNsNU+
XGGyhpULE41HeGaKFmcuKDH+fGW6Hom+PDJW1udncWltIpxKQ/w8nrtwf+Uov/foNwhbD3doPjmM
0iY4KDrjQViG5GvRH7p72mChzI3oAn8umDRIvpZ5SMA93TGMVOQuZR9Lo4XlPdITjhqn4QiEw/RM
hLNAfBeSQCphRjweHnsG+11XHPe5CnzzQ3RIzqjFmdrvKKYVb4zd6QYAEjaiFKyQT4JgEKRqLmIc
AbxAytL4m/EV2klWlSv8G2zToB5FhDAcKwBBT2JAja4vAL74Kr9oG5vewCEjmE3p2mNk/aVFs1T4
9S9uk+RyEHQ0CLnE7wWpDR0LFei7tAtczfW6+C8+3jN11rc5vnFghu2OdIy2peqKQ0kW1O8iJt0T
r4A1Z2AJ1XCaAhVYbjsmKHyc5qzswgSZyOdpNP5uL1qANGaZWbhpS6WYvCOaLxGIBP68tnDapSOv
QYWymn2IRLeZrNUxJmzzlq7On3D6eSMZU0HVz0LY87QI9wXwGzj1MyajRqjKjhxN5SaDqrdHkBw5
6oKSy1NR3QDopA2FTSxuoiVkOVJ9vb++Xp1t1NiYecvHZR6VHKrGNh+4wbnUfKmVhn1Tr1Psh6vW
z4hO0BuhIFbDp6HCN8DrrzV124+KxZ2/JYsHmDIwL/I2mYVH9WY2ZQFYh627pO+lZlSqoY1mIRXx
ZslhtuA/ovc+wZiSOdEEAunG3YTWr6ySHmLf4HpvPYDmvq3k1fi+YixfBZ5cQ4Pbd0DFQZ2qCAGj
nJJqvH6D09UsELEBqueUvkbnbaL/f4fyXlZs8LFI1i/ZeeJbRwDO0NWYc/LSaDaV2TiRWmmjlGWC
an6gztj+JFY/XjOyEztng29Pl0od7PUjBoWwwG8ihkqXBq/fbRVWoCRVAtRyTC5JJHSgqpgXbPMQ
S1iKJqnwkSqCozoe9q1xFgBb0Nq9VXwGeASlARSbyPvMR7KWcX6EppH79J4eOHxNDCMu2UeYTiJy
WBZl31si/rbfYyxHTZmmVUVlMIDsdp4TqF1PWm3OvGYrJ/nEKY+hYT9ZTGKN27aQvANH6XhdONWv
3uTtkTMLtZn8A+31Wn2krKy3MSoi6LBjBoMH4U8bEetm6dZo6Xq9bTN3C+Bc9exH70cQYM9+dXlf
OmN/A29zNqhuHDvbVF7W0uQqTgJIxvvH7HLrXFMclhp7Qqh7fnJROfXy9WtLDhEmZI89AAmtLr4+
wOf1GNC5pK7bGE/GCv8DSYf/YJpgQJ94x7L4uC6c63JmGE6RN/hkzLhzjtpjVA/I2PSZuDGHmXye
gquBhT06JNeEvZFUwv1ZszgGTP50CMRr7tpJFzauPY5jx53A/FIOiiujmnCvg44tOxUrdgEIdDBq
L/FcV1Bn3LX0lD4CAq4kLAVF8/QLiK2au9gmfqVWmtYKR3jKzcvhbs1+T7/pgGyxyJD0Fl0E4MC8
NWZxP7w7SZ8xSfg8ttcy0Q5mMws9J8gZnWJst+wErDRdjAsT1Gjt1vKChPZHyzfgVsHWWwNptGWa
+Za33RvmP8ygyFkAG2jzdVpnylNRKWMcvj/92BxV2x+QJt6ZfjJoIl/5NCm05LNXjLUPdRMmBGwW
/0fg/Mh+JWa9eeu/fSJzKObDngnKTU2S3Hn9DlVdJUFYybvqfZ3fjzK3/lirvqrSq4hgkQAWy54/
huqbr08rATfW1ryIElS5tUGnC7s1C/C0GFayDL4q6YH8wbb82XAQbWm7Bx8xn4PYj22NgCH76C39
SAlTLWuynPxKfmeJBOLzwtQNZOO0fcGzv9z50RcCzYGOqAdFoc1pU/3E9qiFTGArhlSyPGS2ZZiC
L5QXRUC9BLiGOGiABfK9pkN9fkxwSZ5dIf0da2AKYX3HkZxVF4I2x9lnU4j6/kOrPPGHx/mw2fQZ
yPIoJ/KQprsj3pIlwsE+IPzLCyu4JkCX+ZdAkAuTNtCH04CJdQK00tv09SFoQE8ArZmerSrq9pFX
8iDc1l9O3jUyWq6FRI+8ggXN1dsm+PP+VeRGIF9Rj0mH1IAjhERpLPL1XPBDOgqzyTKLayL2Xh74
Wg8TOI03/v644wE1oK5BirLZuMBrWr0wmmxWU73vJDcv2vJrzpW5Qj5eEEbz8cnflil1IfpwxjTZ
TxzidBy17yOwwOIuYmmyQkLCm5m+XcIJyTuiQ+b9ukx6jaQfiuUUU+2PZVuU0WoCHhXS38S7S+lj
xIztarAO/jvd4vmszqNJBlmkSy9DEg4ThzKntz3B9QtKob8O57oUqfHLlk2XjA8HZzibHd8RrdBy
U+VnHyY/kQOGl3/5Ko7BYWt9seXn2KUvPf1c+Gl4+lIEB6iguXo9w9TM/gs3GYQvOeAUIaX8ULmH
qMlzrSkkuP2L98w8AWEeaP1VAzQuvYyGe3szTPSWsIf6wAx+4isHaIWkgdMY/0uyBZciSBMtW8+U
tzokbcoY9g00wpJ8kpc7+VfAbfA27z+Zbd8XDehJn5vOeuSlKMalbHLkhxOsgFEeMDOEWs7Bz3yS
Cl9NAKB8ppgwrv83abGtfKMoDYGm7NfAxO445tlwM45ZdXMnuaQHdAVgHFEJCV8qXgU5lhajV7YN
QtAb1hlqTdYSbPZqw10cPoFlbFO9W/5T+GN4tm7Y7PZlZUuljjOeBI3ezeMU0J63LFnqO3Wv1sid
xMF2L8J9VgF8mbJPhl0cFPo3sLl43FCxlzNFtJlIU2K5BaoiVPpDTBswrNMREQZcqe8Py4R92+KT
yo8ZH46zm/Jvw8tiEn3Ig3A1q6qlua5DquH3zqgXCXFv1+wOgQ00Yw7pbMIn3AflL306SgchOx0e
ArXPL6Oz/Nj2NwMdGCWQ7l7WyPx/JDQYbaZfI13+TlyM+GqZcUlBBRWh/oCOAnFY9qzMuCVjqD7C
4kMj2uI+S+gYw7ABqxCy5lt8wqqASIhebOtfXgf4raj+8l2fqz+uyewWKDXnD/zxyuFi/AQA77ij
rowHRun4P1Zr6qLWPAYP+dkRrHG6ijAAeI2Yjth/qpPg8KdPLLTyg50YEPdhjbTdtHTt8qmL+wL5
n/yoS5v29mAVGP83Wi2prvS/nA0CWmNC02qHFFjebmQgC04WCNmi6asDcF3r0UvUO2Z0pqqpW/KK
Hn+GH7u0HlwtDCj4YbLp/j1HFM0xcT0q1i+PycVbvUA7xgfSjb0ZO65PTiXsEn85ZpnUP/diHsX7
SCFIW+WMwa3njv6fbp2twcaAEk/WdV3/11pYJj8B5KyszFqxBE2wJdP8c9ud9neIFsH9xqGZiElh
Lj2hElOCSgMkqVA5GRflI0+4fkQdIntbub51mXGMnn3woysrFGMQtuARavJd8uaxm+639IocimVU
kLDofFI2I1TIpx/Y35eWeOAU4Loe7JKJaozqdBllWZUOcR/q3QGqPIPg7VhjNdtdpJW5L3eRM+PO
10g/rGBdcN+LLAnJ84ZRT9tbOqVaVD5tjOSBN2JifTSjieZu8SivEZctJyp/xjmJMPvsJxJZ4EA8
sPwA19OjE9ZNT/VnJbfxp9n25sLfsnmYWdnmIHJVVGHoaV5Vo2x9L+mg5xPQg4HJUozu/g7Rlrra
S9PYGW/8j2Iy5+T4HYgtnLk4SfkmjgrEaAGJWZ/9htoOdbiH2cb0RaW6JOd3QshFQet5MJU5Q3B/
trQBT783qiHOuJBW6W6f7juuNvwEey3VH1NBYIteto+/oIlncVF8PbXxuGPnfvkJaF0ZgzWuDoK/
s+oxYZRO/NPXswBK+x58kShsEsHPN3Pmin7gVD3tM9BaOLc2nlebI4WjilUiUMRWqRlefzpGJAbl
ygXlj/cdUbezrBw5tcFb0ic5EfdcGcC+NNaK6EFxGlOoXrwGD3fb8zEjbrZgCiJ8l2Dh9aHxwOKB
cNqOVL0pjoZRbM7CskyWEBgEH3Px0yaKITAUSk2VEYTK3wHP2MxvEXbawDpChncROZzId9sWzqhR
KdoRLssVBz5cdxrsjBXfmwhMbdBikhkZZLTEOccTZFs4oL2KqZ+kPMT0nMG+7kpXU7FIG/KAjnUW
o/YW+ibx7KTtWIgL/SPbZzwb3l6C7qRsQ966j9yR31tqTOk+JJnBdIocjYG7tVEyeupD4lGX6OjG
Sx/LrWTkNQf7orWZ77DNHcLaWcAmV2U/YKrkblhSdIIcVbdO4Z6gn5a2BJGgSB3a4VyyErCuoOCO
XEZ+K+BpAGAvGJ9yH7c7gXu+zR4giBV+JUkD/AtSu1OnZAXtkcbORGimr/C/5DK8Ql6uU+/6i4kr
wvVDf7cS1MsOmN5jzYnDdKjjUCjd00LI6ghNAj099yqm+p4vt4vYAOyVhOua8Y/Tu7/ls9hubWUw
+eQJqrykqCNp27GWlUfCtKQS2hHeO/0qNm627Bv2mH/rN/BhthogSGo7QzS8Aq4tM0BHlYa7kayX
INFTRDUa/a0rOzwmuP3xN92vNTt2n4kzxM67NWDrvkzw6OpB49DdxYTALyf33B6j3hC9TdP62IZk
BuCe9ANRSrUyStBdXmuEaNp/GRp/vPJPMAb/baeYM5cXzHbJTxnVpOCAK8ClL1/JL3GPuBc1NTfD
63hCJiOf4iOCpJe74B1gVMXm4+9VC3f2Rt+udrNcylj9djYOWBKEsRtmopYpA1rWkaRHHS7oaDyf
FOfvu1J+Y0ginbq/3OQLxxbMLHPUKA9X+RBSYUUM0Ac5iwFeSm2GA16w34s2fTFGe4dOwrjqxNez
GciDnZhWft5PD8cNooAMPCsvY9fzgXa06HmrEdgCkkm5HpvdWP8Ogo7iO10Bqe+giReSdAGJ+BWV
UY9Fp2Lls/3E/TTXj5YLixBrrt0SlwCjWAfRGHH4+NvoPF9gmEfafhQUKRS1VRZDFZNjDF1F1hIL
nhFH0cKzQNozRvULmdwYvSCDAc7phQbu7EkWMWZT+dBxACbzi3vJZTVLaZAR+XV/k1tCN0mcSKhE
90EPGOfWIAZRcLMabxSNb3ADihVrOxT4x2Ah7yH+bEaoDP/7+BmU4hYLwBpjoch4ZzkdNvzAujNQ
upeDUyULQDwZD1iyX4z5hsXWLJIRepBBAcb6q9nNv1Ps/LOnS5zGtUiOcbbru9NG9PANgIKUBDFL
IhyrkKpsgDJtfwubzlO3TWF4AYM5XerKQJ+afOlrdLgHFzlzewsxWCuJ5v10wUFP2j436tENte8W
YZJGPwYBiK2wJbryXKQ2ILp0QaU6C7Lu2oiUZUxl7j+5ESqcNmcGffEdv2EjKmLTfXcYTxMpOG6F
44cul2b+3Bl3+tqT3mNY2oKqqw8+agyMxMHseceSrlOYDDU5I9PeR6TX9Fm4GD/chVNknbIIo4ow
Ri21mTCez0J8DY4yad0OEU0iyPmOXH5Do+UIVqBZGL02jjwuZMbq7McC9vCKItb+dU0p01M/liH9
LIO+5pBw80TYG1pSTiLCejhJZNbIXcNfn3nNkkX03O57rdajaOrkWKJneuIoKrxvacw043cQXbR8
Xg8DtoSL0XUZj9LpmrUrAmLSx8V/JKI341drWdAuNdiWfy52ZzKyK/HNwnDM9ms8dzqQtdnrWye1
EdcDWUPKPWdmq5LRHscItVXP53VLGP6VblSR/YPsiKdxUo/RoP1X7FQEqUJcEl6aPIM9s6xjQQIu
6BN5HdY5LCMaSZfRiboP/Pt91KJfdEc0/q2jCR/Q15Wy8CeWU4iwiG7K6s4AAd8ayrS2hMQeiYJ6
mkG8/LXkzXmUM/IjCNQMFCCWRHlUA2K3IYnoZKNg2VpM5L1wKmzgUcIv4qZRQtxgVA1t2FZvLqsg
u6uu0Rt5l5RUiaZ+QEMwkavhPGo2Zcxnx2pGASwPwU6Jy8f/JSKy7sfBoFEDWbr0HheJrfk2I2z4
T3SOLy55Cfm6Lrijy2QdCYOtnFB1Duy2Tr6PvoVsrQyz/vo0o6vrlJBTTnf0P8f4ugzonRMM6jCO
bqZ/v43qFuST1ohQ5oGEvTNMVAnGQr0cU4iZ1xqWEQkoJ7lDV1gUZumriIG6WFWW/TS6j18mNMCB
ImyvlKvyv5ZOqdJoZCQd3cgdrVDTqsmi3p19xH41ItoijLjf9utUBjlPa8IuqhNWSU927/lu5jiv
1bDbgiXXSQrQflr3j6uekFp76wi5yVlBNUdSc6t6kY/z8ANEqDcspDkDKYbF6cv19zRRbqlAJQy8
JYleKxtLyvkQWSOgZ1IgOeQIU24YURBMacfNfuTe1o9WMLPSOpIC4/NXkIXBDzmXETnRvJhrL8HW
yTG45KNOAIzSxbkGWc3zdWhVdzR4FN3rqTfhj9cLvDBK8Jdj8azoJP7v1T7svGNqvxDfWYNDkDrk
VCxivy+/WGuX+YpjflcE+yAiTOJ549laeGYaYeQsaIvNDGAnW4HYXDqywV2PEcjbggGZxXYj8iD+
bEUuidqtFGOAYVtZ2cKVxu3n0ee7NkQKh5LlBVD1l3oPPnhJs+vh6qWfZcfaFpZdnoL27ckBIYiu
I9yVhZspSRt8qpEOMfb56kBTManayXpf23+D8k3/VmivQ6CxMYjJOXnvnB/U3W8d0G+z4Ac9OBxP
zh578CDC4RXOdyJtqkRUqqq07vMsLE/guVL0vKXvEqAv3VYELuTNVDPY4WJNSFm0gp5+Q6Te/263
wcb8Jcc68TkV2zzswdoLBfVNEM4DT3n1PTza0BBq0GFxPpmv4xx8JvUwTPMGLy1B+Jbx4d7VOKq1
uZ5sVaeJGU7jfGtkTBk13LB8dCIXJsUtUt3pnHpsizrhUhjX8srHGssdK0y4bx2fvGOgn0Vuhqpq
uSMeQ0ek2WZB4BkfVzNBZCX5HHe/vecYIEqfdj1jbx2I5t1UJwr9tekrPo3iFBtGnf92eFYGCjmO
DgRzDVaQ/qpKMANag7PxRzk3QxhLKZOZ7+2ILADHDHGPRSrCsUjh7thwprVsnHKxXt3f5ODfxkdf
cAfjR5dARzrMnpYTseqKQz42h8Q+9/fIEIE5EhSrC+mhFHMq3Pxqg9/7e6swdMXp6tPJm8L1sjip
PrtGpstbE4goGFiSyWSRPE5TbSnyNV+3eOia00zuKpbr45r4sXMnJUJr5UxyInqYMClA+lBRP6tx
KFxwdqH6ofG0CQKO4+95vYfSxOmMraVrKM+qR6mkZHn8zx+KhEkcOXDoFBWeibXNV+LwZaqXqVDd
MdnuOA4lblrWrPU7DImDx3qXM47fVwZXW5c7/Q0GfNqucfkGeuceHtI7Ba8Rfx+JtK29gCy5X9PH
tazpi3YmgKi4Px3tgTM7lKfVdu9P2sfCUkIXCzK/DLHiJ+ymFLe4Rbx/RzO1fkop+m6HT+cbPtQh
uyU7YEnjVwRt2Kaa1T9uLvoKSxZrWp8Sid5pNMWi+HmrFUODUUj46OGUDo0UhU9IeOaeQSkuQLMC
udbp3LMQdeeqjO8qHLnZudUsu8CLr1i1CBtFnhJGTtqb7V/NDGHlrv0iLhUi/7E0/KYXKhtp3Nx2
dcsdvO4hn0RTLzefPRWGwDSvc109rVIt0yS86Dpt6JhK46HpIn0FlF6uLEqsT3/RoqOfA039P+a6
BdhuHspj6wrdlTlgVdmOVQzweUxyjcm+BBWiRs0hlK4sMNNA9SnHx6buZKiMujZgMR4i4EN7yueL
yiXsY73Lf78zpomH0Bkx7gTWKqb3F4cXeb7AeoEf0DuKUy0ydyA58IuV6nP/NIM/SLT+5BZOEbJM
VTGYiYOAbf6cUombWZvltaGBLnWzr1rqm9xBuc8WJlb0BNzcdxM6ZUnjD4J78yLurHfiPkXBsFIJ
yV5ai5bRemsMcsrFC56kTps/GGjBJcDkY6s66cT9kSdvS6gCT3jOKenI7TKJIvz4WfNrlDshDEqa
MTdOlR9v/hn2rGQdIavXo97wUYfFc2Eo4HqyUhLpdDt3gAHuNVrQET6RZAdA+avXpnqzE8l6rcVs
cd0J+pAVnQiWopWpBp/tqieIgi96/JuXnoIxKpMFRuroYy9jtonoxqoZ48TadGtjG5do7yvdYSqU
+1iTMkxb2cKap8FSehlj8YT7GKYlmN80NQs3X+qoPscIy7MgnhsHjrefLvd5i5jB4sTYb5lJ//9T
GI2DDZeR8xkS/T0naQWLAhM70Ln9jm0h0sbd2tJB/G+ZhtOAM9cs6EpoX11idMQptT0XHU4L8OTH
Y09M9Tgi0TCG/+90g+gIseWPE1Nvl/n32KyS0VUkwOuV6mkL9rwVm/9itL+GdT2prtba744lGJwR
Qkk8/M+eh6KvPjMQa7cllPYTy9GHwzXyKdkNe6CJf2fjwwxz+eUcim9EbcuzBF3usZzaJn1Luwlg
dN2ip8qiDvlKTWWa5DBMTvYYjEv5jwSYIxKntycMjsrDSfiVmw3C/Q0h9BAcXYJzt0Z/SDOP4qXq
pdj6ZizzH4GOUdj3vbr3eB39LimAXUyntG52vtvttGi5UmpV7cO9l3tLsGVeOX0M6B+SIOygJpis
hS/Lq+pca7m9/e1GMf5I+7oN2nsg3FG0Y+rjNOJfjVGxJt+9Ou8crRuQi9IiooPSwoEKfIO07uG2
0HI4+t93knRQUfjVpbzJW3vMbGPPrE7+Xq5ktebLTaT88hZYwfAjsYAeSKgiuT79zTAl/n4RDXEu
ekLOpl7cAokNIhvhs1c7vb+EHVGOEoMkXjVZbs6pvcpg71447rgSQmOlJzyjNvVxy8WR8TsNwaT/
0M0kUhqqpdhemWOMXEwoq5XZpKPMRxVchKsCX4a8J1dmaoI764oSS9Hh0WW7KBqAvrQbapFjd2AO
coFovXcBXwPzuy+p7F1Bx9e5M8u6zH6B5E4J30VCxR0YgWihbCuDfZ7qg9TyLMmIbpRLjqGTrE22
3aYqdkjCX4yygu1TFVi/G7u2KXkD98401Bmgf9FvfAA0dZnyBknb1M/Ft6PxDYFyGwBnaUNQIoyG
RF8c6lwl7QrnvcU1BWnvV3jiJiq2XQfQzHCGDC8l3KzCas2N4qS4cR7Mx+rhfD6CUTU1db0I+wnu
fyJyjE+277J5mNxoN30vv6rvYKrMGVl0ZuYNm5LrIEotZJ+t22TgbTQqcqKSn8B4+dQsVxCLpmNJ
EZFDmQrVFLBY1IVw8ifVmZ+czxZMqKJwaJ7TZM6cJrcuK7I4SHsyERW7MKeyCzO3AuInK4rerq0g
SbPCbWjEBimGzWzcHCSWScSHxZQUncQYZOC6jktGa7zjEh9N18BwOKxS+EUlxF4gTkTSt/GRfWl7
U98bu6ZeGu+edsH2JEBaoFebV5tKSCvZVDmWbwQ+hH0LW2D5lDUb1KKA6BfRy97i4tqnBMaNOclp
5z+Lz3Su+tJjKhhGgTJu0gQf/qcENPAVL3rmwXiiAzn40GTCxcMsfWhdr7dwkjpVjb9t8xIrimHC
BRkjNtHLhUnQPSCtOkjGt6GdbIa9Wu18yjKjymwUKMC7nWDj0Rhq8GsQcZ4b/cskn0pMhqcsC7+r
JbJH3rSod666bYPlBZiiYcE4JRvNZz8aDg6C0NAd51H2aB5KqmTfiHFrNG0a00Z8L8H39cZKlv+v
eJBeqpwXVwXyhn4VJfvNo4PY4IPErwkHXU3vqCkHnlwC8xJwtj3XhJ2iq+1+2MWZj65KJ6f5zFnZ
/itAspnyyynZ5VEfi1y4i+UsTkqGoIO/E5pvWZ6F6nRDxlT0prV8pdqNPr/6lz98WrXAeV750SxR
ZayWsO4LKcrG6HEpy3egaKVoDOMbRTIoScL6oFl2swaoZNyF6M06ie19F6KFfJ2wONwXHYzeEi6y
QOMWxQubXClgfCvyjhvm7nSDCA3VnvcWEQiC6Cyfex4isIXOztNOg1ZskjHgjYiZmfDI+zJViS9i
8l28Y0+wb21gnf9yTmWyw4Iu1aJgEjBekCmldFgFcLLccZXpeoSaFi9Qh2PRF1lMngZbsypuMjhI
UBibDS4ozbblnQl48nyfDbpQnd/viGdyKYiDBwS562a/pTcg2iIadma+ag4NNfeThsMLSqaZazrY
YToHoVuEhfDw/humOHAhojSHPKbI8wg9FwhLQMD1pZVzzSeDYhFfcjFGViTCRnTV2DfJ2lxahy/G
JSZ9xdzwqZk4rdTRgCaYvUlpT5C720i6YC+rR0zxjyZN7VW6Uz9Z/qbSuHXPNOsKwunABgYbbIys
KRV1D0aFdWuT7jX9GTKKST+MyLEVUW/iLsFXDpiWYWyqgsFC1602VnEL3oDYsOcq6lw1ktN4yyGc
P/hyZdaG3rClzbVCOVSkIkWXg6+fwQ5/TN0qSXYxW73HtVFXhEiURe2e0lhGN9AKjoNmTqS+t1FJ
iBguFs2O/e3XYM7j/wZdFCqMjtFdBeyCek3fSuaFwD9Aj0Khg2LARHIwALe+b60pVWlmSulePnjc
KKkFQr89mPrWwywX5Erln3FBbLlSGT0eQp+kXaQCuEb32kXinhZA1ToztFcEWlvJhTj48hibFi87
crwILftdmjJaDkA6tMthL156CcgHmyJOBrpM7Qo+N7Caiz8h8AE4CI87IB0gVIYLGobePypJji2v
PuyFpkA4q8mGc03sWc8tS8Zln/knrL6lYMybiVixzRs/EikhpknbhIzaNdaid54q1y7WH3iRHyqm
o19ZA1cUw3XVykilEI8/p4opFHlGlOrX+L6fJGCKBN+JHEuBFS6E255LS1c6JFNnaErGwqbla45u
8U7H7lah8CBkieGg07JJYDX21UZQeZXUDOn/3TaZIHojV6/WSguhPinpPJLszDCO0XbmyKZvKVDl
dbbekUAhTqxC5tDsVJ+P/oQvXQXV7MRdnRQGg6kUigaVIvBmhcYfMOQ6jiG5/DYaMNohyCK7N1Q/
d176HuXl6FHMAhmiKcMOBWSj7AhDK25IDnJve9lB/QSCLQ2qviHZCbTv46wselB/9CGypHlOBdY2
m12CWIsYzrcK5FXt27FxONIyvzSZlL05K1N1kfLmDA8X6PN5omC1h0oSeoQSkdDz9xmAnEx9ZGR3
zkQjPDbymq+mJzT9Syv808TgAj5mER4MZMNu0HaqyOY6s4DZyYK7cUwM4d1WyV5obyBFmhwKRUY5
oanbOe6WRm+94HQPpiRxSaE5wW0sj/KjJF5uLaMQ5rWlilzOhQjE6j3m+NI/5Fom7WchWM8j2qtB
v9WN4EX3k6pFEn5XTwJ6qZk0D8MS1DKSiopgOCphaDryNZObMgtuJtRSa/OfrpU1kzyMOxcyaBf3
SG4qJfII6LQvqQ2FK+1vx36rXQfbiAKPVHK+v8EN3NlOAhbjmG6jwb3vR56T4E1aRsCkty2MoR41
O8mXWJmc1ee+riU/kVELb6L3SnaY9oaOm/dQ68TCpNVfrGPAAOeFZ3vq0WtdypQo0oiBUJVPt7zD
fSNmh9zlZWf7jWrI6Cs5eilvo4TNv2BFSeIrshas58COmDp/HsepY3ulUM88W6+3ImkT/eZZaRKc
LImClbiMHgBWDGtoTr35OsUXJvQzqXz3YxJRyO/JbLWkDhMp3a+hEOX9YbBWaaWWRlbEZGMPRldI
EMMsNqH9vo9HOIgfOc49M3+uF7kDmKkMhz8rV3qzdui+bo2GWtMSk3xFVmO2rvM1Zo9+wRj96ziw
z/oXmSslqjbl2YRh3pSInpw2h/EWk90bo2f3nyOQSUxfYC8AOZe4XRIZl5+xKzDQ5x79E2neStzG
/3Z9kOAdUxRFFoEbcvcIk0+k8HL/Y6VlRcj1oFaG4QMM8g7JvVOGRDItyRXVVJnbggqd+TeMk+VQ
+GuG+PNghZvGBXMvX9q9DQWJlw4bH0EFwSYy1ORJ+eIN5NjN1xAh+IAdlKr4lOygqCQ5i5Vn7n9v
apSOAo3x8mPky6UbB+YfhHrqGDPmj0smZl167JcPyIVNPR2ZC0LF6TqdPtHNeYWYq5pjRFjN8ViM
DNoFXQucaMpRhcCA2fGDh3o2oEdyecK7Y+/CiadmhoWCFpNzxApEsw9O6uLXOd4wjwxKJwFHLvmw
uA1kb2YXlxGypNFpCT2cYOF3t0NI9/CZxpqcAlDaS3SRSPQiWSGxNWbplrx5CodhXSuDnSRvYx1s
5fiQFvUPA0qnU3Lfx/vqsMZdUoLTNsCGtynYIeArC7LT0rBJN31xvJ6V/YSuci38/QuhVzC7sUjc
mp9XGZuxKvzXIswrFNLMtqUO3kn+WViSmTScT7gObYwn0N4k/4BBGJLaTWce+MFmzBw8oC4R/7G5
XSofqRiRr4DIcQij7otAohuo4awnH6QOhfhWL583xljrukORd3zAcDrGchJYwaUrI6VPB4DEcnSy
La5crqPKPQwHK602NweiAYKLm1Tx0Y6yZjLoV8pulq2oWWZRaTjP6UIUpW/kM16ZFj5ULCd4Vtv7
BxlFz7AkZ7R6DvidjpbtqNda5g/YVl+j5F8mG6cvVFIkqYKRywDMa6AClNP4lnvXHh+M+lVfCryx
sWNQsSpIBHfIJV+6zFSIEobg98msJDqzHdFczqwyaMbiPlxiJonhielbaR3K+lWAIlN8rbfy/aGY
tfxvyXtdyRpTn+BoW0ckENOdRMtW2Ridc5EaFjR/25cQCS4q18MWAJgnIAs10XqMDIFORUQmKgaY
AtwcseYnKNeNUi68raxSp0yxBhQ9vBQteewCSZufXQmQp8vVHVCGo0H1wOuFdxbJkdJ0rrnX4ex0
KDZjaP63lnVl4DdT3vVoFINGjAFbYVlpauRvyPvugqRCYj3d3V1oHFwthzjzLAGu6ICt3Ao6vm1A
v8CfSfyijOGwvMlkWKTmnWaVNoFoPLzQaiyyAdfYs9yyKaJrxdBsekNOdZiXeespGba/R7KmWLmK
iL2wutqzwQ/noiFY71/A7uD+/0L0n0/L0ckaXEoknP/tNrD6TP7IvDuicbWVNaKzPte4jLIQ3ivQ
xmBpRJ8fUxjxgMRfeH8z/dEysrS47w4AcsN2d2fOg106DXbpL5dd9MN/swPmoenwFCvCQnCnO2+S
iuFF08TikEUpOO2RYGM2KsfcAJf9r/8rruDkLJpvWOaGre4ZFSMtdSu32/ofBgY5QLMLsHRcSLgR
syxFcvIOsi/qxIrx+KeOzEYceaVruu0dALuGOnolIIcOeqnzHXiQwZZt4A8jUyaLHSLkpkEtHl6+
EG/69PP6XzBlFeIh1n+EQEYRxL1CxYvdHEzoth93kRZZIvWIvxmiLYpXJai+oeCbo23ZVUHrkJ/f
AMHE0pf+LABy5wfyOvXMf6Mz7lUI2hzf9Zy0uSRoAc7HIyLfLnocgQGm2ezkpmucAjhmPWbDVspB
twiZRKb4UVWg+R1zPp4GOGrDerWtk7fuLBhBsEHuEl4G74/R6saXWEBnemMIPclGw9ZMDnkJrQ5w
bMFwgs2E02CIKplAV2bXmuR0Zhu7vyvx+I9Vity8fGWEmK2Lnv3C5295fe2zHfaUMUv0vZoIixoe
vPPOQBu2OdYM40oQ49Rv7WZ9IN3MXxqK8bvUTVU5X6v3ANCm0mSod/+mSsRk1P9QzcoG6O4A82/r
gjzJyFZXr75lMS7U4pWydD+HsvGUGr6/F4M5o4vpZWhAlkx4hW2NcZXjAIO2Pr6Groqfwe6wm/Jw
B1jGMJhnRptivos/XJwy1cPmsrXdOFwTn2B5lTijrffmZTCx4psd/fTQ/V7oQAyQ6XSQ5BLw9+k7
993kd84imS6BNepffHLSB1GdoSNRUXLsFLQe7ys9zZ/+gpJPsJjrOwOjsJVm/dGCANfQgZoT3g2b
RuYo6UZZYLLk+xWNIZsgx560rIR9eC+6I1GgBbemr9oW5mGozz9QksKa2QuiMRAUBjqkV6SQcy7C
72J6UIRZTwKtUbGzZRUMR0IOEZtL9vRugVRUw82JAWKo6RsrJ6SeEN4A4jWes7snIqj9Shg4+2ab
1Vpxx+bcd4+ciBfJ0s3I2D2JyO7pwSNPG79m/Xgkhwpgy0qIoM6ISFh8F2z1xO2s4EYpqbQawgUp
YZ5xilfD3cNY7ASE2Z5k5vLXFSNp3Y+NfkTVNIJ68rwmWIzbSLcrjYUzxDIl94iuqifwSBBcpo0o
vJ9vv/j5jkaLcvEs5eDKRfx8MCBsGzqGwuboKZEaf7M82Zk8v/d9Vpx9SpO/H6eFGhftbZNnGmCP
zlacxX8z5LQqH/HmA8tyguVGptWf2WkMy49SgJmvqotYW+PMID/Xidv5l3LpfkX3p4i4uW+Ybyxd
e1iBuqaMUSGjmjbGHq2ipBLTiD3kKk29EX78dehh+epVb36AWq/lLNFlDIVc6phXwZC1F6MMONQ0
7B3L4C0T1ShsVXEDjdbFaAzgabNl4NqB9n6Mo4Z6o44m8cIAyHuJMwoKi1JXKuWFpKAH8entoOFm
T5LGIMwJY5ZB4JzeBiQgm/bj82xKt+I51ooBvlzMy3XzD3SLSRXHx+yYJxrGzZbGXnvs1Px5LFKi
wF5MrEkdTS27TJSiFRiAMkfkzuZqLF77Nr+jgFr3ikfYlVG62p1F50fSdYp3QzU44+va/Y+a3gsC
aMQntnzVTGacdgPeVXqNijGpJSqrjO3MTdMtsw74k4fW/h+Ou0zptBMI08VklY4iUY+i4+7EDU/4
xdyHTHrJM7OhEQwt4hsoqMAZTH3SkUpEv+HgRG2MjjJbtXl9IGprfwf1hpll1xebwxsVvBkXvpwN
UdXG+VOFBrF/gPn+O8G5Gic4OA8BWl9Hp5M8HGlzcAaT9MaNRig7CxjfabaH7CBZJFy8vdCXEMiz
itk8oNVjgqN40CvHpZUw+stKSYgrnjOn+s6vccXU3HrfaSqcvMmse19JzxsjBGAjI1+CojG2y0RK
4MwTBDiu5nxdTWzpkGYDaQfB6EHZ/V8dsb4rRDEpKZ9owXRobbY5AuBUJ2unPNUGQlmpdGXjuixk
k9TzP2a0py6Sz1Fxp0p+NpAdwro8Aa7TqzoesI/E1/GxYVeSZUmn1HLO1coybanpQnnbjk5tj5SL
KiO5bYXjl0l/icOzQTwiSf7qjPtVeN/0m/hp6xQ8KtvpdvliJEThp47WIVM2BJ9Ondtx0hZW93+8
hL/JBk1bJ9rt+bAzfkh1uTm1TQrB6jre607NRe4AM5ZPppqSWODxM6IJvqChG5v+NtT1QPI9gpYT
/AERHv/3r3DpycGJhnYAJtzy4F96Dblb1YUe/PBvCiGjxNzRiq7ETShnq3nvUlZK08zx4DJvJlKU
PXP6Q7Nzs63GhOZY1NVAzZhKELDe5HBzra9rXc6TUyUUTP84K8ikubDiYQcdmpmYb4hHsgpC7XkT
fUHptZ+sf/SZsGYzHL9WLDw568i1CDo9l9P5dpfGm1sNn7jON8z8pkGlnP66RbZg9bTPp0z3bhgb
xM/IEDzPWOtLnCLKF3d5xh5JNpFfe9IS2GLifcwHkcSm5pxDxVygdn/3MbXALdn/jpY/geig/H6e
s6Cj9qrfGjvmEUw0tm+rui49KrD4j3YkKWd4dht8iqoR88tFSbllFVC3Qi3mdQ91Lur9Sb8lChLH
8quz7ozqkR4Z4et7uYlrCIuhrWksUxTOzl/eTSiLMVW4QtQNcx1IvlU4A2x0j9Wi7R6xcGULCa+d
aaTS4IILkFYjjW3wm9hxU17l7KT+ff1NUyiByTIb2XVi6l2frOo5dp6FcH6u5N0q+pAezMN04urR
6s/iL9Hcji1V960XGvvSbQj3i9jlE5Zc47NAv9f9gJkKpgnhK+547EGDcM9vtfqJLsAlyaSc5HK0
lxYp/Z/lC27rrhqCCmrKvFoNoDh8qyTHPDKYQi1BhVAkvO5UJSTocRIChaZJd2huDNtBu38tjude
3GCWSd+7Aix1/Uk6jhpR4UuaObnLnDREyRLnoJBldbVWsvXfRSC4zisznIWP1tQChu27qCG2Y2o2
QjUbVrPQw6jcwweUyIXBsHpAF5rcVWWAAVG1oRPI1orwx4nDyKEXlEzuBfbqDc2E+PpRA9/MOIAY
pQxxpJrcEv7Gcl0PEDIooiJ0WnPJT97cNbNkufvVjh/2R+mcFjf8ek50biSYw23HTsfKCFZuo2Ww
q7UIy86VoO+UD/0q5JKVtzyVurAoipOSGtiFRpL6WAA1wO4bK6j0h0HgF/dfzXGu+1dlpdeA4ZTT
0NoWnspxcoiKMztHx91bQ6Km9pV9qMAhMI0SynI9xvd6hlBOA5L3aFNkRv/NnOcEWsubmqFmQHGG
tE/Ej6ykeTxmpb5tvfBlH+cH259U2G1oqivp4v3HRX+54+MM4LMOVpCF18pCj6jE7XbqrTdrqb4d
0qhTAmzzWvssx1o08uhphtDZjNgM3QXoxZVWuVh2wgmQkYJsl0I3OsXN7dJ43UnW4u5T4geQNRaj
0lUxgpzMNsIZ8frs02yydqpFuRj52myyDLA6PWubIHc4QiDnI+sFnHHMrQWImgBvSGjsnQOGpyUi
1aYSQwLoagIVZf8TCdZJwFnZEHz+T1BkK2dJMv0nc4ZVv0Ze0fXclRqlppJxDCKMT24BCek12e6P
9G6Wro7fR+YKe+I4bXwXSNlMSyi2yC+SQBeGirdg+8onTe3qhYsQjJLW265DJcsxpBxZ7UUhBITN
H57Nf6TXUTz/y0nb2jCnppC9YJ4Kes77/NlKdK1AB/9waBHEVcJOTlt7kjqgEx1ZeqA2D1N1X6lY
j7AxHWKDuFcDnG6JnNoukJiBbrI062K9yq2VlzJ0TRCgV3+aO+kW9EEkGgjfvxbSEHji+4B91xxi
7IeFN1yYvBEbCdd7Ygn1mV25cf30WHdTqddE0Zqn3I/JcWq+8otmiDw7EsegkO4Bms9CyVhkk86e
KEGmkkhqt2xOuGahZgD4WyW/kQkkYKiIYX4MANkHFv5Qj1xzJJuw4oVMaS6uNGqnURCH+RVfgfn4
GKTemZv5XmNMSVAvaNkzF79sLxvjho/NZ0XK0mt63BtBWXRkrg80Kn0Sw02nM43W+tTCzyWj7auc
RsxZfphZcRBifvKzH4ExWMm2C9uHkfEuczWXDscMVuxeTDiB9NfhE/WVL3zcmzpWTurJhBctzsqZ
JuoYn1XtkBsm+9z9LadS4wqfuwGaYuK2PEeS8dZxqgozH/D9bhUQgQQjRSZbN407Gr+4wxnsjZPm
4QBl6cyrfE9lnFRnUrV1ltz6iP/OleR/QcAYYc5LlTBnr2qhZuwNLEYCoEaL9T17daOXkmP03qer
LEKsd8B5mTxbh8SfLp2rrAMlEDzSC3MW7pbB5V9QedgLUBqNrwPW18RY+sZ9cYLvL9CbkHfCD9jo
n0kYdSC3BEpIgKnAbosLcRTcAvjLLwY2ckfWO6q9SENYBh2YaFD8eVCYIVU2PM2ZoN8A9ZD/J4sn
nJaYACsczaFUwLKph9zVbvk9rKy1W5R0RtJUDKww/isxbED2Z625oX8PbbyRGoaB8XrRYMURto6/
IFVpAEqDl7BDEd+ykiqLuNEHviTjD3HFOhyR1ZO+EQFWcz9pCOBa7HzOEN0h/VNgVxbqBXnCW0o9
ODrrk4UsxZD9wXqQ1yXTEHVtIR3skT7CGwyOtl3Hjl5xqwLQAoKV86jTXceJQZr7rfJDjmMwPP9W
yHybdgC5wx8r+i/w9tS/iDGl5khcixRAOfb1+vhEaFUY2IPJ6bvFqAIZ7W1/9XtruKUKm7zwR/30
r4NEfyaHrCdLkkjyoeH1Ss71EgMvhhysmjrQkuVZm22b4ndMg8TANOCgaGykDPaNqc/7iemoWYcj
Z3zh/NNhM4VyIHyCwjPLLYYDvZfmGb/o6CA0OJG0YyNPJn7lK7JW5FOtsBaXnmWUT0MXhzbBWNSM
nG2lalznwkoZIUgvdWPpd+ibK6C2opjR76ZvkLN3z34TIuZl8kh04UWit+pjypCqYYPm6fAQZRc6
ldZ58FSQAimWFHIaCqe02iyMavAk9HSdMls9Sy17DWD98+BpU/Gqwvrl/3flh3jMKwZ7i5kB6FoM
/9virCHkvYYL+AU9wASUalA9U5fWNzHkrZR6bxwvLIqO9mWMmP2hMQyvsQwIsLBq2KZokrgYLgnj
lavqHKWK73O1FkUCW/S8wb+RvROII2sTTs9qd3hJOBJlj4vU/1oHbavF4rarHV3dxYt6smY3LA5v
TZkl6VkPMvkTi6EwdlZnlzLB+xfTHuNrNd0B6HNKQ4ASq0CxYkvpk+8pflw/4z2cJTPa1HKCFYPE
+yGkqeuzwPwfEpBLZyApxbfeQ3u8Tx12SHkvFN+Qmo4vO2Aqcrqeu9u25KOU/iblnhCVufn9+uo/
G8plsPxS/GLdGncofEEmbyaYUFqfDC11OprMtsc3F+ApMKGAV1aE/v0J9FHYBv6jaxGhuq4d5y3E
m+2SZFb+LTAErCJB31BoULVy9RpagvXEVqK0H7LvlOBaPEG9s5YD4adyzc7ivYo9u3aqg7m3U5xb
vZGW0aIuruwWaVwi5vh5pe34bxI5DFTglwdCliuiumtboO4A325mRoU0tuY7NFYjAhC7b6Xjf7W/
RyGE1IAWpNwp/reKOijcdt78QBARl2z7XR6c/I5IJCjRwuh2VMP1VgHNNDJvJtfR+KRMZeHjyxIi
0BVygcO+gKBOzsF4dmchS4MFGvUup1qwa2hnEgMXsMATNYwVwve8n5Wxff7noh0zVpe1N+RkV4Ol
2WryCmsXJ9Qx9EdAS3z7lZTrq1gxM3PNt19jK6YfT/ChW69qco3yfRvY70Wd/WgnhhW1R61Q7yK5
XM0D7y+gy17TbZ3goSp8qBC0GGE8VSDqn9PuBgtOJI1mAETtToXOPIvML+cI6X+biM1wmED63fMI
gAqK2cFMcBT98Ffy57/BAq4Nix6fIt8PqaxLNE6U3q7AwLHa0A4ZC/prULCVz8HU8KeA79D9+e/I
1c8qMsrRxVWcsk+lrLgCXEcODoUU94Eu1bSd2UTDfv3Avw7i2jzOuBTGwqm/VDv4/vb3U8UrA3lV
e4v6ze2NyAG7Chl+DR6WIYl0L9kVTiY8uL6cExPsKRc1L7h6eRfmUKkdqSMFqXM84/3V/P72peBP
GvRzvuHwwo5dxPCRM6OCK33WjLQomQdTC1l68fN03xFFMRSvlV+Kmo1WLc4utSYxM+Tu4EPulW0z
jO1dxloNpkRDuLi9wCEiKQwpqSdkpNj8wa8YmJ1jmtZOz4jf2HvgWb6afItdHp3ewlkpqUfix/dI
6PtRyhGIZ1kpKWpW7vz++P/h/xncz9iXsPL8X7+p1OKQZliOzWXkgP79mZ7k+M80RvcA8Rj2v+Sy
G4zbFWPFk5WcVVgrxAzXDmoRp2tUaFe4AFi+88i83GFTvTZ0ZUYm0sjGI+bhnLP3V0rtdzuyNpob
TBiHfqFpf1Iy3c2oMG+HPcJrBT7pCBHJ3Zn6ZRQWKNn1WM2z5n+La8/HN/yHqboy5jNlplCxCLzN
nkvdO5R/Ma48vJ+94rrhnV1luEcnN68oiAT6/bHlcD1ELEDNMQbYb78vj3xL+HsH3fJLKpzTb++M
8GyLsjDMlzwb6mnz2slCIlNJLxsGVJqnx1tvSWINdCEtZLbWyrmElEauI+zJMbZbyb2TC7GlGRiB
l3DS6toBQe+BPkEGh/E40p5RDgqRUsRjNE4XdgPsOUKluG4jiF0KurZM/+kmcxJPwGi6K7OMqSKE
5GjwE15UL1tU1VYacj8o1VME/ZAoIL3o73qytZSiYDCasdCA1uTM+OsoP8MDIlP76wW6bcbEc31t
MKO5w01wxoZeX5SsbG1bNsSdtQiKbtSdQmvkuGsOXOoB3zWDp+X9kNIWftN1VI0O9EQ7OGp2p8K0
JeregthCETD0ZCumxE+PjmseIkI/LuLLjrkzg+uFWNGanJfL/ANaH+mfg2tC1v/jPboWBkxcwflv
G6rrDN3QViS/wTFlMHhh3ls7zaWa2k9ysmcXGbu4GmjKa9Ap7e7b0De83qmM36ixRchdxXT2qWuk
xztA7dBNWgz687Mw3sONXBBSk0XTdQTLXUxNRidDzZkPAfQmneAC2Q2iNEQQP50DGirqtAozQ2gl
YN9Ogq5o3BObTOHXNEPeHlssaceyqQQ13suGJVSSkVEOm8F9/DihSGWdI3ID6uF51Bg59LNRZ8hK
OqSqrPuT4XhEvoJC087i39oWSWLTtNDKyyNVO4Z65JjJ1eMXKSE7NLARrGANiZu4DG3LzQOHS3jl
r1ZVtjRF03LEdxltF+F4P1sOt2/zlACCN/VtUzqbwLk8DnInTPCjFvPaoK07Znq4Nt5xhBVzAMkF
wm/gqnKqIFrrPJ0fmBYzNEgUd76Rd/HfHr25gGigKEcnDDTM0qJJQySxbJSdTrHDP8qnaMOr0k2v
krf8zinnhak/K0YjVWGYv7PB8Eptsf5R2qvzTMafVVMfUGu91nsQwjjsrw7drfqDZOlz05wKqcKW
4+ntE5fxsrE6UYZqUpvbX/ih+KhbS8+bzIDV+nRkSrkHh5jwqtbo9Pihs1AHOVZcaqDq96IvWThF
ycFKuBPMtpl6hC/DeZVJht+aLGarZNF4Lbd7fKA0nrUWvZ63omMm6qtqYKklnfFrRVGrM9yIlZPl
H6g46/7Fq86nXro7tYY9BNkr3tZ/ox4q912VnWmZRiPuvY9HGxQK1sMlQ8CL5nl4+rThX37c1mAm
PZbwC6q9WcemcO7vTLxkCqKEtNHKVLvrg6HFQUndwQrv42D4/QmpBLskYUsGhqtgC1OJ13AT4fic
8XcmJxRPiwg7cSTH60yueY4ELo3qwZcgOnr9fLBNG9iJ/zbUKea9bXUrP2ZGNXK9Kvo8Bz4Isy+b
/rw6jrhspFZf2l7KyBXxrxVEqOONNmc9oZehm5UcAduHOcC4z99eAiBmDtMXsft0GzyvZG0b8kwL
C3Zmkjq0vLoWfdcsIP7mdCm3Njd8lQY1EYCPz4u/fO/xmxoAQD/V4dkEp7FlBrFtXfCd4n1qbKPe
NnbvBTn2jOF+/8fk2imDnaODuKjHE8xXdjxQ1JE9rrBYi9pvBMkLWlym/WUgmBncxE/NnzWzRpbj
Dd2D6ZyGLuEMi/k/rAsu8H/1G5fWrGxEuYxx+l54OMqRcoJcbYDc6M5KBNv+ALll3Lb/7Tl29Nrb
s2qBVRBk194p26GS5o9iiXrtKE6cHJovDTQX6v7eP7NSpcaf4HnffzlVQuQ1ve+6/GipQC9Hni2/
XJUrPYd37CAZFkZjZ90dSRHVj8wi4DqdilwbUvvIMS2HkSR3kcfuPNerP4TggGriYIMi1cQFztU3
9TUdX5z6Z+th1sQSuhdk/rX3YJCUmtURGIIPVrKfmjOKiDMN0/2gPgabMThglM6nvQLXYHCFGuTn
pdiLugAVuJFpCf1Q44IU9/agmihhGCk5ZwExKV3kAGS/G627o1YviDgtbL03hIE8O+T1B1JqyHOn
DEj122TmqrcrJgTW0+sjyKk/2xGulFZhx6C/njGNHLaSL3QHbRrKjx0vVUqiJfH60zi2B73DT7f8
/HIo0VblytjAiVElINsWsZzr3xjU64tTWZ8ceU5DH0je0mKfDjDq6WPJrqxTGDa9f9r5KneVga3j
F+XWXjhfSWqnYw3mb9SyZHnZCI4wvpWKgG1mOeKxt0pvrOz1oXrlGrdHSYi1wOGVS2Gp59QsDZOP
m76crYnrEbibLpzXeGhJ7RD0X/+gyOfcVNOjfws7dVg1sdjzvypDG3g4YWG6y0TBKUYKMhgaszzl
SLQTNO6N4lAp/RiAVUvn5CZl+z/Rn4E7fZAuSHvDIv51UgG3/htUpSXsBYQiwfFxb3JQZK2VTS7A
RRoK42nv8T+XteJ7ka4BkDAvcg39mFXaR2j8hHtTetnSYdzQ3MoeI89mj2SVJnTr79UT9o8rg92Q
KEQo/EBIpVSvRDQ+BoE60FV60X66dTc7xhgFmuoGBsJnvMoAweM41skiZnARFdybbIgVj4Bh4gq4
O7s41vJius2/XhVhGDLy7NygLMDJLm0I8TAeeA6oPi+CXX4Jjd5v1Cx8R6kjwBHHZhUg3qRY6A4T
QiUoa+uOstimtOI7ZJqCEo+uatbNqoP9UchuVCysRMqbsGYWCWUHsAr3IW36gQRpEbJgYrxL807E
ESsLGvOB1ZDYWvwklKeeWVex0/2ezYOwFpVPPUsTBSedpbd0yn5C18N6EybqrMO7aonFsq0A8JDS
CDQaNTc9fasVMdw7h8B+tMpt4IMmzVIAHdfEQTO1Vmvwr9aOmwAtrkfyhSWjt8+COIz0EsNS2TUI
AaYuKbVJTVqSlepODgH8yoXfeFl67/BexNcJ9V9dTAC92+Vjp+2dxHUPJKNMkheY7y4XLsHGf7af
BLaJBRPkY4RBUMi9sVvynX+A5cZCy/o1SDQuiSipGQRMTSo0a2/FPw/42+cELwy0Kk68InE8d8T+
CLFjwK63aslDmqwOpU8BHkvuZtBXyeiIAL/QcwJ6uZSFksMRkNOzCSUVGe5FEMo/3pc0aaqiFKYl
D+GNHL7A48+LErGN4Z43/uKg5D5o4PuMPmZPPt0yKr/+HI+dAqJVZOzcetD0jNYuXOVEfB8OkiWl
TLCESiLtYdKKrmBV1sUtIorPz4mZyQcmxJXTTnYjaWZPtqLV5XhZxoAgQ1a5pIDtxtMaaMts7iii
ZWnsmiJay5KZT2JRbSUSzPeZsMEYRD9yy3kX0dL19dJjz6I5AhyHo5HZhSp9Z6WPhHCcc7ifEaa+
igiajLHFSeqIBa86IAMIwcb5b/gXsq7ldFMXCNplub668zq2/OJsZ/t6tWqwmeecwOaEQmvF8hwR
CyTlMKVJSBqIKyxSk+6vA6o0LHEzijawmZQI5YYUr3rt2wVjbPUPpXYQh9zEVnA+yfAD8/mOFIWO
Kh9FA4/qGfWKbk5DCV7+iTIIw35iEZo5y2y5bDJwL87TIKQ2bIepFmyXTXcPDxK6FNGiAeK7gVW1
lWQv5OHNQfbofDSHgHMorKrO3fsX7OAwye4/+6ZsXmho0IMZfo8w+Y9E5HQ8F45VOhxCs1/Fe5zQ
qmuODHzAanE/Ft+m1U7wE6p2qntMgOZ8ne4b1a0ifjkSSgdqAifhtMyWBWG8ay6o6XD9S3SGo1BH
u6TojsHc+B3fuc/AWzobR6gAH26wiQjkYecy4dUJs36mzCG1jSN0AsL9yu0xa5ccj9Il9qR88rXU
lgW3LF8S5SPgNAfJEzhZwEN2JGvL8jubV07eMdHEm0TQZTg1mPsGDqL+6dFxf/ugQtahaRN22Xir
Z0lnUSpklBN2mzvw8Y2z4gwPNHYRg269Dl1SvogiOQTLDhYbhl/a3/fzeku/MLkZ5NI3Hods6huN
BnwHgQQXwaAqJb10k7uNh0yEi6LYh7JECcnwuJeWllyvrzG7KSt2SHoE/waayrq22PWscNi/B1Qf
8L54ZvxDHaQ6zPySUHLc9IN8JpGXjXjWLoNaeES0b9pbwZaX845FxW3NZI7bBXdtG5NqdAahel8P
pnkvT3TOHP3xAARa3SjLEyNGgkwVOAgU7x+tdCWQmjzlajoHM1VTYiQQmcaqgg54yB31r3Z2ExNO
uiYyEKjrnEDbb4sgkO6bj56YG8hgbGEreNv/agxr2HzYTDZSIXk0H1MspVSfZzwgpKKT4VT5XOHB
liDDg64g5hkeWzOu3emIzvzgFn2omxEcPsrQQYzLQp2e0v8H3KA1SXiNT+/YNCLCQOXlAaULjRV3
ocRihBv8o+5QMUKGIFWvSAd0UaS5cTvpQFxDHVroKZMj5/tZf7tbaLb5nsfADhbThTMTu9ohGuaO
dIklBCJ7uSylXXlQTRhmUeTQZFjiq4jH1XV4ccbUJb/AR8PIIMh+V9OOq2eiPA8b8wfykLfl3obU
jyWOHX6cN20EuO2lWWU/+yx9DQyiBe6O2DVJkghOMM9I7/8AvNkX4ExKv8xdiebkcYF5Pceel+dP
+UVRG2/q+n5s0jkMHqt45g+YkWtru+f46xwHgBLEn8Tze4jqRcnSiy9hxPtuDgWtjGm38glpCXGP
tQddkV/KI8C5IGhUo5CWO62NrEkCh465lVtXjMFrNPdPtp12Cinwd6j0zmawTIvkF4Qpu3htMPYJ
dGI25HjbWzhgPKj+5ICjvstAEWGFLV+C/RQzVfnAROTo07+tVVfDS7d728QOtNu+mmksh1YoJqk7
gcqoChq5IHS3dajd24n4tctt4j2Wx2rb2qVK4YqJMA2gy0+2UQtBW5/waYRFlUpOBa5RpxRXo33n
rfhEnz0s2Xf7vJ2kJq07wiSHh/3dGoqvYJJLZ5v8IXsXjfUX10d5nKfS6JeEFwpti33QBfZv5kDs
QrgZjvrGzfGuZvaT4FckWgB+pWs7i1GJIA0mfZqoC80K0jqVsoDnQIE5FB+a32agN7+3D8KQ65vt
q2xrGXti+sb8LUAtyNCYeQ2k1jrB/7oD7Cs9sRUaIUBXVXp1CTotu6np3fHKQc0frF6r3ktvxpMU
hYbZ/R30x6CLLbon4Dr4Ae3OaG2iH1sHXTyXzOm+eDO1OjSwG6t25vagN8LyMIoKjCqz/VkErYZR
OcydepcZ0HRFKPRIc7c4qyVG1GRY7KIUUHcHjuJEmitEHnKdr/M8996DoRC/XJ429MihjLbrqh9n
KX6BdbL7c/2Z5e3/7m9ks79TUEIwiI7Kh83ieS5QuBhfCXo0rEkXRjb+hKRjFKPJ0GisK6MDstzv
UIqP5oqO39/AbF/fUnUPp4BJh/lEfEiyMHuI2m92/KdM19VXzUjAEGCJ41XWN9O4Qk2MgejTCClw
b2ajCpMpJNyQvQymOOG/4ZNI4GHbRmiwokpaEXHwiji85Sf68D6/n4YEua4X9U7CYNEVhe1TAs3S
TqccpZ8Q+zIW4uzsRA/8BiLedzyTTvH6wDTRyYnPjgPdcuT1DbHnfQ0O6i1GNDZeQxa+TNQp6ads
90B8pIjfBX2tH/sbEv5XykS1iiJ6+b9LYlIBHa+PrCvj2GUhfYEivoKRBlQ3gK3wZsNbuib3IFGZ
h6BuyH2Jh87f2PbLMS0/CPD1o2ylI9n6/2ii9wZISQrEmI9gZI5Axn0PwZAyh640St1VS5YWZHN1
QMD1RJVnDfJuKG7+YYmJ3XNq9pg19FZ7G85Znc5oNNYJilxCVPN2KdnJfo0v10V559U3sy4qfh3/
dMGNCQ5qYQEm45ybwPKIDyiHkJCd959FE6bnZLLmE0k3fyM5VuJV/TQK4Uao46c13C0mX98TcZph
+95GAT8RTaqtFEJmjWucGKurvkUJXP6eblenh/Hi2pWpA55F74EowA9RJE5bxpQHfbQGLmK5feFi
lvz1QmtTYpZzNLY7RHFXP87+Z4ibjuXw6xjxSyOIm6XSYXWww9ILieReGZ1jDVaYN37XKGsfKa5W
s02uyLY6eRHMhDD2D+DtEWEAz/1vxciRx+196wmUsubqdUq3Odmyn3H/uhrdVW/E2zfyA/bkcBUG
wFWWNuRNaKvka1ygcyqJ3Zs0jRrICM7RxTUQna8l+DfabuRHAWSz1cbTrncD5Q4UJaL5lIIuVelU
OSY2FdY5ZQdwzA9+xb2fcQOK2FmSEdXWNJCfQ12/4cTgPDglQzursiveGe5LpAMUKDx+edMN7min
ysN4vjh2pbg5svLSpJeqdgLDcFpFIZJlqjcPHlsWZyjq7wkGcOpr83PCo7UbKEfx6ey5Wrse1fYY
dsWRELRC32tbVQ5+Kpr3ADxNEyXJH5rbOXVtikIaDpkWMeW9bxuAI6Nn49JKlsLiwo6kmBJhYWzk
mxttKd5uI7qq7sKr1/2hC3PkSeTmqrcBKk1bvCvj3AdYVzMipYFHUBJb+Aqv3EN5gkTkglOQEpM8
RNasmL/PDLXx2Hw57rPvDjcLnkVMRbI1lMT22GwjBbP3hxf5t4OmL9YC7sFfATIiGvH025g1zp+4
Uci7W0xnCrBx4iB1KXFl+jMiPICk3CDqj+71l0i7BGdjBR1xHX1qvOIfLrnRk/xhKuutfk21tpfF
7/AKjTN7qTntIHCsJrwsZdHxFJRymbQgLoOKODTFKssIroYJpxuRa3of7AVFAIU5qtKpq2KFtJ/v
8/dzEs2kxOZF2tQBBZTfR2FulT/PdzaWfQoK8ORlwSRBjXbsISHa81DIIHhcovffVIySeyN17uF/
hA+dNY2fi0+GCcGPwQfR72jGNvOVKFuRiC+Xyx/wZnfHohh8tvkKpDA0bigbW4X1t9svFE4NxRzR
yUFaIw2cAAXLVvyQtj3oghOMaYTNVyZZSP+YtN6eUCZLvvRU1R0xWduFO6Cx8zIvKEvLsCuylacx
eNu0afd0h5F9W6o4kNwacyU73/CwEyd6duZMUsOinMpNXXwbqMaEv2PfTjJhmvfgo+axmgqj20Tb
kl6dHtYSz4rinVCy0dbNlryVvkQCjeTzRVDEZNIGeV12agDGbG9nzTUhC71KxBscvcIZZfJXJ0MN
Lp80klITbRAZ2ahBhshZsFrL5oUR/Fo6Bs+sCON3RjUtfI9gto8ulHoGgVlPR2EmvH6i86z2iaYe
Omvk8nTV0vDVU4faigR1zDaSURqWOxtnWNdOhDSWFHlTwSNO51e+lpQQfGILs7TtHfyB48+ZALJa
LL4kUAfMoRcKsm8iZffpboATPBwKO4MjrZzidlz9vw+AWQHgcet60S+gUu2IGSJksaeNkovcGrUA
rHT01T4RebGbKr7czl/XHMIQPmizHBeCGnVpqOE6tiPBfH+R/hmhaZvaX7sVFvEOTouJniFkub5m
xWTYf+N5XhCM2KxS0GgbGa9Cp+ab0FYDEx8H+5npRjzx/WEfCB/yZZ3q2JVMAbhC3NU8MlGiYGaN
2yxO9TjE0zXQbqiuplh4H35Pohmvy+W87UsR97dGTebalvj2/v36rPaVNTNTdIC7m4sEtYIL8jVZ
YRsgaif5DftBuWWRO3GQNJkN+4gPT+eJ3ZodTsonlSA8MifMjswL6MHMoVCycdduS7T2sRsC0wa0
B46F9UjDn6W83TxnnpCgCeWZH1w8jg78aC8/VBgWKedv4nOA4ufDmoOCuKrk1mgGCskYHURm1KhG
b/MeBDKNvlY+17xxpX/0CAK9CLoTL2WJ3omVvm3ovnqG/No0mH0Q4nyDV5XlTg9d8tFmRKXqIhYi
aUJdyBxB4UNEJgyivXau2eW90dJ6mLFY7RmJoQES6eKe0nukox/EtZ9AM/RSnU3mtZ/pacjuUmo4
fHguU9bdFXbP52UkB/b3K/wP36HXwd/hB02KRPJ6sxocy3dBjMAByPELbT6dqt+P+YX8YTB4XOON
GbM/VQeik5++uo7lZcyc+jDO8j7rO3Gu2LieGBJbebJLl820t0nLo5Egh4QOjN0dggvjF35BOwx1
RvEZanJCZd7T7uClCthbGsZUOqtW8Wh251J6MjK4TB4XTf8v0WOLKF9bO6V8XavBnkTbQG6Bp9/w
ayl4t4cndMwIjyb7iGu/OFuLu1osEWPM8Zk8o+9hPdA6JUTeKFAbsvYPZ50NIllSlDwi9qd8Wu4s
LSA4PEIo3O9P/DUvkG0MyTQ/oO+6YSodtbNsINNFcVA65U7o7/RoC+cQKD69SpQdOvJ+Zpnvpp/d
XbL06GcDo/NF8PYXdPRzsfx/74wafUwTNYA9m1yRZrsFx+kkbvY9DkunZw4DRYRGrtlmdBz2Ibq3
CfkAULUiNSzLzYrRZd/mzlCBFYiqYrzSLWPSDTyodkcZxjE++VhMjXY3Mw+KjdJNhK3NTEVyzl81
um9Q9qdT68HUFVXBuCHLpAmo9+Jjt/2U/T/fXaUa9qF0Lub0vfNoKmi9LoBcuwfpP1fBYzKzG3S6
7cdqMenQurnlUnS49q65zMbiyS7UklnbB8oFj7eFeYKG23u879clT1ytsxHse7AsMB2U5IplnWS0
B3Xl2gSHz8Ebqb6EUfoIkKpKTfKJVAXaDVdj4gGaHVsptuE9yRP1cZndPPlkaZHD77hT0k986+8s
KT1dGE80NxBOy2/etL/Zb6gZDaFr7Xjbfc8Eeu0juw+UE60rgQHSHQkNAVfU3Xg0f2fHVFH37YOt
rFR5z3mIn5R73jBobN5ZOfrDLbj3vO2InFke9Xbhvu5vy7hzbX48t5ExTP+UQoqDkGnspeleOx5N
UkTvXw27uagQHBi7z5v1tADcmh+59lsjldexc02S9uyUE91UFnXKFrKlQ5gc7IkGm+2dwrAQXSrP
QJW6ptiY5PsUOafyxftG5vvRjc786vCDqnjQjqI92sftrSwjPzZYrP/g8cHW+OoRmrf1RUTANdED
NJjIFwthrjiJ6Dco8/NN3UeLGuo5zp+QQUd4S1GAw0A+BzyndIo+WdNKspXxdWOAa+P53RJ7H/eF
yXKNMAP5aONE+EU+BFt3MeVB+rzmAckW9/JhyvuWsLke3QNOidzxfrcu/oA3bU0k8YmgTb4ZGR1P
ZChS0/FGw3uVZwbZSlALsl0QoQI/U4pz2ldvhfHcHNJkNXW0GVzFczavqn0jHSNIGY+/ISX2psBQ
+ksT07O1NdOpXZJow/ENcZYKYqdxLkp4sSSca7trKoZBboMQiKruO2c0+yYKMdfD8azQ7+h7HV4W
YM6UriTjwwQIMr98ARntAYGERkEqPCaJfK2EOVQVr2misRXE2v1KW7gx46toj+CL8Xwavs3qapev
LXXbn3QrT01XX05TeRpnEyBS3/VK+tdi7989mSEitiATJurLGpy+gIa03FHDGW+7PncWhIxBOBLf
p0fnd8LY209OAJlY8lueoU2xEIRWMf8GVUOclZgNIH70vJdJ5lhEU+0vfGE34mPPXVtN0y8JBFUX
2ysWnaoNGOEr/x0/BPsYwyX3pq2m8EgCu1EiIv+mVbCrO1zjPnpruPiM2aBAxacnLTZJ1XYPTQiQ
X8LHBl/bfgV1oyKdZ7v2XthnvXSeIX4H7gfYPsYr2H4jTOK6w0izUBMJRjrY2JQtQcPjaCU9zZ85
EbZOVM3qWsQz+OF4vIe2uQk2VgfxHDb2j9jsb9Xm2ODhr77F9HKR6jEWvMN66pgLCJVJXVxB2lOp
8306Q/yshdR/KDwdnEsWbV2urUfuVhL4uLoxzoprx+aB5iA2kvps5LWGy3o9NgmObVoXzTGi3ZSa
HPdaMwGBdp7WcYTQqm9R+ICH4QK8TEgUO/ZeHYTW2hjJXUUtfh3J6q8BOdRDaYLino+GRYfBealN
cSM+feku6i8g5ao3VvJFZ9FPGSFbc/wX8bYVnhEkYJdG1P1KBgVCrvPd9ZZHmQkARCcKySAeVome
WYr3Wrza3PY9YGYZtKOxZ3zYJDCfCbB1epMXtcRL91xQyc12VCWOWBoqb2fJDVfGIJhsfSVHCTiL
5h0TYPZbMbO2GApm2H2MSVkdqbjPyb6v1OWt7N9VuZfVz87cvdSSckUdQhAtkjRLzRKDj4LVEthD
i47SJOSp2e3t1l/f4OtXkwp9/Gv/3Fz+wxdbDjZ+sUVcIIC/ZfqTwcqIzFRY/O+943aR+p5lGfLe
kFXyvCzytxoIQn2FRKCN5Qmv+9Q4CULuWYizKfOLqyEzQE1SGZLPymlrIpBfpoQNGfVzlVJfYgQi
xnTOyuUxVOjrGLLtvuBdpxPrSEPFUAmpREtjWfWf4y9UN9kzfGmlbkRoa/hvLiNi9m6fvRlaWXdX
gGKOX2Z4rTaDNIuK9v3YZzQsXkkD5wmZw8GLE+XMMmy9GiIB1zQ2dDkT0J6G0jg9DVUzOiLoxhVx
S/5xsCElzqFG8qEcxlQa3UqW3VGI/pOcpx9lLWGCfFsExvmfb5GtNkG+x5hdCC6C4XgFl5Q4oMBm
Y8EM2Sli5P76MgU8QMNtjO7hPpWLIyXjbzeqOvRRxahoCLq0woPpf3AT+U7YNKoi1Wu8SjrCUtKl
tHGMYw6r8oh4KPfyL/WPgEF+C7nFzWW6Epqv0LubLqiVhnIZl9fkWiiRQCi2y6I1R597efBH4kTK
vjIsBM7aV3eiTc/XVydnlJNU/fHArWhBKiYehi8fN3C7GXRIPa4ZSaR1Mx3dHuyhles1TB5QTn15
PYhY3bNgpUcv0CqCa66HqZ+6lxb+IlWtZBZGFy3wQLBBnyB1aiAaH1FrML9XVZu5KYwGTvmsWgCK
XTIC+gsvjpt2KEAaUk9nqokctxz3inckF3oYBK8RoC4HW16ZMonSETJp9gCDafCCkaoBvpAIiiOj
dJXsTOzmQrAwwb9a3GtKna9iJED+w1C23zAKWTE55zenxqE/csDczPHHewD+yjZuLAHG1X+i90Qk
1vFCOY5q+43iwAJveGHoCGCCvJPEUMRkQzw+y58YtSCZ6i0bw+Ss2zLERYzYtZybo9NluNUwYkjA
H8gN1b1ZRBn8LNugaBGLcqCojS0yYq8/c8Z2p8TSGhUpMYWuWIezWKt9UfUtXeDEKyQQWx4/XATc
9uw7RxvjJz5/ONxl84v+XU5M4ieGkmqQEM8fKHzHkto80YGzfuoaIvgjvffKmcsY9L0NDxvGU0+z
+pdJZVXPGSHB0VA83DrHYEWSICxa0oeXMcXwsXIWBE840MjvBjTT1IdN9cGX8MO++dWn/sCsy8Do
qMsnh+p9LfwFWFmeml+/kLkCWG65alz8uYQMSYkoTOuuJEOPM5j7mmqF5JZQT/lb4G6LojEk2DAB
VNTTdiqSgIS4ZyXs8Ix5ONDqRmqd0csep6a9BQHe1uI/PtgQ4+tRwxOw6ZvWHxjVjC+T0MKc3CvF
1K3aIOlBpri3dg5wKPJAvrPxHIQvEFvLkHo2d+JBNW9YN2V6jH/uIY8X13AaP8XtQt1JJqhQB8le
PBLPggFrb2iSueUH0demgGhMg6vgvOzKN8XhN3D9A0PBeIyWtGV/5lHu/82oaQVthkr3tk4V+uhH
kP2JPi6EZTapihxHpPHPzP56YgM2Dq6Qsi7Ajz+awjEcp7DyzhoGOwKxuTaU2UgU8+fiEd/DkSQJ
HzT8YhCSvmjJ5obAnEr37/5zdqgkdguEdCpxHfT+qZUNouGKat+2BKWTClhOxpDPJCdoGlEHPltK
gZ8KwAlX8zIN8eT3FLhGheRYEyaRj7G/T/IczVyLGa8LljSa1N2Guc1Rjwc5VJiRMqUtBpT+Wbg8
F7b45SXAP2665DMO11D8mmRKOxlEA5ve4N6J7Vrk5ScSyZzVFHdCDtqk29gwE9Q85hsLYZBLfrbG
0JjX4EM/+aqKLdvp6YiaG3X0EujfbBM3Rb4zKvGvnb2ApiLXGRyjItZBCSorD07gOiiTli0IOouJ
KEB1CWvD5+jt2P1Sah/wFH8lAn8KLhtShrID0GctD+kXHWOfQhDnCP79E9FYk5FA7LXsWlr+3+UK
HICLRChklOlOE27tpQMgyVmBEfVa+8yvjf2gfc2jyZ0hMoz+jIrmySfvt+dbOM0+QwNTv8NUCBc8
hCQGH/rn9WoLrkli57QdvY+4c+9UncwObEJQ7bJDKTaJ5OeKoRkh5y3VSDtNNDSTjlcqpJEH22bB
ZGrwBvWhaempzotJYeYoz+LrUIXfs6A1aYGjqAtfENv3MdRZzEIfkaRbIQvikEhZTfJhUdgZqfL/
o/2XYIvGchoXwaGqleznCYRRefMlBu968s/lDNcaeAKLq8vLSzaouQApMWdGZjQlvjuqqy3qb5fL
am3Ttqd9M4t/1kgEZzSR7cgCU3XintWVT5hIzg7pla3vX7tv9s3d1ICb5X84IzYRap1fC3ssZaTD
H8S1nypYR5J7X3yZveWakN3UbZWxl+OWWbeNGI9BtNZ1NyBdaNOvJAOUCcU9prxP597jHvIyxwDT
knpTMRs22F7aR9CCc1WJAtyKEXyCL0DXpDeNCIdmRhV8M81wvwsHLWtMMe1k1tMu9nr/7qoezCUA
yE3VX4i6st3rh51TP5+o6zad32oT1VufQS6ZnAh6fGFcdfKgi4VfvGilXX/1lIAWtEjS+1UZ5VV8
xudXKZmCpbk/cZCvL9+tm9EPKGVO1vBi1yE2OFHLErVWDSd6YdhfAIkKNGpkl2aC2Mxo2Gsuq4vl
C2d6c09Ya6WJX+O82e+H0RniC9NsAqs0ruflfDfr9MXr77NqcRulKiuMWQp+efPBr99AthOQmI35
OALT/KDeLjVYldAuIOKqWeZmke3hmQdqeRwlh8JBerKTfslDXrnCA8sdAiaVJxe+Un90RxNMTCxg
w8N1a+yTzcEMaIBLmNmuG4GhyO35YnGUYH1G1V+z2/vG2C5Z1YPyq4shdU79i/4e0TZPptH2TqrJ
QAZt0muRLmF6Cloij9ygGjdQmwM23XT8yFORQnoSN56MoH75xEfMxLc3AvEJ7z8bUAmkVs/RjbgI
9az6Zz0ZR0yAWkraxMNwK3MSJt+zLZkh+mLai5PIJCeUfRnWMgJej0AkIVakG+2WQITo/cUO6HXn
AOGSv8hAZ9vJSSa/5HfjYhE0fh0aVuCno50bDyEppdvP0bwN/5uhLFeJQ8wLliE28sxD1XQR2G2Q
GhR9Gyb+RFr/6liDS7ENB/UEB6AYmfFnDYMjeUwpNFKAAMbYB8YjfWVIVtBKJHeeIIKiMnVPsrtZ
UIIVK+/dpn3SEAAF2sJtl0Y6iPfRepZdQp5GOYE0ctTjRhODKuRzcbWrbH19/ppKlEZ83a09ztf6
F7zItAkzVrDCB42m7KV0gAMqWGfRoZHqbebIfUqwpja39VU1rsk0S6OCGTEAF5yJnGw6av4luD6m
9VCbBm5ZpHQjjcHF73mHtQHezPorHD5g2NBtT3R1jib3vZMJC0M/YTNBznhtGNkKYuEYWojSAQM9
+dfmUmjVX/eyPU0i4vyuwaDa0bdUnsEv+XLW9U/8OB27jCgGS3Cj8c40TR35c8Nlb9JTpa5GVMmu
ywy1aHNkhaObHKGIeYJIZtKehdFthL4CPoppzevbBOpVNg0MhxWXSoVo75uQFinfVn2rTMEPLDMD
KSn7n/XYJxz3eYVe/7KZRDur5dvDgznfBLcJFMYUbBzTKadNvJ9QsSuJYwD5j3DPrnegmovm6KuR
nOZzbRdYkURRmLbNMVqMZeU88K0nVaPZQdvZHy3uMfq1wafXrtvjtqvfCqQ6BsLJizmD0CrYHb03
6zuaBBj8oj313B/eMugMa3yYfaMWKomFlbFTaCuHVWW7eqP+wTWg/kil6J6hZj4DtRQ7yIWDmnMh
k3N6Qa5Sw7RJwoXDRBwFI7v+eaUV57yaEB83Bl3JgRL5ptdP/dHsZENhi6a18sR3CWXZKgu2Kl41
UFP2PosT0YY8/hcwfsfSM4EtvNmZwGPiDpF8b5M7WB4F/SqyQqSg7lkOar2UmuaEcP7Ke60ISBP7
6NNeHqr7gA44VPjYw2FFpjJWmJ9fiIZ8RBPhIiYw18KZ341B64P2e3tsFNnSDcBrjgv+PoK1NUgQ
b5SLzHwnzkPLdt1Ljcv9/1FirAZ3Z8q+re8OAIapcF/m8DiOfElMCSzlWzG5sxAks5MtJi4niHO3
yQrorU7jPuBHarwI247zLrNEHOz5nk9RTPZtLw6jRvjrw4Sf12oPI7qsGtvbAcrQlq76V5p5F5CO
63/qDpdI5ZjH/PdGIVPvVj40sSK/c1N2TFSrXm5k1BrbOyqxMvnt1sp0wh2NXzTtHJQLg/8ZxQtu
3MA5eCkSnB8/WOkJYz6IORB3ayIOaAVeHDw+hkLd/OUG/R7OhucLO0W6vmcbdnINMeXAMd3HM/lB
HbhmznNHoDnZQmB0B8Y1CGqUBvtFKqpKY2znw73bRHHvOSZNJcLu8j0k+p3Uab2nS7nvm4NdxPGp
6XnP8JU3KgbwoooiGuR014gGDhsCJr8guN6q1c15/kdW9Ptl5yzBh7p4IlQMkxxbOlUoqKS52em9
FIDqwFARWTCSukh+OoxO6VFv4QArdYv1FF2B09vaGeqs20q6iDaoOPGE5uioQmx1hCxURirOmxST
gN4dxWNqVNNRjwQD4WB9febkxs8Jx5skhgvWFlTWOE8c6MLeihskephrh5MtkuDjFwyit+t+Minm
P5PIrgXP471q9/G1H6C85j/CN6YgL7pW2WXjPuAlC4OY+U2GZ/3//cioP3v2W/vAsmj/JSOwN5a3
73/kYyu2/FTuZyA6bqH4CJ/jaopB27hwhjiqiGdt1E2aB850Hf4ayPT9a/9kf8QjHRePHG+XauPn
mrIfxFWgk2r8t9uU/xtVVC2nttWBeGLlw971wcdIUttV5UJaGU2N/fWxatru4Kkr8snizJsSqy+M
Xe1n2tl1YDESVNk0WqmK4zd5baXRr4jnK6DAXTkfX2LGD88z09WwyQEhD9qdDI9FxDr7AUEGCxvr
nARluqcgw7kuzk00UY8M+KpQ042UTWOA8eY+n+TZG6u/mQO4+G/RS3demJMLkQo8eQSKRUeyFyEU
evvhcXePCK1qzh/0hF5HUgTgqlspNU0MjD2810OCnFg7zIAVREN/SzXX4+KNIGU071KVutPY+Yka
ZaZVQsVzbt0jQaIhPw1jGMo9ZAhKo9MyMklBOA6pbgu7vFaCOjjlU6kJuH3v8aPsZJSwXeoYagOE
MrQNBSpyLp8F9h2g6Dt6zn4FYb+PuBVV/GUsPh4/600EhMriRS88wVpwa/ZMy9Stz9feCf6Apz0v
hYo7SLohEblAEXvZLsbFgcbhvHhptWRlkLuaf7ggB45qFZxv/X09rDXTmn+AEXNpnaPPHgxiy+IL
SfRucgRl/c3l6VL8uDrRCACmYjpqKG8fj8fYInUONyuRiWnIqLGnx+gxPVVjrjDNDxt4mc6zWuZv
HnlURVOYXltefpKrBLWKMS6/gWZEUpeqapjLvW9YvvH5w7JSmKaOgsWy2Img6DahpaGKg0UFf+Vg
l0BQaP813QiGiAcPohH9CcxtAgk9mgs3Y6WYbUAEQDFhs1Q5mmvh5tfxyntgRlfYBXfhmtOv95PT
q9jh4E65VCI/voiCZGYFY7Ji+6wCCCT+iJdbTFUtY3ZhmZBehaFlsWqXUnCG/q/ptgas+2/cns8+
8Qj+eqGc+KMc/dPIch4Qu4ogbcfA/mOnZb8tVhQzqryqnhCgSJBnl9eiEETxw7eHj5rfOTUSA8c1
ggv2OTu0Np/OKkqAj8Cgcdi4dp6OVUQ0wcXKpH1J1PUfwjtZIq2wCoxFwMwvq97a576Y02aASNZQ
GU1vTnDr4J/RsT6t6Oqjks2RgimmlbnoWg40p4HgIIwQSU7Vkfb8h028tlwrg2hnKnlQ6DBEhWYk
GrXIbbXioH3ZRYrvpj+bLZwdO6QIqkU29WGEmsER2uq6fKZqQ4B/qIjB/+MwAlOHDn47JybemCyv
+yB7lwQ4qvUqStvTawUfTq4TsI2xhDBNRTV590ADgPGSQ9Q15kPHmTYxacoCHETCMZihnXjZRZL0
GuZaq7CGfVsDrau2bmB7JFZj1Fxux6dG6yIGFbFgIwfxRnLIOsKkKnf4FcmC7F6Z42AhwVeVRber
znkP3HKI6S52idDaD5S5R7T263cM9HBbEcEpTMLTPfCYrgefBW7jsNWdRbZNJfrhB29nkJ1p+AQD
yf6/tyUQLDb4aldJMOtI5zX/9LtrBCnOboY1K4S4qdvmhp7F/d3JMWcFYkHc4AI0zVR9wZcV4Yti
YAz8i1omcckfFsn7FC9bnaJUA4arPvBWUwY0SuGle3B5ZL36alsLL6nle0oj3aOkaNojLSRhpjod
eIfo3LqmrXe0fLo/3+JoMUlnNSup2h6JlAh7YemrEC4YpLqd4jwiRlKAknKzWrCtZS+phMoWiFPi
l4JcGhUM1swjCfoB+rRqCswwt+dTusohGr4IF9yWlyDLxvGV8yrCWO2aLbZhXgzeEC2BtnZfohZX
lgnlbrTTWsqxK7NiKbOu4/q1BOjF3zEnFnowvNSkFrc4R5Js5DlXundFOqSlgOOipO1e1BKvmMLD
JAG+OejrTqcsALIzTudovwNjtx6wvVm2ZkFtjp4v4bufavAlf+sY6zOVzbLhOKxHRPjfqKOYjAbn
LPfbfudR+NW1IFhS+acZ6WmY6P/cwSV6WsngsdVcVa6c9kgyFunvRpDY106rJLbTqjYcPYon17Yt
CLeuIunWxh+31hBcSH3N1BoSLgC8kLCv5CYzBNokTQ8JT9jqmi5ue3J67odI+0sR22YCIbN2sL/w
5IvWxQLS+H0GUZKPyjtAXefCJgVVo/J8dYGDX/YUI/C9syNIpagDHM9n2FmDrELBpM4a6K91VgTJ
v5zJvjnFcaCUWad7bEH9EqiC+Wu1praFfFdNZgU27ECRPBFvxATpb+4pfBZr1jk5GAcEvTlaAiZE
jIydgvG3XR5Q13cUW7mXNzxTeW4a0Uqg3Iwi9LiexRvteCXuHAcGUpoaxH2O0iMgKQXrFNhcc7U8
bSPnkhCRm4KiebcKb/BJDNNU5tBTKPqXNJQ1D7sJuW0R4nRgfBtgtnIDwimpwSfAEyflYk5MpxUh
9/kZgjrLjyNCe1L7++Mptby8sFAkt1FeKbvKukH7ADtsMLwe+FRjc/W+nx+nDn3ZIXAg6JoQhLYc
6mqZS04p/JL1bqjbX0nr9gRgJQIKIxw/etNWG3b0wZYtW8UHIE56LxdFWfD11k6OkAQix6bUHG9D
UmNHv6nBqelppe7CncwRhSKsa2DP5CuloEKysdYPtClbMPXG41U5Eh3Ejdua/AH1c6X5l5V2KxDz
+4QXtz7tjfXnuSOc6yk+aU8Gx2pId3H3V1uEWb/0jLHG/2uxVo5k0AERsVOUhmsZwikqQNGDvANX
6vp2NYCgob/Pm0VJCOnpJdNLBf5EBmFBAEXEHkHvGL8pCQ0Hrl5BVrSLOatIVfRSWxq1KpeocLRk
sjBUQaROr1TXLfgdPjmTjjUyEkrQdPksvIQh772CZSTGqllGIjfmpZ7MkDfi7RDjNOm9DnRJxyAi
jQP9ogkzirM5DmRQseyYNnnZgGnWdc/ywTjAS7KZ4IJyPQRhWS37fu7k4pfNJpRDu2owpG6XCKSt
DsQ0JmLJlNkNHmlYUbtrJpQkqK19fRXWH2C4wKtLeu0Ua8vvyRqtqCOW73ph986c1Ke4lE+Syr+J
GP4h1DNP8c8KRrWrkdoleNM6ZJ6oFRyfiPRbZEoyKL8zH6mp9SFXset7zTw1QH40qhEJ0CvHoOfo
CPhlTZuVl5O73zJ35io3DiFhFYbg8C+IjSGFMPPL0yUAART3zyDGYBjWxM3b6j7mk9H6gZrFsfQT
ajeP1aN2EkSRCFAJbPgSJuspNJqmgiTqqEfGNizDiFrHJHNP3Q9gbbLXsDl3D0Fr7KeS4g1ztsLE
T00KefRkUkqwESupUm/0vC1CPIp4f8MUsfr5H81GpDPkyEUqFa1LzzItSzX8Jkm1HIH2wkrilL6k
vJHXNHc8kE+rTvUOuLb7M6qsP1M8hKiiNZ9fpKveaUGoRmzO5VT6K3Aopmmigdyu5My4k4XPjLoL
rrM3MlgWjPrqxIp+rUpxff0IL/vZnSIipxiMWuBsIXwR12NTMzp+ZPOS/ZqmlD9lTPqF0odlb1JI
RlWOqveWJIfVn8O9notVh2JKU05iNeXLQ+Xa9jGFLOqMgwP9ZvwvP/IvZ1mQqFCjl+/HeEgNy5A4
8Hsn/7xQjMdbXXYTp6g6qtlYekKhXvKesHKx3RvsaNHah2HUgPkudr+LWbn0+ZC7LARdqarR0uKx
uRPcWFWJQWULJ9EpMzUQ3DbXcdiBBvfr+Yn00gZZeYIx38dcXBfpl3U55D566GAWjDzE1LIsWpfY
grGXQSvGnp6nr7iP89GDqOs5npKMDEsmzjU+83Q/4SmRF4zvNG1AUJYmiYWYFiVRBv4F6uPuI/sR
+YJXeqPMdBXaojANLmi1xhcshKIQgsgTGgCj092vtP5cQZ45B51vhc4fShKoOvEgphErfncbpgHH
/FAbcvNYMgFPgPIq2YgH1FlIUJVCmbymyM/U6Jidu0EkvZys1J9uTY2qCIk8uVpJW6o5rPEivwF2
QUpM0EbHjjCAG0q1PKAIw1mtWRgES3bN+ShG21gSv3RcHczwzzQ5Z7M2fHzQwoQuYX850MRjxXUf
VjdSpOEZbuiWAL+UC0cdT5utivnhEQndpWW2IkrnhK5oGrPHp5SStBoVu1cqEt+VykV1RzXQIJGp
58bpJ10QrjWUq7/GLEVxua5bPyjl8kVcQIY/xShxiG7ltnB4637oJ5quH4D3d1SRsZmPuMvWn20d
uKQdPcW+m8RT3MDZj4WqnlQgEsTW2zBiQjb3nXQSxfbRU+gpsPhWeShTYjOwk3pQC/EVs/w4pBEA
DMRsGtZjov0zk4aI2cfK9HnYMahotD+sRLXXrbLzxMAv4I7ToeDKVnab2DLgTsENStuKStEMMCBt
n0vQp0g6494HUQbAoaYU1D74BZZbuLSv8d3rp3zY9UqpK5Uhr/7V+KYFUPN1/jH1Lf3s0JL0AETz
70YOENayYd/pRworfcrvqFaeE8Ztj9EkSsoFyAEhyHDMHIa86SUBtWN1LKrbFLB5DYHQEi00K3DY
9id6VIXrESRwvv2qNIOd7KXHo+MM7OCFSaunZqCRf+U0J+AzD81NaTRhCPcJB9gs1zBRs54K7F5Q
vFYYJQNSX6xHaisncs4FGlt9IdRvIAwq4/+YnOdjAMMVbtDJK2CXtr5hOlNyoDrw85k/nc5yD4AX
Z9WfhhqfExaRxlU3VeBl72MIKJ8SvkJdg5g0pUct2D8dk/J9Ur2/cNntjM2IjUAWQdBgM6Pdnam3
ssCPWL0YGj9ZTvamT8x8NPRVN64hmPIhLKBgcbyZqqqB4irgBmxVVTUAmhi9LBC4+jD79lRzNx5o
Y8un8+i+oE1KBJxe1qnI8ENcp7X9Xie9tTwHbNz82wLddtwY5TgstKTejKmCEBe6U8XdUp2Sfcqh
cHmLKA3MWZoep+Ecb/M/yWwQ0HwupT3OMRV2Fl9IsWTIlS/hnN/a2yDd6bhSUFWPslny55URSpLT
/qxamOpiW4f4B+N5tb1rIKfg0aDIGtO50H/UxJmjzw3KhZ+3avoLzZehgYsRZaKmJncGyoxvV2Jw
MczTEquMvrw0W3ESgqO25LBmJQM+vlwLK/HTYZSXiJAY1dzpQY2gwOqTYzp+3ykop2/892R0TFqG
+r401y1i92fVOEIk2O0sY+ERm0VTao12xlfLnBXuy/Rz2HeHh4dpjirTnQhy+IDa0NZRp5rG9hbJ
jsfgjEaRB4lLRwdDVi+rXYSh4SI6AiSUsy7+CI7X8wzHIxVpm5Kgjp1yB5ITeUCm1naEakuDvFjT
WWIso5hLRjNTlpc+ZK+Yq2DWmockWy15BrMmV6d4tiQov9K4ZJkOPZYrzqbUSz6OZjzu4/zoua45
0zpHno1U4xHYnnSP4e5hh/mK0I7gdfRUI6NJ6u4uIyKvxvWncpuWd1ERJpuiU6GHY3Siz4JvymxJ
MljJsBm0X88sAg0tVisbnUEhF7xQLRJknhC7hhZO886gxI5XEQGVzpe7lJ5GyIkRW4e/H028ytuD
A3VaylCRgx8YGA25BWnJCa4nCqcwB23fOpH7o3qgIVjkRahXHWSM/E9u0qU+TH/8CqWDjspJ/4r7
68v5eRUVQPgU8e4kB7K596/GAsLi6VpE5wgqXdM/E4ei/7E/TLNpj1JFw3BY6AYOAsufXZzYFU1T
zxrqR61gUayAOP7p4HPZhEpfjWn+FIPMyO6nqNl+/Kl/F3BnQPkt2DFpgqdFCRFSQYvG4FWsajWV
KbjB9lkHF37SgwWOJW32r0RGSEqS7t6AOp+Ddem8UqkmFffE+ef4y1vAfJ9Ogw6Au2rVdv0wrOoE
H6ZcozIvTNWQfmEBtOhKkAq25LFnhDn/p73MPbLZg1SOSS0xPPsDdgtFTI/sb4BhhjlxHJDOUOHf
I2UnADBHfCV9bGQ+310F9VDM2dVM7exROozVkgUAQRSyBsbZu1nv6xRXma8IAaGFggdxvl1A7Rs0
vfn7QLKdFMzGuL0cq9e9htPWowZdneXJeAF8CFiUiFUBExUoCvd4hdz+FzvPgBVz63wgQwfQxtgM
R7cMybeLO41h85l6tijZdoeEYT4cXIrRYTiz+Nol4htVNjZsm3OciM0tRURgobEVbE1Pjwo//0XU
CzL4kfVxXHQ0WkiBp4BB23toSgS+dSSCK8MlTUVea/fbY55wu+TL3JXXN0XxH6tKKoaA61aGl582
rn6AIGydeXXfI6pnHSz6tj0pzM8OfW6O+0pU/C1fI6C5RSNOp1KAH9kw9BIpSiWstrRqONXcj4ju
zvHewr6i8OvXADbm6MSX7cZW0nJX8HOg+tPHuNyG0FcHvOkY0tcDQ3OUNkzPl6D+RT4s05jtAVg0
YnKJ3zySnYSHXAoyW75jE3A6XoynlS8TXcDweW0GIMd06w0z5q6DevjbzewIFrjr8be8G/vvQmEA
sOri4cnWAs5OLmaHQEbR8aZO907Nra/2GflCdxNrTHgveiBTW0JnLLNa9bcxCz7TW5wXIa8u2dEo
Hqhr8nB3H+1CO6yHep9bbUmmjOIGJRkLsxsept4rTYBE6tqGiNPm1cmRwkyoHcl90UuVEWdVmnwT
edqTLdMiV5GNJYTgmC1/0Gny1jI3D5ncIl/f4X6LxYg7ohkLlfdlVVQCl+CBrOQwx2+unu4ibZVN
WdNIpaAR9uq95UUkm6tU9GKyr0ERny6kzYIOlWYgzlfPAckt+lVJuW0T6kNUDmXl1nLDIfqW9zI5
yPZdfOJ5htHIlYVcj2/jMDsrZSb9JLRZiGYD8rIIf3a1W1PPk2b1hZmv+FlenjIWOB/yuOkjt5km
S51dO8MN+Mc6MG3ikKwy4SngNhP2jutudeKcHWUrJ9bPdPvQYqmHaKfzxeS2kqJofOrMKn2a497s
+mq5xF0FwspEgZdthOC3aPDlI5i0aSw0GVJ4kXqhIcxyc/ZOHViRc2p5aqDoKuq0txNYr5e+cQED
ZwZdvuqre1+jIbo8v3Pt4Y5mBj9HXzbcKuPI2F8RXQFgi8gZdA7bR+3wk2WpLc2LFo6yHXgmj0IX
jnk6kEaILAn5Jei/ikQkC6JihW6iinOmgeVp2iWJOoOsk6u3mUsOeWcu7zi63pTDQwhP23MSypL5
NuC9Zqz1wgWa1QSXlgTy2IMinX6YFtRoY+G0Et3u2hcWBajAIyDOYJB4e5bWns09weJnwwDHq5Yg
8JU3SWUltj7jezlzSM2HBCOKvWnLy1dpi7Ksw9s0kjbzpep4dS1IkQbONDC3neEBY14gKXd30WRy
m/OaDych0d8frrCwdusLNRfBEH61RsGKZmNl+GBZVht0d9HsUCWNb5mU5oa2YbZDaV96YTCG0EC3
OJVjMv0XRHOe2ViSeh99K8A2ZOs+RrGBh/9oCsboP78eJ/A3egWvZ+WCo1xZIfBfpsgUaw28f94U
c9PMxVcCWdFwNiWEMVW5wSM5Rl5WpL6JUrc9ZFZPdUzJ8FQogOgEXWKFj8zNRskcLYTA7sU7Q8Cf
NO2jebESoUGt0tD7AfPjUzlv3b3EUQisH//xwMP2BL0+ZeauwIXINXv7Xc5s0wvruYXkXWNmGDbZ
TMvQE9SH13/D91io39DBJHzq7Cg+cJZPeYZCMPSzpvoEB/Zy9BfkwOcT2hcsZ6/BaTgPeEU1+Zly
rjNvMsjrvrdpRTnh5ZWJrO41NnQ1olnMRZQv05A6qiJIlEwVGU1HqF0bUAi0Nm3the9KSN7UbF3/
6vq/Pp5rSKD3YEd0zfpC1MgJuQC+K4vlOeIZpvoLp9v0CZJC5oLu+PZAHJnCmhYrD/4+TJS4DzuM
racZSRSoC5MJEmPADJ6vbCE5sS/dDCw+lDjNU5fjZrtfmYEg/EBfRW+pph+JyG1dhFYa2F9Ggfpa
s1sYSNNa7Kjdw0BAIf17u3Es7c6J9oSo6bLj1jrnrzLHeEGDkeVDfhQX4wRLa6g42/3h5LbFuhOz
nJuSpRqSPCRKm1r7QNJFh9XyXLdmZLqOTOGx2tT+Y9lt9wgeBXW5Dt6aOmdFftExmbKlUOGvl/E9
tDSeHF1mJtjo3Wg6h89HN/+njryaR12xbtK6hu5ZfBvaIa9OXsh7KiL+iBSERHWhI93z6Rlg+viP
0T43r5h28pMBucrS3KiDb4jd1Qogl0RK3X0u2NqynyogeTQinMuJ8+hoYn0SZ+GMjpEVWPxRf0km
q7s1NGNc5kjo2LlAqAW0bhLtwnAXKKoiiB0yMZtxfLSMYxwDmMK5hWHlK4OHBFpbvla+7Gcyc1+M
W4C4UtoEEStvXoPFXzXOj/9Eod6HnOSiEDRR9zpZMGPlwNtV2hjA6W/ClZ8kOyoZbrO4Cc9W0eNk
ydTX63uCBqvElWK79Qd090m6FYpBDzXpMY9ja770Z5zW2VYaBDVg72JtlrfWyqzLovjrqE/8HNVq
awymM5urZ5AMZExn8/dbi9izc0p28hQq4e5UwfmJklqnBpqy5RPCIeSiumhM9Drwy2LAJebYEwjx
Ka8dQ8E2m7d1rw2J95rBJ0E+YQTfep1/oNaoS6IQYvP8qdnO6kn6lYJOt8diKbCeCucvbPHvQ8kA
g/XcJrbUIUAPKo/6oHBSQeJMu9WBfaic1HCQ7Abk8i2T6V38cCr7C5OCRKuKasR3YRhOOzd5PK0j
GXJVfuMQYEckhYjQ+zu2tkTnOe8PxDzce984xGYhq3JzS72Or9fjxWhbLyrujFE7w0IUhqn66tgR
g8zPlzXh1DwVLRah04zi5Lg2rQVm1JA3+NrYt9dCibjJJ8FBALG68FOIUO+X16j7duVE91Njnbjl
AVeTAxO+YOF9yDjI3qfIbHQ5GmGL03+M9hoVSX4OaKbJeCEgGHgKBdgwOq7L6z+dHkUcX6IptnPv
8HByVomGHfXtdq/VHATTgCN3nBc3XbVs6U3hPV4s1XQuufPdXXHOfWQBKqw8ODXNWlrAs/tl+DVL
2k6iEU4C/Y3BoIf/rN5VfWxl1PjkgNwvcG2vTNbdH99Mw+tpq+2oF8guajdfBxHyNqYseogTCBYD
Myvnz5zONup7BrG46GEtHKDAX9yg/hkiiIYZHVUMBKL2ZVUDLY4XSCvq9ImgAnhCst+ulRYkTi+G
+xKVg9uZKPcEpaGlYD6zImqjlykGlhjNmtO74sFsAujPfpYZswGsAe2fvrjyPh5ul/OpEr4H2xHf
4GFKkRX5VnvOfXfUmGbMDTWaQJH1mm153U9vmYHPAcQeFQzBdg/5ESl0ohOPn6DTxxNUHfnXKnCJ
b6RYEZSHSMvicc3sCqOKFm9RDuWkQcmJSqCEC5U5DwpZ0+tkwnYcrejLK/+8jbUKylBA0wKp5CEl
L3vxjTHmGXsW9z1FVwufA7rs6q/01WHCchSXwU+ivx8equuf1c45z7fwFH8CY3KoP+PqjGNEfX9O
Cy3fRiEtY5fqLHC2v35s7tY8sjz/HDV5/IUoTkRs2n0Ls2p5nL4cYHNPuVPUpDR+Zv3wBIMxihah
4GHXFpThLcV9qlGazFGRNlzsduxftbK2YgxZsAOsVEA1089imZj7CySH0+ddNNYp2xc5RHVIYkn/
iTz88atpkTyDbOUabBtUnXpn36FNJd7nG8MXhNRMzbUuWWz4Ogp7APvbGioYrIehgcY6M7q/avmp
6rcSnxi4qUc+mCvFd06hct7KGjFr2WcT0scK7zRYOaD6DoTmy/3RbsYfYFJdFGi48ahxikzU6LOc
unyE/uEHXSkXh8tD9opcmAIm1w6IyTGcxAEtPiR/qyoj1sZGruPzulWr4Vsd/uJqNM4AkFcBjHvM
0ibItz7+uQ62GlPNlriL3Z6LDu4Hy6Watg3UuCEAr5YRh48lReCeySy8e+eTXf4srldVA/ObDJlT
QncHHdRDB51Zape6bIijcSxFI6xPo3XGlPm8kgQDDlfrvTclfwydsCAf7IRR+jPoje83eBN0UH+s
uA7gmREvBQQGOPlNQZ8ylqQzfYjhj5LktrThhAcPg6N+Z/DzWZFJ0umYWXu29yuoEj5HkJVK8+I3
Fgch3gZRxBPm5p9UvdhnNuB4xdfYHsiST268GGhJnhbMa+KvCvkaO1umkZKmy7TUrfmYaTg7qLXy
w6gBbufFw0rln0fGNh7KRh3CevnmlVHl7VR3iP8E09/8U0q0DhhFVxoIiFCZ1Lj0rj6uXLLz/WhL
yqtwtbQk8U+t/Wfo+hEcm5oX21Qp8DbNGqCY/qiyB+oKYvP+QkTQufznq8vfjdkkrNsy0keDNTNX
Dn8tTdMx+3rtxqNLohPLFKbnZJnw+ixlSJrkoZQDa0/Zf+OpzcLoaAslb+5ExH01gax0Zry1i5hq
T2MXJF10fSj97A/IlauorlshbV7Kzl5Hr8lclrwCv9a8hlVtTlp6hFy6y5NQ5xs1D24w4+/b2A11
HDaeOq0XCf1sIKYnOh9zh6dJqlewDIv/4W+tQtlJs93hNY+9kUJlV2TMJ6oe6WJQypuQFLmtLme3
uOfnOkuYqrHHc0c3k99xedgX1EFnA5PiMSOCKxf8BaUV26TJEK2/zYEeNxdpaiIrdjoWMAz5k8e9
wfQTvG0ppySIRP4/mqdXrkLz2csfXvbFcoMCM/dox6LhsYNFggXS+4siNIHrXOw4fCInJwjBOmNh
KYAUjqMY+46Xvl7fdkLp3JvJS7jwusWdzzULQgGshCge4FBil5hzKfEnMnSQQeUi7Y0Fwh5oq1iW
3mXKqtnbLhDwwvzP74gydHm9Ns2h6Hpk/Y3AT3ySGJJAlajGBOYhdii/1IevBpdmmTQ+p8sxVY66
0BN5MrudO+DaUXFf/mIJILLdRAwTe5CTszZaWaAP5oznFm4cjkYILfKsZThSOpSG02pbI2kHx6sI
l1UV4xz0baFIqCrgUXkZYAQD/XCNfVG31cKF+RtY0wTeMbA79qglMCACQZbej1oiOsqz1l0Mpl8E
iPoNwVWZYngCmNuNBPehTtoJ2dulvckG8UL2y3dl0zbAK0mHUtZQyYeGBJr1pqtzD/3Ums4OeWuA
q6+A0ahiIyamXs2Q691NCFlOZWkt0xtO68wkfdmyNb9JA3fHIzSWad3OyPsXzaybYVti4dl14T/d
AKs3px11tf8oV7n/Ji92vWIdX8CkFJlBIIFzO3xfxH1oqyTixLy0coIIYFTJqxU54kfThRztN/Ni
5IYWeXX+VNQjyE6Oiub/nJA86TP6b879Ne0/bhLTZvrAAyTNu9993gzVUz+g55NrcIpuGpOo8fa9
3A8A8qogzT5RIgMJjwM6zef4RHRjY+40iToSCZm6+dMYmL1WF+j9lrqg/T5Y0rXOjxxKqLstRHAO
ik1IY5AQGLjJvoo1eq3izgL2v4rMKZL2a7lOM8a+Ye69YsebIYOStfEhxuASxP5/XLKN93T0YOko
9lGkTlvgaMowzibaVayCHKu/6osSlTlG8HZ/KaA9b+Jtl6a5ZTfEI2gFUdXlP7DWzsh8jpm/l5il
apKo1EAtL2bgvD9ieoXRyTqtvF/5vhI9aVjPzXlznz4rMqmcC/On6CjUrBEIqPSib4F6F9mcVZzS
8jdqc82COaSvUAQcP/0yds1fpjjklm4TZQuZ3T3Z+hvjMCA9uEMSkBeXPeb8g0th3ljNIJlJsb/t
8flrmtW9cH+DJwgSAd/fDE0H6lDqX15ahVnyVowdh3ESvHVDkdyCv/jUSGrE7dUORirq9X6LVPos
U+MmXXE5VIyavmAtYTw1T+/dQ4sgwobl8tIV1JNPjXgpcqT7lZtHFQQ6J28Z6YoHnor5Ig33gXjj
BsHjhFNWIdqraUo+h0i8kpoZxxJWb9LTC8k8poCEQFsah/rDRcgH2ThiVSX1ER88I/h8qLeEsAbs
jUZ+P6ejv07J7K4gbtORKKRmUNTRvrvzYDSNZeyMhzUxVil50G2qlUYZynErMuIpY0qlc2iS4re/
TyygIczWxvDO66OxFUlOV8A7z0w1Axt4nH6v/TRrqPKIAyyYbuGukYldgdEmkmiQIfGyyEM5qGiv
WULGP9UUR6NzemolgIUtdBQmYlDh7TOV1cSv9R+7DweydRsd/GlGulzGs12B5XhKzAFOX/qK/yA6
zyJHifQLNQU9kkXPqjmHRu6SDVvut/1iM+3ZyTO4my7QLj9rq7A7lUrchs5Imjh5R3xHpc7J1kxp
s6tD8DKudb589yQnu3RtsaF9fGVK5PDqjTjEaxlhgNLczJ+g9G3wpp7V7rIqEBvDVjiI4kULRV2S
yrdiR03ixrRvf8bXbCxXe4o9197kfpAAaciD+i8Vq9JhXKU/J+P0D/ka8ejg7PoLqNvMw2p99uZk
zrVc2pMpZClV0VXXijCO2KBlr5dbZPbbKA2tcTmFloaOheJCV3AMO2AqeLiBISMPXrsS64tz4Gzo
rzgKBMsRYTEadQdvuszSj8evgSAhIzUpv467CohjtT8jFHHuPa6sK+zV3fAq8wSrt30l96zkYUQm
x5C78ci26qVzNba2obyLmiExAJ+wUxzuyQ15uJrXOb5A1SRpfM3cFLxz/vvqf3i0U4NY85Dcidkn
Y/tXslTyJSI385unA0mEQshCuoS/qLHriYt6m6qVdpqnXRdrIamLHSzJulN0T/1BfJmY4bGz3PCX
0qLpzSRn/tkwOnYHm/TmLUATk6/4rOT6ssIbx0LR3y0hXNhvKRtrhDvz9uoIF/s3UsiNJ95pfCn7
Np9eViNrE0VRc6NyKl2qTIfqdkjVScr1sXQtxkig02lEYweR+sEAOtg4UOWF08F8xqCUgun7SCd6
WQLO7c+c80eFzmY/AEk3r40eJ5FLGzsGckcB0l46GvQAip7RBrVyvcw0+GuIj043ImmO9NOCm69D
tk4X1GgoR6+30bkQI8ZeJV+HkFvkMds72KZXWy5J7tzRczoJWawm5aRGM7eWv0k6mGGCyy2/QJ9j
Ji71UbjyWPZYurNOYwBp7iVFmItISUPB3W9I6vouuiSA60PtVMBy6zWW7lA/yirwATxkddW2d7Hq
K1GfrjzjbJCTnzUX+M+z7mVgUZZtOsrTQMx096WJBSYFfxFQ34xGQnsIqW5ZnkJlBKtbHVuCApwk
VRKBMUdSGPkrUxu8xfjGA5MfVyk1AGitmTjdwPJMdlmZHXffNvoKk6/2RNcv8QceSPXFMzwFTxM4
E3BuOxE4K7UISlwcKGjbcqF8nYfaS5zjoqiGgimp7PdljMp/RtnPPJNUE7B8+fNfL7dhSPMFyIW3
EcdtssFJDypKC2C+XwTtExM5pvmh1IQEDkgHwztiGCqEXDFQhr0pWi2RW2WjnmLNMIcGhhPkUL5l
H22emVxr9WyBcTG4tIMTf60YhJoQdW3y/0lc7wDok/2yBW0YkuJBie7xM1cCxHZVqOLXSd0BQr7j
hljz8COo+F4S4LuM7mdjnhWpcfzRX2gL7aDUMF4hxubDGTXRFoaAMzV7flfMa5Z0mX0EY5FFX0nB
tt2QCgiB7pPQnfH96CrIxESYFPZOICv8BtIikasi5+Rxuce6ZH+9TkWTbWfvMsFVQiMNnPvWKKTR
APBHYTYkDA2TODCS7n6OfLnRa2uE0SUvRxXLdqoUs1Ztb3ZC6e6y5iWIKfdk86kX+FhhunkDa3UN
fhPeGgj/88mPn1V7uvGS8t16JBUBvY2E21ENKwwBuiDme36Ct7AdxB3CiDjUX0Mo0CgSGpuY71rU
grEVIsy/dcLbUgdshQyLjT1+F5UGWOeYaUv86YjOwfvo2rCs5hQburm5cTZYKKKdifiEZ0cLb/Y+
qBhV8E+HHzREyq35EPm5WuSnDNKXkWVHXtvkj2XPFseBpWrOh+7n0j9k/0uePhlgb9Y4sZ9+GjF7
e9JD5somncBVCHFJr2+3M4dcw9Jb09ynH0vCYCca8uXxYL7B030aYFRl6n6GgUCQz77Fgw0rtnm6
3ZXZ5yyARUCXINc2hnQ9o6QN38SsINZx8SuQDBGPKHYZ9Up0akDyBt6W9+Pes+2NDjO2GGp/JNDK
0+33ZECjQQjBHitY7vFgQYZV0YAcnxgGJtyb3yxpaJJbMX+RCcfrMR2+TZCXSR3WAjLbNTdrPjpt
QwnOzHlo+IPoizN4LT4euUwkh0SCKn9+rXHag0Dfj1IryFtEWHSNfRaBfAMbAFaAuc0arkxg2/xQ
TK2JeZ3miFMm09dEc5Gz7Gm81nBhIzo3GfSu69iWnU36NIlE3gAkzVvT8pcORBtmlbeIPV3uYeIW
IWFXUPpGUdxZC4TUc9QeyPLqZiLwD0VFsd5+mF0tTglyk/99jz5ammABwDobZru0NtxttB9sEU6z
nHUaHxtv6bQUljzR2ruHSee5ePiF5dryrQD1Dbn00VG2YVoEf4fdga1zN9JbtccMYo1eXk8XMVFB
i8V0XOvaX82vt9POs6I5BGjjvl3E49RMjMd7vx1aBM04ijNAzaIK4BRmBrPD50f7BGNmrPJg7j6z
4VMm6hSHUXnLTxMFqw2gZ2O4tjRCyFtAPAgME/eWeZJOPyFaDCyl6q+UITOQp1QiHExm2hpCJjll
pRsxn1OObfPkcikOfiVkgTffEy5u3fB1tZrohmJ9QKto9hPjuKgEUSm8s2bF0ypUJq6QwnbfkwdD
2ei74EyiQOjVfK7vR6makeOHOT3u8wBfO3T6YqoA/G+Tq6+sjsEMpbuApgcs7LMnHTDygvVzON86
sRjb2kAPhvk1gIv5u46+4DhxRgQjZ54mTIiW5HHk3gxTvdBRAXqxttiqMuVXlPKTXTj1kDdBSRpK
TSQzx3SnVlKwppMit+AGu+/ojU2lmuCMcbTc2qrFjEln1xLbfXHm+/66Pr3cc8dJPoUmx5dCTvh3
VNMTehLzYj+3A45LsMRmdCPm0I3qsjL9EMrCmDRr4/S8oylmojXQfZv4HiMMgh16pzXUbZuz/4Im
lDGMNEcgwJegp025hYMGG2oPH59ObUZSRF64jIOE8UYVhpfdfJ1/eblUNGbT2MW+v2BLWh0LSRV/
w1I5Zuqoco8BAvWbk/w6RDGVI7TWAMRAJBaJS0fcGdhbXvhK/G7aME3w0QxdiXjToQiQW2wH9MNt
PRJO+b+aJ1pygQ4it483ftnc+VeeeizaTw08EFQErGDNiy1UTvpAHqKuIPKFPXsX4YTOGd3F1VU3
9TfI6qDAaatXG4818bwHuMKKjsLc924GOUUoGfsVSEcGRTXoPXE12gVUvwmOiURb8aLA+5mJYrZH
2HqAvKjbYaX8V0oyrkggDgmYChtBUcJBwMJkD/cn4DcbqEIZZpcfcc+GDSGtPWLTWLxqORfK8qQz
Qe/+U7x3mb7jKvKtVLjgMmYnkjgMqGCZ9EGSN8FnD0QvWOBIM6rv0aT64osM70pqAWoZ3sNhIuZG
Og61/82gke4Sm++MnUyMLTBkbMBE+jknpVa5yrON4YU5WPv7ySETeSpmr97KeRIw+zFJEqn+dehk
0LITa+5BswHJdDQbwONYIvHtLaoE2HV41Fk4j863/YkuTvyjI+hTotZBKb2eV7gyW09neBOQ8iKp
YMTcpcqCSLmstLWE/Vris3HJQky9a8ykrqL1hGaA8zlOe7Nio6E4WrOYnuMrJGksCZ5ZPXTqkKCQ
2s0Fgat6jK82L4+M4aG5b01ZILaHXPxRXZ3Z9/NOleoRYX1ruH1hJH58+1V8A9vwn2ym1Mlig4M0
TGKgCl8CXLVmog45b7QmVsV3EhqpWzs7IaI+x6aKvZo4DEi16Qmctqk8P75rNza37aNr3TgRhRin
5jKroD3hDUu0YoYYSmDVJJGAC8alT88FcSx6IfpPLjte5IXkrnVw44bCcVZg7pQgAdwXK6nLfoDE
rC19QJ3aPmFrz32Bks6dKCx4/ZeEEXBExZD7NxygVVuyezDRPIGcIBubJ88hdtzqP2AYgA+sHdC0
p2xVBqrMOiVastmpFOO9757rlIR7f3FFq/2iDuKU5SN80y6S2IGah3LG4QxlCj5Hpce3LZKUYBiC
2CRu95bB/c4J5cmqLepOWS8A6YIZ/O4CHDYgOEB7E+wnOie0goNd3Y6/dwQEJ88s+/QgSvlfl5PV
OBCwk1ZkdEClJ/l1senIYvkkNwwL2ydmeZmwLuZaVNO9FKcJ5oX8cRUEjKZKNjssbb5hVSP2zqyD
7HhXj+aVuHz3a2UuaNvDBLcMLcIMLLSylk/Tbh+LYaESnKEww5LjfDpKqjQ1TGXaUpG50yXtQCQq
7iUtiNIWnKQ4BXmYZxS5adNiOYERCQR94Iuj+91WRb8Px2bmxlsgCnrmUPJeGsUuDL1HcA1Ziyfp
vmTv2DL73lFPoR32RfLukafhwGHjCXtA27TQSpT7QRXI8HX7u3+b98zm5xGmezb5265x7UYm3wYU
T8hWXGSv6r9fcCKi/h4MLIv09rqSG+K5tSu2HGS+BTFKy9GQI3Vaoi2XIHidNErqJXveZkNcDJ/M
P6IO/EPld/h4L3UCZo1Yavp04fyly2/P/iCLG37kLApW/OCtJIBINYsR4QVYG2r/9N2YpbMLgvuW
tvI6+sSh+LTaRKd6m7Q9USIwmD5HMg88NjP+48UwVQonfhtnAofk2eC/aTg5WfC6Pb8FBGc4z0Rn
uOlf9pZxOkw/dO0/1ZatV/s263pxnUyqOzQb8kDkV5dbHlsHAJ/aIuUoPXGApsgQYQi/mpGwCtkU
JKRkiAvDnJ/ChH6pqZGtn4ldlN43VN6vtXR92PxE1SOmujOCMowTtE7AV6e+y5q5JnfePv/W2jTF
BR9WjInb2pTBgoZ5gn5Y2m+W4kQqg9pGQ910dj7UP3dCxwl1YQl45jQIfC72bMJvzJtxHBSDKcM+
KpC0Ys5nASEYf9vHH+I2T4+idp04zbOvZ8R3zpLSR8sFXRvnxlPaN7wTkS6vSJ5gBcbJ491yhxNu
E4L467AubJsEOVhhmITfNKGl6AzA1MvjT2W6lpcxEnshwqt0EfhjuAOVnbeuYA3HwN2qjmfuSrH9
q0sSvfp+6O3PQFxuHs/W0/qJaRM8Ts6w9fy+RM84hkyBJD1x1wSZzhELYpvswO0OZT4ujuFSlu3W
6jSGsy8+/JwPjHBv/DWjE4BQqZ5t5cCnh7y9QBISZr6eEtGXtZg/qPAJYhnIF6J3MDQ60T4LPxhW
e5ZbPobqP6yMu01ID+clnh+vY+X0XNLTHw7o8myZ9GdRielnEfgTC6ayDRxdic5zr0G6xcfCgN8G
7c3O5Lj2pVBYRPD2mk23Bb83fdldYpTbz0Yn83EUbSdcI702+0e5KupQxhF7Ptqm/8xntjWSUxyT
E9/zFrKuyOUfLnbo60fIXdcX8l8Xxecuh3ypcfEfU3TOFCfsdro4uU2LTFWJsVpc5cdQEen8xBkS
uVCegFwIcbD1/L+n/qWfRIXe8E1IGfGl9fWz4aGBeIi55z7EJ8b6/SdeXVEIxQRYMnhpqajtDC+d
D5ofyV6xV5fhRcaAT/fpNTaFevYYw7Z4hgaCkz1OclQ5lXRTMZzme9Flpa4DmxWFtq3gxiuyKjID
mKinsjtNfj2vqBjRnpRIzzB9XkfxGbtQw8f6giEap7jvCOE221QJtkO7975DAV0q33mhw6KlCatK
LXbuBwz/Y22NPuwaF7MP5ErLKZ/8Rwx/Oh/lEgDlv50fMzduDdAzuzYBMWZMFcE3y64o5kwZ5AlA
SXRNsq2l1gJcNiD0PFD/v+L3rHlwp9Jlw/KCUQy7uAyJPQn8MXzPzbmzHSuD/syf0AgAJMrZvWQP
I2uGP5MSjQeIt3FbGa2aIWE+i3nD5ynEN4pOab/Tqx5X7mp3UpPLTqXklxYFZiURgxdjuE0QNzrw
tIVIxq6GZJAj9xVgzw9/cwQ7WjbScgGqSkOPIPttIwQr59pesD1nuvzr3+u7kHIVBCMtWWYQkKv+
dSZosj0nK20aJYxyXWPm4sKrw+b0W20OgG3m738+XWuFP4kaUMPyiZRY1Nqqc+zjLxL9AVhVVoG6
0skmHzDJW9BVGVFLxlN8QUjZtSxTf15EthrDyv4hLhGcVvubJAZtZHi9G0RcWUwoKzrSIlw24EIu
CY/t1Gfbg+xzGOc9Gl0sznAYGELtjgs0Rt+n/ahIMqz5+2hLu2I6JG7DtNFj3CYyR7OA0J+awJNx
jF4NzyFKHpgKHbGovqz8q9iZx1nKru4uTPymFxU1DQJN1Mw2eWAM4fdAkYDtC/2hPYtkchPYRzvF
589EsKCyO53eVFwn/33wVJmhP1GLsoj5XyBraUpk5A1Um4P/F/jHPbGmxU57pwjEeYGyb89lhHm8
l9tQ44PEQEkkKxJPs/enOzT9ffGLLR/Kw8Dz5MIcTU2/vCZX7FaRwzBHvIo0EbuYwZDXSInjiz6T
NAh65WDov/yhU3zzvEYMuaWkJE3PUPajzKI76DLAuwDYmE3jE56LyQ+Zx3sZrp7aXHHvP2bmYfk1
p05b/G4aidc7iChfUk2ERvAGSQD+7aA6B546nDssT/6dGV1HnUogw0PZzQhNRzjUIuseXm0RulLH
tYTF9wjZTZM/+l4pTXnlolmbDcROSBEW+I47/F39AIPvyN6VcLTWKNVtmGXPG+IdKR1JlQJawgqr
M65yuujF1L1ecTBMiZgr4uQtIIJ/HIbWqjcy3x71fl47pUq/LEdZNPhcI+WEZNZ4I6Hs5/Bl4NDU
ifbhfkfD2QVkJxeeXDuWF8DCFhlh9Spc0L3fwRH31tw2NAyEBA91vDG9myjK/3NxtNf5EznG+KL5
IKGx8enjzPrjiYYZclXfyKoIdwPP820uupj8+R2khXQv4wD8hwrGCORKbMOisp+xg0WMCyHO/+ST
DsOigRNEy6Qajsg1RYCZVOIybkBlHUFVpn6NnNSljOlET5hubBcxI576FCILsiUupG3JtIT6JU3C
UsqMasVdvRir1VqoBojB+OUEtXLjrFbFEtbbhVXNp++f1pjSlKOx7FUixni/YjXPoCrNLj6418pf
iK7mZlmvGZ+fCBiPRq55XChgSpzQo6V74gTD8A8XskIy4mjp9dqEkWxkw4kZZbKuneOGXYmmFtEF
LyvqQmAzGYvaZwL+CiN9sj7XNF2aMks++7JiR9ZjY8MPznw+DTbncsurzltxRmGX1qHUATnh3iM3
gaLNMYBKccD5/gSGXdKakKP7hH/h1FZqlHkW8nE4AhGFtzJFotH2mRhyw/o3o245hgKiulk/KsRp
tpYaX3lFPmj6QNl93SKEOsxheLZ1FmW4sdIWorR4HqSgXPOMxsx8OLvuBBVgZ0HvDb2RsIqgs2D2
lZPgps2omSlRax5ZCOzGNRrYHPVoM4KgEZ2oAa3vHTRpWy9o49WJ3uFmcRHNK7LNfxnDi9WFhrfn
hvKvc/iYBnRiwdv3UFgatudkJQH4Ts0K+2ihCtJNLhDRUqLwibGWhRj+dnFfNr6+kgpWLuUahhtQ
EXfLJi7Gxf6tVKzdmvm/ZCpcfkZQksAMoAKoELWaI0QHPQVRAWpOqBXZdR+RnN9YLylusNn5kg7C
qX9mhkoisgRzQqF/7eWkZ9rR/aTQDqHFLh6VUDFBMtRbb+RAgLZ4D2EfEko3LQqjxGaZyrcboWTH
2tSjwgk0Gu4mjALKNLQqWVycC5CSHFndV39qHaucNg8D4m48rWHdpNkYhWKzlYmDHFhPgJiPEVfu
u4PU+VeCM96Fh3zSi2/7a8ZuIT8jdNLtih+gVuQBOCtfbksG8gZkhoUsX8Ti9poR7YspKFuaC3RP
WcuyseM+xpN3sR2NGKmF0P43NkpxbNixQv3s3ZpPiKpXkv1655MDeTOalievluFnkD0W4l6HCorS
ZyYYJaKbH4x2sv3Sr9kX7tS7zuJEocdrtRf7TOircI/89GVGO1/5HumY+fJAsjZURHOE27yS+Ue4
BYO7LQFF05kS5zMeRsL5TTP8O3DXx/fpWf/3gIyrQqyQySEli3negAEocgcs59F4quLc5GhJrz/C
pHPlWZ1m0fAmBRsmutXIyRMvSIuWE0UPmh3H3GGus72VJ0h+3dikKmWNZkxotkis60AgjYTJhv//
vXdXiuebOJjsYUqZvs3B4TdPMbGdm2wvt+OnFCVhTiv4atpi4SIbVRAw7waKr/GGW0pa6ugf9Q0r
CpVlMO/ehGH4ziFMg3Fa4eFLIBlomaDw4nQtlegGzOdazF9TcEXVL3jFdGFjQ8iBx9vVHexKd+Cd
FGUH2R6e9NxTV4shHZFW29Za2PdOUvkjEkO3+0nai7LShuQYRkB8HUMa1yF/DWJIVrAvau4ry8D+
cMZ63XaCVYOw65/nZlAAtsHI1PMn252Ie837bYPLBxI0qFineghBxWw896gDW4gxTNRClu0V6R40
Mo29QPYmqygeePlG6HV29LVJhex5KT5hMaePK1BqcWpZm20FtHkQu731jMOWz2oQFNaAZ8KkpeXE
gYdz1FLQrySdiUWOJfRrS21nu1vGS3bHscAGV7JQRHSrawV54kimX0wmwsUATrnSeuyDMJLGVqw9
Z6lAk9cG5j5fvXABk0y+TjaQlOJ3cMDl373ioshzcys8jwNaCLNxycaG02GKFvM16dRx6AfT7vvc
lCBNVSBV5+jpicjMIemoMb/PzSvkyHnt8UMNTut2GSuS6PFe+Lo4FVDxc4U269ZHTQ6BgaRmlwwG
NERCwKunMGKWpyh+8OrNE+2WCFGSqu2JaHxAvQvhY3tfQqIG9eeFhn95ZTNYN8zv+DNPzeC1wn23
Tcrl6cqN8gz4BZJfWu1zsrzYkB+rcpghEx+vNhc2Cz3So9z63dmF7VeHms481RjH2Q7awMlBlJ2N
9Ug1oSuw8B5u5GLsNGXTXMz/M5UcdziVoMNf7Yc6EMiz+tV1yc0ml7h9NHEQDMxP2abkeThDn1KP
oSVjUVd0iVAW/lyV8IKtk64OQl5mKJJDS/x+FpCXyz0JH6dyfl3d0XlyMLIKEvjvBzjZTmTEJyS2
LaNfTKDTzXkWPNbZZ7nEpb3G3oBFCVNqG2TLKowjUFlDBOIT4UhMazAo+JylKksMyroCkArpkNG4
0c9rmyFNhcwpBahKohsocum5QroJSgTxKbDNzBfZ5iNbvMWYsHn5ED74zkJeaGS4g2ITz3nBrnEK
vcTHAkw+/ULA9frqrEQNOpE1Di/QspoCbfKMa2x82/PwFDz0W/4L++2tMB1URBjXq/myZfsStzox
3yMKU39TUbt7Yd/+5L4yaShkoNcpdl6PT772qWRZRPkBE9OUiOW3qSae5OOv7X7Jv79vv3gNnv9P
g3kYOzPPUxWxCKDVU2xD2075i9zZll3moOTe0hgV1TI4EssMlKeUIRMdPQ1EbhpHK+YXRTQTCQun
A6J5VVEUnShM3XejB12AQZacw0WhguAXqlkqcWETiOUZKgVTJm8D1fkihKwxF4zfWi5mbEnd69J2
qsxgQZa96V11CA1C+8W4SAJ1py6rv/i7NMHV44qBu5X0ZXJYHu0FV9R7GvaVAvIl2qR4G7rGNFdZ
GgcWwBc5t73r3v2H5Ra+3H1lFfyHwMlEAFD5V/c0FxMbUKeJu4eT1i0ejMdjJDOTdb/mGnUVluTL
ZxG34qN6c00ap0+8+gJWdLUH1E3ifUo3ub8iR6BIm9TKpPSaIOg//knbmMTfuSgBEVq2ag2aRFzb
cQ3rFZx/k1NarFnNrRH/S3let1ZQHmdpo1pQT6QkX1lvz4WF8Uio+Y7YKH1gzFA3mFc4tIQ6/CP0
Is20Oc4oPZxO9+mHyFmB7VEfV2dqd4ljs90D6ACK3V7hcM1KONWshgel7SF6h43xpI21wnb7+nEt
YkuC7voJw5tUPtRwQLiZ2iNh0V/XgZeF+WnsaPg4F2pPFpc5fX1fA6ozw0RbIYmQOS+S0G8i+eV9
Up/KfkkEZpqwu7nxrPA/hdYuX6+uRw1XuQVjlSejvImb8RWdcbQvXLRxIGI0q6fiPa3cjTXiPGl0
TvedpApYsTGNzqhLQqnOpImd9lbOY7CgH5er3Cxamf5Fl1FRfjK51uXFB84CxfiCB+pxwiiGi/Ip
AwvFYp9AMGgM6txLXAjZJqE+NmQ7LPy0ZOrIs4pnQgIh+dSjdGlU7P/8WmmWc+xrroIOaKvpwOVy
OBe2Mr4sviKi4lwxcooU83D2ZxXfK7SBcaghLNKKKxshOvRe7o/p3LiTgIIVM7ahhoNo5l7ISKLV
b0CuDx48lHLZBr7EfQh10wJ0Ty/JDY2dLvEtAZqgtYy5wRIzusxbP6fYDz8CFOzTNUnn0mHtnjQB
gn+cfCfgNqDGwhz2QfliPEFGyUz3jFrIvK5pS83faT0xWJS6BbR928SjS+h4Q/waUSi9/vS669D7
jdv8PL4So/kXgMxl2/MyvNIR2/2fjJylrtxVE0Ltg1IH3TM8nj6ZEyKJT+KGVRrFW/8sE2pwN/ro
+ySirkFJdJm0OTP+zTX06w7ErgOydEnmTnT2NaC2vqj4rwmInGhfbpw/LcIC01mzFezLQuqBIZv2
ZXf2pwKGCCs5bTgD43WGeVLIKiRQwPjcPa6Kgu+vOeAhn2DFKevQk0sACkHhLq2bDBsya2yQEC+t
pMXKVprLvzvofoIkcFlHlRGmllm1r4iYhkQIq4W2lhfUWM0geNSxrTOlqreE1G1Q8iBNX/0aepKn
Yej8drjopGKYGdvmRsaH4S04krAQ8aXgPuvArNJ36BnwdTAAS92nVvIhBFVBx7t12QX9c2WBIasn
QHvSYhRwghqiM5cdH0ShtvFiLvi36SMarqosEHaNFPYskVmT5pYiBoNGyVIrmSKS1NqlNbrGlWGG
+Y/lrDHdUx7cM5ZR7wL8orovVnhwe7PpAZlaDOuqro2oIBCo5+JdjyWyA/tRpwgD0TNjxJ2uYYkn
pIMNYmGvRsL2wC0mBfumJXox44PrN5kOZAt2k+0bZx8FzbKc7PWq6PHL0gKqHFdhZiHrkmcjfbqp
8OYvdPGYUq0qCC2XCrgAaVAWAhxSoj+o//bAIlBasuqFw3os2p9P9F47n0EfadJaICCYn01la40y
sc4PrZMn25k5g/ThSAS9FWrQ6dzYZe4xeup4xbMelIVG5NdYuWkRLIUgHTatFVU/+QD2yuV0SnRv
G5YQK7Ls/RWRK+6sHD09jMuF+AqgSdtqIMJXEiy9eAlaxYGVZafRVg/QHDPK4HAzyCVZeIiV5c2I
evzKg0XM3nnPbI9f4yT+asNKC87s2RaSaE6jBQUg/j+eDXaV8MbxI4GQqY30iuG1Rp0NF0asD8SY
aHu1DVEDNFD37LnQW1lgZ7yFa3lsqkUnkecSZoJvfQ4btlq7YIGCsMO5JsQvhRFjlaBp+6bF0WCw
M3FiSBIsFkRY79kBzi8NuwuBFql6C3E2/63/B1o6UF8su8Q6GshF2y+i+ENg6iovn7U8iY0y1BJk
+/ECTqjSpU0DgjQpdK7KPqFlAaug/DaHZmU8qdIyYGpPn66yVApJcYlfdpIub8wVzcAuTn+h6LHW
ydIThs3AeWCeAOh6We1+NHxi6h+dyNe4cQdq+stuB4SrDJH4NU0mgrMf8Jfck81FOxsmWNbDQkHT
SrJpqKACoG4ewxaMXLb5iPOEnXDbFUCyD7as11WGcVeu/hGs9MWy4bOabOOvtWWjfsIs0s7/3DOq
7/BdWcQbJg7XCXx8tePgnqK3/j7yX6dT8VP+RrBAOg7uspPKz57LxXeNHCX6ZKecgz5l5Ai6JxVz
NlQKOD/67eH8ElG1xDCg0psDo1Yd2nG+osvU6HmtukVST2XrEEjYrnpg4a/XxGWUUwZjGgDNQoEL
8QmEE+ghcfM28TiL9oiVmUPMwBIj3S4B4KIA36/F1ekmea2MzJqIzHwQ5WXKJKbhav01snu368qK
qDLgkr2hbc3J9dxFfT19b/vLVu1ls6Is2Y++uWU7+wpNmcdkdtVre1Z54VNwIDZLYz60TJWmpgAx
mp5uysB1TG6Q7LddiHazb95C061YIDn3k0DdlHmxXPufBOMY/oxLMvQOvh7yAWrO5tFKvqgu/Waq
DWDG9ld1P4OLnMiw9OclMJH/0+WUxd5rYGuB8tXF7wvXbCis+zRDRQWQHNF2+QbIeCsoRYr3qYx5
kwRrnjRdNgfMi7ALKD1E0mg57kxmpLLFsP6MJi5yG9BBudkNLOivUi+e9i8O11h3ejjOsFn8/4U6
FfJQ1SLJebJRQWPJODRmvi6ODI3JjOESZEdYHm8zwPLzbbZpado6vl3zAVWzqRX6EI3IXxMuE3VY
GmOLJu5+bJPmUIh8+4gFZO7IXhE9FhwOAQ3Bo/bRBtnzVsvgDMMc2B3ejDu/r9tUL+FPotJJURnR
k2Mr3A8MwVeptUaZ5zeKM3ER9Dd+z2yBhLkuchPwhMKvnvmO24jS8HVFczcOF4OAITtgPI4vXUyU
1FLMm0scjujb/A8feP7rHzukqTH48ThTjI1u2yYSDCQJ33kmF+uA/ntbBaMW0bGVhz2ogkywCIuE
0LfAiPVPoyfWUJ4m7Du8rzyXfITdxQFF8NLPGM9xb/Ooz4GE8VZ5fKlpCbfd8K4qopbGtmsozap6
dyaRUEdz/3p8MDosUjErNExS9PsYV2knNpfzqwD6E/8BdK29aWts+Iqbi1p2eIro8xmLKEpwF770
3T5TRU/7fPXqQabsxBeH5yjGDbNxkb4cCGLNWKsfJm+brmMXBEA5pm7sLBC+IyADPnBGJRUaQX0I
GNCm1wP2E70D7V2xQUHPy0U3Gj6YJvCs71DiN17iDubejN36WQkYwN1E69bjD65MslCPKH0q+/DB
VaWAz3tnmOlGlmm+a4Mhwur5DBhmXtmuwxgK2uykh+vL6nEP1rFv0XNSKfXDuIYavT5S4FN3lX4l
xO6LWnh40njAWluyYIhPegxEwAifzjBGD/zlg+uRuDmNpA1Wg+ngDOOUuOliXywDbUo7g0D1EDVz
kTLOoxP/EOxmuo6Vxuh9947ZJfCcgsSrRtJbvFNSEqo1t7tMq2iQlgGV7q9j1/bkHBCYDxtlqsTK
eduAhgXZNAfHFSB7M8dnChitWcK3s7wRHI7IU1f66UsieDjrYqcaL9SbNXbFU2KrakzvqdLKeiJv
OghoPR9c/ZZa+jqOlFcNzSj312YPoGh4ArexvfjKzbQfzJNOtH1uVahoKp/0QK7u3zXSSyg1wYLB
fAIyGAH8knv72ocC8Gc0k0jmp2vgTGuxUSFnFvOXkZB7yKpXD2TUNPAeZ3gByuoeO0Tt5dZJpM2o
8gFnLHkvzA7UfucbQcR5rh7jegkzhfDIoXlF0JCnDsfYUfSecTK6Sfh84oX8Pj7bespGwSdPBlj+
+uFnUW+nqAMUHUdtOwSrgBnvzAwtdlEDFAdkiwuBjm0WAUdOTYv/L51041fQ3uIa1nzlGGVlUMwi
PAvDGD4lLVTw6jVLi7WaIWejnkkoBsdwhnxkNAfLgH5xdZPTgzc8sKTQvC4VRd2w21RDwYiP3nYK
l/FfsCOTP7SkE9xCcreDvCt76Ze6ZoQ4KXvqNN3Zc+20r5pEA9095byTsfHvaKQrKGan0ieoEzPZ
8hdcyHoYDtvASMfWgtFbAUll/gxaYwmL90h8MfoUmxDK/XG4k9fI0TKey3bkXY/VtOpkk1gISs9J
Gb9jQJXiFIN4fur/xOm72Y9LzFw7r15TPZ01EgapFlFSNMVWcAoNUXhTRRbQqJ8D9hM8vU5z5xkn
BS1xIEGVZ29yTihfVoFF4WNRAAgUOLlktprkU1MQ3ZGg3iFwG76T/ip8ZEF81HuhAo7ZEnQ8ZD6C
DTf7qkvCIcSbRSgcgcPtiQk4W4eFWhM5rt6WI5FJQZvv/YK5rufwELqa/Vl4pNeKmCqUlF8YRf8x
l+oeFMmJbHJ5A4YFj4quH5uC1Gajz8aaoX6u3bX+paxMMKA4AJOvKGRpG0SMeMK2gbNbjOf94A4j
YIMOczYw2qjeuK1+zL9jOK+vbO8K4M/f1VP6Gdg1LVzcKFB9T/z/AhjcKhdeKNnIwyIdB1/XGLhH
6AQJDIXAq5wSqj4anbcPeBjE29IKnuLi7Uj+wcs+OCOO4ULp9yqyl1v7M48RepI0pJ6Np1jYUfLy
8Pcbhzi5coIDWz1Vyl23oO+ox9oDywmt6B5W4v2U6kYhelwkOoXked6r+Nm9Inz7JvTaveCOBpUJ
8D7/P777oh/SvEvVv4yYABi6xzpo1DriGbM6/gyIfD50kNAc0HxyJkOZq8qRKbv4TsiADLyZhIW/
4+eXmPY9NfOaDMQTrw7BDYMT3gKbs29sPEtgwn1RT1IXlX7KdaTWZVPEqsGNvWp89k9E/il8us3p
bi72DF66FBxfoc7Df+uB+UcwGrKlxfc7fJ1CWGFt55HDzV1qC9wFlIjQU81Q0xmk6UfxW4DYo8s9
7nUppXIzuKfy6SFy4HIH4SidrlAj3MTvTHPNUEM/rnRkIGhgeXbrlM9hFv4mfM++p33J6wbfbtv1
3oDrYErrFujxr4pypAXa7CjLqYKc+Cx5hInn9a0Xfnu+cPcHCfGf76ZSgE2De7yzRP7Iww/8GkBz
IvcHBP1yGiuwWuATCq8GP5MNnWx1T+nPSrdU/2Ni7LfmT/lRBP7Bn6LjIuI9sSHskDj/oATtAzWx
emG0adJUyKzMnHu3ciLtrIg6pdODVfYbXyH8iuH1AB+J1+jZas2BJrqoGzhDnNovrCGlhYULctZi
NWnWMvm8xfnDrJeRt4CHXPHuCIUOoQbiO0wSV2dAAkJHUaEh4dVv/Eo5aSC1en7gliaLo2uTsrpJ
tbkiv03919u/5NXEyY2V+bjoOLn5TxoRNlnEzZYZknMmPJL8SVSOQjjazMXgY1SQuLXzAVdDt7Ot
E73cGO4zCU2lL8ZxOvclNpKIPEaf/AMeGTRZXf3u1JokNBDBfHdariKoUtiFPjz2FuDumqsas9UI
Aztek6Hb5/vC8OLdvtmH2GBSoVu7rxnuG3qUQuPt+hU3T58lt9TIDyaqKNNd5PnJwwyJFLiOt+Sd
/ykFnct140K4BHKc64JlKIjL90V8Rb+SmSiLF/QSjkf04tNISW74AQesbsKBnusfbgrqeZzKSOs0
EI8pmM1ot5feA8Jxy4maUjqRmIhK76ZVMaPr3u3oGYauSp8hg3Jt9UMdVaaT2eCb+nk5uHA8dtIA
51HWFsbuuakVKsJ4DhZ7zL9R6dC4qxqrwAWTATl1BF9tEV+h2KlpOBTbwWo4oDYpzi1NqdrdHPtk
l1QMJxotuQA8EYWzlAv4NQ6xOcT2TlfL4IF028Dr/m/d4YOecw5WCyW31NSdVkxcKp54tEUJcUin
SYEuwjXiZTaHh4q2Ptekbyq04/K7blvYz7RK8tZ7Ty2mjBZyndBy+kw4gViIBYTyrUOWzA+02nk5
yUY89C/Bh46JOLE31JIywwbaSfM8qXtY5IbAkfRVMbxnAChj1JrMKmoI5YLU4HTo0ABgaoNjDSM0
T7yIBWrbVwGXwwID/Kii1sFyfN4s0zaTbEbksOzOM76x+iXwpz+eeC1dEjggO54jG3wDyjrq1uuC
/Zjq40D+vKb5y+xSWj9JWn79PtS90W0t3w1ZwIHqHC50ZVdnUJyNaKmjatkWhvopPQp4nDL9XwJ4
QwQGpreFnxISZGxCJNtGtMSAxR8M7XAsJPEx0qoHi6iYsDoHpUt0DGnBBtHb5SYYnadbdm6+29Dl
2woCZRM7GLIM3t188aJ++BRAjSOuEX2ShZfiTKhUkQehYur2Mh7WI9WhVgNcikeYtPaamt85C6Ql
uvmcIkQyhw2qy89bNES9IN5V+0GwE1gkZd3chk7znf1+6GeOnUe5zhgDFUGGpJOEvqXAgv/cmTaT
abvTGBmQ546s1ZS7puQaeGpVHjdMoSv8TJ7lLSQQMTz01KTSWpPEGnypffnS61UW/+Hn5zR101pf
GRSZ4c09ndKPhHrw3NMS2iM0D0xht6cyjCu2UsoUCt91PxVbFPwB/DAA7HUudUbR01/22uJmiT5m
EGU229+NAlfvQ5LTXCnolS7nnoSoGOTmZeM0Goh/YXB02yHnUPxfYOnwBnV+gBR3G+nc+875RTe4
MYSUSCmzj2BCvPSsciZ6QNptErpIKugT5LdjB2bfvyKnpGXn860aaQ4UDebij/CJOUh90CUuwQvU
VBxaIpYk2hnRdzzFbXsgEOTlXOoiuqq/y3ZjxIbazkzt9kouaHt8z3aJYtCIsGVxIA49sasIZ5uV
AXZs/c40oP1I7gjB/ZSdtSFAvgE3XriTGFKrnnuTkOVR5KmQ9BR4zlztaekQz2CWRCqLAvEl13Tt
8TvUq390k7giBzopo7TE8uSA6ADiUGLhv0bzOXiks9QXecsfxZ29JjLn1znimJwhJLiMCiOTGY+2
p/jN4+QSkxB/oIS/cXHIvBKlIyUKqmssnL32e6MY02JddEu86lLcfWKD2PTr/wsFjvCbIYB4CfT9
EFVU5I29M9YPtd6xjgEXaQ1Y0MEYjMv0yO24hcXIRsmcDSsxzBcW902B8zU0kBtsV9Ny3RCReM9l
c8HFQAil3497eIUKpzr0icwoJTzgvguYaaRz9AwKl+75k6H+E0NmDYdHx8T0x70VxapgnzZcWtDZ
qt8DNg8lGEUhSfhp/+m2498YA9QyFxTp/PYA6ZVtxKrdIIbCDAMA/yDKwZHcxGnlFfe/b/mrwKjR
8c1lCDUwuk6O7tj+k+mMY1pL4UncO99TEGpGhEjmKt/ijlEo03t+e9funG+7EFMGLfmi8MKmKtSr
+dql6JDFiqGp+o340+N3qB0+ymlyL0Iag3MgzkIfVuoG0x36z029hmVaar/fvbdXSfmYTjx5LhC4
KSRTIkT4WW2GLWNLRBUQvhh09prh1QmMnni0Z5GWTs30QoCaOcu0jCZj9vDgXA6ciwFDo54rq/Zq
OClwPlYhOjYXwOhCuCZnUteL0PyeH19pUwTP/iElg9VLMrHMjRRLG7/uigjvDzWXkdezCYcFnyLl
/gFFg/avqeyOeyv6WfqkXg67q28CatvR6KKw0LwqIi9V8v6Y+DMCFl9ZV1rYm997gU0OfAXtTl2I
Ys1cWhlCkVvJ1Nh+e1ujAb08aHkgluopHbiwemsLQvxR2o1W38iKFhlRFP8R5ZoMPsVtqyJtl5RI
JGX4KzR5yuR5ZXyPKXDiXcq6b2JI7jp2dFEnFim0TL8hHg7PQXTBKr2i+IfIQ4lnao2D0niDHJhr
g6sJUqkm2mJmxr2zvIPPBkv107XJvsHxsuXmJxC6Tweky6SfMe9Lbu4AVfNdLzMdUcPXNpZup8JB
xysG2brzS4eCcFm94iLBMx31v5Aj1tdQBewVNe6oDTwIP2rAjYqAbq5bhzvQ2+ucB+giAAvzcbTQ
3enkqzgIfipeKibdU6ZR2iP3M5T4r3/h9H+hZ94jtxwcwA01zWuXmrfGO+41ZToEQGb4m8MWhQCS
x1xzQLXkRAKAvnDqjyYipqXoRXnbUaKlAXVEkqmGEG4fIbrHmzMCDWiMGUOGILvamXxGR1bMmnnW
Kfe+QxAqzZHotf7OYv0WS1dXVEG2rx5dPcN6YeESlbg+CfpPD3FBx2ytViRjFRsxEyb8Qa733cHy
0gZdR5k+Z5FThI2EK/gGC9sL5eNURuMI9s9Ps6l6SLxFJ9phEzBNMbxOHTmjmUrL3Vtx0k3pGZPC
TuOYh6teibZ7CjIc6ccPwlaOE4yK+N4O6YToB3A1jVw8JzcXyEnJkCNhy4O2C3jydLybff5T7Vj4
+VV9wgH74mblcfFPeeBve84NRyd2b6cNZ9bWsft5+ONbk3gD+RYG3dxCcPzGuzgT1xGooyrbz1c5
/p8TpVTmgH59U7xmRBQD8PfP/fyvFzypqva1yhXCcAGNUQwhPx70HWQMcM2mFI5E3LdUiMjSA7kK
C44IxbvpLOESUAQmtP0eGGnAEli/ta6sWhEahh1+VPu7j6IUboqCq0snCYWZpNty0wLBl33zPnW5
q1Us3zHx0bq3c6UhbKPyKGly1lLU4tfIRU0nsg018w5tmTapZn3gg76nzBpGoDWu/RDzaM44tDsv
mNsuvgHNuoWAgHH6LEq+v0uZEQKkWGy0ti9PTMFLtAhSWIvZg+GSNBXHcu1ooO7270ZR+vKlngGc
Ty8OMpDWYH5wE0xzGnnUz1FzU5ode/fs2j3EsX7KQQah1Rp7GDtansKqxUQXqe6EPErJbsO39NtH
yi1oFr+ewPJhikZzP29Dk9aGaPESWnOejGgVSymkG28T9vu5Sjnr5GcWqDftbIpXmbUDFyFWN9kC
DekLVoaDU2hh9pexSEXXiE2Tb7AGByzeykNXEqWaLPjtLmfCNCvA4SaXocKeN2PUNL1ZoWuEMXV8
lrP2+0//ZXVtCpfykh90orLyCciWGsxOVXFeb+fZH0nyr9ry3u09kzuWivEDegwIuHTiACbxxH+6
d0in8ImSe0GhooOdNhbkuapge4wjlquwjXIQNZrAQRAZtg2A1SpOoRH2FEF5x2NlQxDzNpvnPsHq
SBEdsnF5CZwzpSOn9wk1yd7fHu7AqWOGaoaoiioIIvn3ZDyEGFN0fsMygOeh7g1dQ4mNaNJ/2XRK
gKLbUMJaJ2xl8ZZlgAks7n7c+5M5xK7S4aJuvoi9+GYAj2gnqGy0UnCdrtb69lyGPKUtoKTzxobY
vPzSPc3H66aa4N5+TXq+viyB/osB2CxjiZ4CRy3+AvGwXPTl9CqovIVQsMKGKWg3hC+iPqGMNfyy
+icCokwxyKjNqsxj3NJIzhaypaU2YFvSK+6Pd3ooQzsrgB2pjlvBpBDzhiHi56reocmSDQRFCaBy
3gH+qfpstFb9MBypbGwhxAz9Adsil/uaa6OStx/nqjyMzm4eVni+CD13R7DXDcpbk0npfEGCnf6a
Az4EcMUG4KyIq7zxGHH+J8E3RxfdIE46iJwFgiDm5+edZRDXmvr2dxF0eA803Wu/GuanPinku1HW
vFnivmd/NNTq2uw5eODM0JtNbYK/jXtUr60OM6LrC9815mCgmepoo9MhXp6K6DTiBfB1b/Qldkci
ZrDLbpGaJZA6Hb54UHpDnBOrGBeXp0O501Figv0IP3DUfgnIpOO77XUM3t7Vfub/vs14KRsWGnw8
RzaLbPdkjwQSafH0XKP7KpcbVdvYQB0zQUWctsart5d5RtymWvi4p726I+zZK4ye2MhVXIvLVafA
ysmusllROjHQzrTzSymvHD15jZOHm/nkape7Lo53crG+FguI0WjjlDxVHCGZB4xv8CoE3e+3CD4q
Cu7urCe8yG7sVc8n3b/4xNeJKlhQT0tCX4HgfmipcR6tgWX3EC+nWY1ElMaTqb4UKtVvkyE1ggur
zPk9yjIikZ4/r22hm1dpsjuMExZPz2uSlBug8SvTnfgRofHjbUlXzML82WQA53RJ0+Trb3ZRHkJ5
rRBIWHLYs/THtHnXjFQPkiU0W3Zd8aQaGGWmRKdsEwX7pe+nrPYO7/gP5FyrOIdFdx0i0A1rVeJc
m3xFkAtwSTafEkOsEnVtW6iUsYBgIj3r9MxxqmB8zg312Oi8jcWkYfLzYoQ+DPp8+qL9/Esv0Tw6
sG1C2lvVmO6/CfohfCdseWizwXFePaU/B87pIg5N7SHgUDR8qO6NGK8mIq0Zt35+pV4QbM65wNmH
+fckWQaWAQPI22JKUXF2mpIg6PVjc0n29IBjX0CrHaatV9ydNpZdhaSkksrrMXRxk+K9DEJWQaAl
p1RVS+jpb2xhE/QzFETt7xyQE5RV9HWZ878q7DtjHyaRehbG0l0nMu5/5AX1gY40Kd9zNrbhB8P4
RKgs1OKoWcbUtLCNnS5gnZw6viVD5PPnvPqXKOfUAXeGS6IGpu60Yl0x92mDvxavz0CufOpXIbiZ
VBN+6wznMnuvwdUj+o+Bt0t3CQia1Vv//BtI/FyHjNofjkPSowqVjK3UJgSPpsUOnOOx8RxNYN4h
t35XxGQE2gLcpsKN2YqdJuMjXx+7oN8WElCT9nRNB5jgwnMnF4IJ5x0zIZEIhLNYaGXWMRDpc+lS
TTJQLnJd0NmnKZX/ERy3vGwIbiiuWx8DTv7BPTcnGLl1K7DPAqu/TEi7qLfnujlUKwbwy4TVpE6C
9Sc8XcOWYDE4k1vtRoBdxbacylL9I2wxzuLb+rNwPOWiDPIUo6n0RBMDMcjLO2Oi2uR/3wK+j37D
9EyVlfJa+kWLWD37oG0jvrt/zTiByPqAmKOX/rcYw0IaZvlN1xlT97yuHN6kScf5EjDBGarY5bkk
RKBwrPPWpg5lxB1RLTgN8+xwEOvsHX+637WsvlIWfG4FSiv91Z8vLitJpMt83tcKtvScefB189Ly
In7Dn3+Qkhm55etjic4/iInHjBTSJTPCkIoNk/H/YfcrKXZKXWTAsaxmJLC50L835lWr5MKzW7+r
OXjmfqZCOGhJ+BbimsVrxI/LUPXsJqLZcPaBmbH8uCal3YsiyPvB68qGIBcTD7sLYmKLKRcgchNT
6Wk8yuj6uVobSh5NZqpj150b0p7VzaB7gpTezfnk5/UX58LV0rmqIAkaWBB9RCqs3J1JUmrzii3p
q45HfhQyEXXxS+za2drhh+5mgoBnACXxEZ4WhJqmJ1wDJoKWLMLJVpmkeh3S9xSgUlg6oXAu/6Jt
K56b6F/11KaEwvK7/JGbEPhSVYKYixeIxAJ4yp++gW+qdUB2t/2/sJ9Be6NoNlqT20FXrOoHDgQp
w9p2AaulNPpu0GRDh8EfNE4We23cG+nqcEcOw9giBgciXkd/u+JO5mnleUM1tQxsQNf79c3zoOFN
woihBgaBPp1gcJZJnDdRt/lRtjtJYKyt+8zRnM16dURtWRdC237VjHwQ43Ei5mnGBgOhiwLv954U
6NzcJDB5kXCJkO00c5TWxWURae5hpqxVf7n095hmpzK6rPpNNkm4rJRxRA9psjP6FqPz6zuw3C7z
U9qD2hhoW5+fWdO5fg42b948gEODiYmK1ijG285B5kZ8nbUbEa/sRGz11kFpd19+FNddUON9OZH0
ERbuUrm02dMGl/cWdxYO9sSe1eCDdC6R2sJ2OW02bBA6VNxT98WHUe/HWJIYwuGV2pdJbM7DQToL
owJsBMHnahTFFtEvb8JG0SzWbNcOhNPvfikJIMSwzv8JF2KAxo9GOnp+SPhVTt86zVEEXIjWjLwg
33KnMF6XSuBTMe8vOU+QkAlR3oFf7t8maUhQOPEZlQFoETebZWvMdmlEBBzbu4ZsDBnziYWP+RSR
fmftoZyvaqQ1PMAzGs7vE12tLdQJc29XMAvApbrCSREEb6B75EcoOxSzYz/EMdCZUIhbO441+Ijw
Q0lE5cU8rJE1on0JdDSsMYgNNa/YZLN5wp3B/Rk7AOMXgosVnl+pTkZldMqNnNLk/F0O6GIS7Jwz
oYVsf9WbEWQHgIvdocH/mmhWYD+GyR8SDey60xfsK26DUejWR5yK6irG0VR2KvCiVnp+Jnf8MMuW
MPD1DWpe4vy86yfCc1d8hhjVkfrX8AsJ7uxzTEYGZX7OesEwCVBu7LNtWg1wze089S6uLdNyxf6v
/bFHs97prSSzn+2fNQN+FOtM5G2Pdng21jvLdtr6Ho8A9LT/p2L0MAnpdTW18Fy3pYEj+9wLiJyF
B2EwiA9l2X3RuiZGQYiMrf0m4aPnVhTo+dZXXNy272akERhjO/S8KWmF9YOLuW87vr2HeKoDC+tr
dhsfM1gUPMB1b7iBXnZQcbJvDIEY31grJOevbQImOXstwO6XGGR1q1kvDjNHIz+aWxnDfmdiIbZE
fb7WUgljL7JibSUdF4zstd/TW7XUXNcJiQlg60VBmrIC+E8VLeyYp/tblmA9gSpGnZrfQdff0HS2
nLuRP09ChZM6veLPCiBecPIj5pdlrWpwpmkLwsnxHVGnE6+jhoqnkJDz9GW1c7yV6r/yRrXV3OMf
XHcR7r4Na2bpunfYVpk7QHXSnse0v5f3suuHSmc2giMLQKSP0r8T+oXwnqWEuKg+NjubV59Dwf+0
NhQb1iBaiqgkkTOGluKUOnqo6TRrl6zqlv4Lj02AemlFciykcis3eURuI8inWP5mowUK2/lj+nPB
jcVj8CAwOJaDsMNM3AzQTZTCWSVKn3AES1RH37yhK8Et3SUB1DoGZHllApcZOCAcCrGtVhs3tJoB
zci31tweZPkYZvuB/yzDtJRxlZDR5lfzRKWZKqrafEPg6Wk78x4AlY30l1v6uk1AcsbzEFhmGkei
zhCVC+OAnj2xdikX5iWeeJoteBkginqyBdPlkwNVYKRqOdWAGX7BgTtySnWuNgLAHtCmoQYmPZmd
yBfblFYI6VlDZAVgy7agewawXbMKGsmhm1pKpFmNLqKJDEHKQEXh6ViHcBRjweznukQGFFKAtVfS
QVujJmxA3w9quXo4n6I5GJfMKAgSVuZ1O0fIbzYrwWkpY12Gt/PmRhYJssevWDWDyFg6AiwU0NPY
Ylx66XoaaJLHyTQPyMRmvLxJPzxHOfF5+IaBFPTw64cErY8LCXzWM+z2YCaLfvihfc1VVrxwPNu9
EEljCj+fJ0JovpVFR7MUFZV2Bw97vsGtuwIWwmeBfbAp7g9giTikA1Oaz+zgqWS1mbaj0CnK/+mj
SBrP2DO/LLIzXu7SS3v7a5kO6yPvAUpe0Sx1Mx7Ji8GvVU/1QV/0463cNJur16XCZQgzSM82mLK9
lJMgWhgaRj79kJaAX5TX/FohlZRX55sU7KAMnR7/OmPd0UpAgo/UHFFD5013BO85b0RYi3sOC6xR
unBy5a64KDVaOBoIFGHINnJ9++i4BoG9IMnu4PWS4yqDtBzbyYLaEImsMyjgMNZ0V/anHXIOzGso
xnI9A8AlBs5kiKa1Kx3C385epmldes8nfh1f6DbRonWO3rU7IQPODSLY7vZAeSiSI++t6vcircdg
+gz2Arq2BEziOOfOUfZUBjuly+fw2OvWxkzGyr9aa8xR5sATpyPjevvtCdR9dvIxaaNyCS9IfzjL
xDaOUF0vzfw62AwMgFQv/1M7I3o3a/rTQMpDLT7UO3RECBD8UCI7/VNQpjR6aJxlS+a1IEbKstP1
gdnk3IOSEEQHEmFGYywX4o3m+BMVy/sEY4STYrCnmoiBBjeZMSwYdG1Msdz6s7hdj+eXjpCDEGLT
UKQi4xyjwJyH7/JF2QcML+X4GdSS4h4+TdDkFjV15E2R5FfJbUlOCruTRHAMu+JcbBYDSdM/Y48T
5zxpdosOHiPCtSQl8WOFfwfczVVdNvrgEa7Krtgvv3HqBZHtaRzwRfSM/6g94+geK2zrDF9fmjyX
wngqicVbR9QZQV20KoDkVke22zdjpk984u65+ovMBswrAXnfJ6RU921jGl2g0P1L30msVrmNBAQr
jEMtFxYa/gH5dbJxK6hR1DbDNTHGXZ6t7CmzsTV4GVGq4F8udsv54pC3ywEhyFMyex78FhUz93tn
5s+3x8tNiCSeIsQnR4qZlKqEvm8shJ1GDfRONn8ZodEENRJESN/CcyonC2FIO1fThoDxoF+2LUp+
5xkh/V/gwIQLij5Yp81m5MkoPolZbmN/mAlsCAu2kTzy3MOVqWpxV5fMhh69R8dmrRPOdZl4UZd+
OS3d2XN382NdsFwAK5KKudQsKlI2ZfuE+ov4IgbjLTFUQo9q4UT3sC8CfxwX3xjfCYo0rCrT1m4x
KUD0vUgWBWzSMxfqYsdLqfiYlkpkwYk9xRo03fSUSACXxTKg9P70TCBNqaodyHiAwEPNhpzortn3
J6P61SfIUXdXv+Ced1ba2daofeWUsZIW9Awu1z3OAmp5z2IAtEhvIfDy8/p+phJH0SR+YyEB2IE2
lgqXaJwI0r0xtCXK8Dgo36CzXK/KPzZx2Gcd5nThJ5KTvTaY6KH/cxFw67buzjJmNS2uEWFT7fac
OM/YcDfA6Pykq99R++hFCFUZ2CS5oWn4yWOj0sbftMzfXRCkWKJkDa7b0wgmOlXPlHJIqF0YbfsY
5Jch8znVkkgcLfcPM+XNf+DKSdXCloyfkQJjZhCTfDcxxx4T2SBTeKsy5hywkHWOBPhQvl4RhpO9
ZZYe0lLImZDhoFvsKuv+Y49ZN9V9bNgPRjWgkIsVbgijL9hLwc3aj/AUt2mY8nMti0e40FCoNIRG
8zvzJq2DO9n5imhXxcw0Fanaa4gdeCaa/BCiLguGvASAKJ82pnThGSw4gLTqltqcITmjM6of5NGB
5R4epzivrKwYSw1/zUuZv5tEjSY2MujNuIF8hPKayx0GUAD5w6KYP46BWzsI+ZPSQdptZz3PS33R
5jxjjaqaAh2xtNH9y1pjjKKid6CAcXm5WGhSBhF4jlWlNVZDNeuk6TKeWptS0HXh9h+WSAcvyzLE
42vbsS5062wCPsWLLnOdT0tJqnD4UvP8aC4pvmKqrtWwy4NDgKRlZ3M5FMA2ooAJkcwtsUJkfr57
Q1gvgUGS7XC1iVy/t9Xyfr4C7fp2nRBNqQkO4Czmm98VjrabLgHIJUvrFgiP2kv5BHvS01vgSkK2
U91YmhCqiXCXgwUVBxqBDl7iLn2eBK/W44VuhHKywfEZHhrJIfXghiEos/83zu1fYspkgfgAd7Qq
Iixb7wKOb7quTJeQxhkGIj6UpLmciYsZ6KmAq21vp2AQ907D2V/R6L5St5XWO85jNXHrA7QMX1OF
jwQvAiBx0c/xqlHqGX/VX7IL/dvW9ezJYyhTtd3IRm9uUR4PnDukJrIVPPkDDfFp/SuGmlQ8GPGZ
GbwQLDGTfTuTvVsgLd+wa0/GI7wN29Mdw9hQQjkSwVT+ySRukCiajTc4cd/wr46WpnlDUVte6aE2
fMR8GTC8EwhuXRFNpOEL7Cw+JdUPhqrWCCWN8JNY9Coy8QiojgCXCgpnIeygTqHWWLjDnjVwSvSE
q1GErBg35KqGB047bDWASH6W0c61lTBS3DsPq4kUMSseSmwBleKk3nRYuxsonx5q0n5W7uxfvJ9s
DFylzUkvuOi4utHWs2FB7YE46D9a0pkRmy5B4o6M425dHAjSrPkG+pRjGYIRTFaLTF05Rha2NINj
pgujblHWw5z7KmFDvgzkiUiWIYgPxjsCTCHZkEGgiswbVqnWSaseFux04zLMgM4yHW9PSPUphM0E
mtdDEtlRu8TnUaESWmtXkA133ZxdSYArnF3+BxWAywqK227p6xgUeoE8xXRAIw8Wn12NOhlV7jwe
JOGGlcrA9pl4kR3UaEfDmoAwBWClm2FK5pxo1xVOnahUzWc4m1/tTyyDUvjFWBi77RvrTnW7XeSq
7A8OBOIamp14xHOyhFVuopywo9hGICll6l6sKFA97l4LpYjbbQublqcMY89NqbX8W8dDh8WGK/6P
40wWyK+9XSCCIFiF8LpVqj3M4Xi4hKN7vnj6kLYOtdT2c/4TTO0MZ5YbwzqEGpE6KArt5gxu6Gmx
be+OBLXsGe/fxrkrvnHYUGHJGNfT4bya7Q67kz7hgJTnj0ZtdHjGCnNt7XP8f/aLz5jwaTqQdLS6
QgGXz8H3j8ieENSR9un2SInOst7QjP/F+a08maU72dEXgTXQfBvvFK64QPExUR3thJKQfbWoVBWq
est8NfInlNVw82mLSm2LCrh5y5lHkxj8kaO7cvOMtjr107O7P8IufhuGhZHfpTUY12WpZdOtv6SL
zFQUdZ5sTifAMxJE5NBvd3/mUIaArXyC1doRuqHge8nG5UVrBqqc/GVj733pSurlsMFz87v9DPw/
CnyQuALJI6ygHKeNXjkjx5HBgu99h1rYYDzOVeMGlN1LlHcGO5oWF+PCuY37Hf90RugGDw2clfAB
cnGeS9dM70sJ64a+WQBJdBz+mzVVUzMBAhas3AHlS9h0n5mCRMl+pN07hox1eN4H5fBkXTqnczkI
0EO+Zjc0b/++Y08Uhf89sLKTb0YuXDwD569xWXCKealFbK8k1Bd2eILzBSczBTW5daVAp0OIe7f8
vxz6yZJErvmEguM/vQArMLHH3FLdGffrasS2ahAi7vAIGIKur34ldCCAs5XAzXi5s+PB892EF5HM
jPvf63PszcNoIufqaPvf98GsDrtVZ7/4/mRWvyH7O8Id4pFmR0xvWO80EwA5wSp/+KLg/7HMZO18
o3+++eLoxUhKjK5ikfUIwdYZ9Y25dSG98TY6tJ8rKCegO48NghF33lzh0sf4D7zwTMSQrhuVDxgW
uKsZqB8dBjDXMRB5GWT4wpExWBRgj5y3Rp6kOpeMoDzIJXtI673pVSwBnLMrbRZV/XGrnb/Z1Jze
U3/4+F3XVxgySkjTBo64fB/FUFzKlk/d/euObxcw64vmI0V7KI1/kZ9K/vZFKpiCpbq7rXyqhhMT
ZpHBBlVsba9MDtH8wb3XtxsrnZkuPHP7BA+AWyQU2p3nSr/CNJJXF4n/AhikEjDzN9O25slie2of
h9oY+FkRzQ2h2o5uZ7UXL8HL/Hd64Rm/I33ph0fr34syGjBioZcGu4BPHNZi2J+WlggSRrfraUcm
R/6X+7vzYepym6g5nU2S6LMMcqAMMVwRnVuUwGZOf8pThNQjNS6h1aqah5c5RlDqPw4e7yakBk7z
6SkajEjA+hxhA1opAOETN+Iso3D7OTIIyV67MarPFZC3m121s+whMIYw+NQend/kGlTt8iJh7SYb
8qtE/V/Fr3kqji3dz6oGg5a3dI1Kqcebs6B8ezZMcypxr+I3+9Vakp+h/wRe43Wxv+Wzvh5rZQqW
QzQAoC/ZebHXJxdVBHZ3Ex7g8zJQkm2JMaS3vUZOr/shN8dc6XojqRbkY0cGF98DA9IX5GFF6PLa
3BtCxwmyYKuWOKHYLOf/T2CP+TSCa8xuPbGXsymp6J1/GlMbadctMeSW8OeGcxRV4J0tMcgFeMQJ
KE1HnFvIEUC1n+th/5QPhOpq80wWU+gLRlP9c5byXgbUFJFjC3H/OM0FnVwobkJKR3mI3JMeRCel
AchSKuygB4jGdsMeF9RKm50LJMjCCGfZW5OR79dPhrunGnM059MNIZRSMQspyRp6btuGvYpGdSB+
l7DZLrZEc0uHcwE+6odoBQdP30Y4vlWAUsKEefkneIDFS6A1QU3SsU8qXh+bOLvreXzPLXBTCoEG
vGcCfAKJdh/VFQPqG1AVplS1l4MlLuLFOgFUizpMWWukq7CxLXFm6Gr1C1xhV87nlZmcvfqgPt2K
vtQhm85ef294wfY5Kgedbns8oGXbMdVRsDkgJ0vVFjGaono8kJJlklT5Ae6hQKOP/HOSWQf39J/l
BqntGx5G5w42+sVNJwQo00xBW2sKNlKx/hRGhL4PRYo0WOZTY/nnJMKbDVWDphR7GIqe6Mh+b2vc
oQIRa4uDn2clWHqlAlO91Akqku3/OUcxGjsLgaj6kdqOchsBKAyrVUoZiXOrEDyDwVFfnC1JvHWh
aNG06E0g059Wd8qWwAk6BseLo0I/ItSVDPH4FC2TUKux1R/8an3p3udou+qAUnQuema1J9B1mkSg
+ld3yA8OF3mGk0Lj50rkJG7FOMeutxy5kaC6G6QW2YYXgARbumaGILrJSxlp7izXSETZ6+4+vX0U
zfZZkHMw23TSsGbB2LkIGD9+ytzXCfsMsmafAw8eNIkCbxePlbvBtrSwGVAE5laMNcJw2tqBhPbP
OqGNL3/ha9myzyE6B5+Mu+Dp7dQoe+EIFeDmTVnKFOhTkY2MMwYzTxwOe9U/jbIg9MMEdf/9H0kK
Q6nc+PJs8wMojix1sj0gkHEN/gSSOWxybcXr2k0YYgILFE8VejLjdDTRg/XfRqkCsM1VMEKHu/mm
BKcgyseuJMH+Szt9zMjJFFmEqVytdXfo/7STOdYxHyfqQeHqP+6n213fWdfR0J2pfnHDURrMIj1L
10Akmm3gxn8bnJpNAmrKZqZa8TIrtJx17vIp4J9NuF16fXmZFrNodMPNeBKCMDVUHRhTLJVz+eBQ
QVtXhkcelRGVgjEmsGOw/tfD8QT9qn0s9cfsYlbJk3OzbgVaqJkPiwJPGICY8RpUduTQGbfBHZ8H
DDVMjD/vYNZrXEjrEzO7zYxrZ2HthEsz9Oq/k50tdhukvT4mJGzyS1fsmPWA03XUraQIx37OWVW0
Vpudf7Cdp5PUtU6kCswJ6B5OgZFW/W+vwuyKCkyKPumhaG5zx9XEpgdmsXrpapEOkQNgViZYeGP9
hqk0924Y7DU5TInub21GGgVy8HyWwYrtjklHOcHxis2Dsr5e2k8ysIa8MF+fcsCITLANfAtpfAAB
nKHXXm/amW2vmr6ybn/OtgQ5YW1W8LQMa4C+PDIj5DI2pHLyHNNyZQ6RZUOZG5xHjF9IFQGocse5
l6p4A8e80Euiqi40Go/sMsjN+Trt0wAFaA9YpVkCfI8SR2kRSKpHc7VqdlNyCEoZzA7ZYfM/lIvI
SVgIad7Z/qWP21372VPluQEOViZlQkV7fzEf/sbxNglWsbzqGS7g8d39KYKoCmyBZuEhhXphciJG
nrZnNqVwA+7IoMPW+bPoPV/umZZBCY9iQKD0h8tSrVjIEfMcAcuZ//LZ39+BLvG1e9mhyjcvPClW
24hNSqt9ACqRoR5j8GK0/o3q3ED9sdELt/CpH/URiQcwf9BBRR0SRMfguXIT8heOnzButhbqv8x9
8JhbPWxe3ajI7a1xbhKOjXBr4M9vydxwz1VwP1sp1bvIiJwFieF1OxO01iQ5TkLslivxfbN4LAau
2biJre4p1aepy2jSiUP2kh11/2djFsOEtY59ziig5dSvjCYaqRSEdvc3fCtDeckTU3qF/qFhRYEu
YKjQu1u7pSem1V9iyK84yxbJi5xz8XYsbQfa/ZD/bSz/cNOnxrrSVPY6Vr3A1brtgd/Wy9vPGOtK
9VtwhDjaK3ZXyE2gnTitg1B9d+UGI/y2ETXxhG1L8xeHtmBzeycJGQqWcy9t21HY/AmUqvaPtCYI
AG9jm5Vzgl8RQPVjDwgKf73j4CnRalw7H14L9V/Sy4oARY4YHosBTOhJOKvaH9EN9lFuWpC1RrXy
kylVfq7r81tu1IZHNpUsZFPdlMojLbqm9J/WoiT8UTA9GmhJbnkSVbCEyVldnj08aIzpZPqQyvIi
tWZvtGBH6m0wXJLWEcdkt5hTZxuPp9kjEvrP6mEqRa97rbOcAQLtJ6sgS0uTSLlb9eecdt+aigF7
DA/d2PCbbocDzu9kxaQDoQrCOOaXwECLkAIqkyPA8WN3WxgZqihi1cWxZYSGAANArXXeKXnGdKt4
6gWJV8U31nbO1gWr8+coj7lxOkylp/ucVPBs8UElLPTvojFOCVKQ773NuWyGpijAsbMBIYQPejJm
0RMEB3IR/Y0BOID7hgfEVfdXQnd0xjfNUUG38ZmmnQR7O/vNDGzJlXwcPlHeOqfuDtPKdo6m5Yw0
oCSnqGROS59d4UIMp4NNhQXeAO+/Ptyc5kWz9iyAdHvwidxLEpHMteWBSPkFlB561DX5V9u2FKXu
XYoT3zF/nJRNpS66uBIPl4fnVBg/XLJ3ETERgjObEc6v/EGej3g0KEIzTfclcSzhtVaNxmbKbDGM
j1tW7txLKm4F+LBKfGsLQouhPGa1IMFWiLjc/rB2qFD4mFT6fWSNgGIscxxpu1/QAaZ5CqxKZvBH
Z7Bfb0CFBJ+IsCP5njozzuSivaHBC/DB5qOQOaWBqbVmfMyTPsdL/7u7L2Ciwwo9SEgetMYe60Ei
eta4yqW+WY0dWBmmF8PWbHrXJO8RtqaGTCAGgDlzqSG7oB9CnT+QVNXTOzDeZyjgLNEVvLNGnE5w
JH/CkzwG73haWQHEYXlZ+8gZ+9IxnLyyDAPQMiom2uaifX1yCbNItiNirNiDPZPaLDVfyHK/uyxA
wZXxjb3kcCrgEpSyIHUcQoQxECkkHduiuvl3Pie6Pe8c0G3vYTGD8PnLFVdyh+1cY1YjoEbM4UTU
kbNS8ln1WSC9E3xqezfpwkAgcgjgDcIKLZMfvXSj1dJ3zL+Ju0WjYzbZdT0XceIbkbAcuFYA7EmO
JKm80AUzgtSNpJM2dz5hXNwTIHiwetsP/A6kQ8cG78s2JO2shNg6mLGjPUwzOlzC31MO3tPQ5v0j
8GcEuxMFD4hnQ7yz5zUG4oExUC6EnKu4wYMPWdj5qMyjfR2+qwR+05Gr0slPyN2nmBvPC232yFkw
zx53onWNnYmmpob3V/mOzyjK7a8+YliX4M3Q5J/G53XK5YJVgvwiRjjIEeWTIb8Wm2SmHsjFt6Yy
IPQHyl/2qQ/Cu/xBqj4I8ttkOyy9BeHUbHBzWqf8hNzAhXVhYUq3OnpPJ1yyizreMbeOwmkNEV2Y
pVGU6HCrXvokzneLuIjpySk8+MfXw2HxLcts+NpF/Jfpt9XZUOF3vFcm6J7DD7fu8CcElSQFYrIH
/PlywXJg7+/JIhlemIQ8anVo846UgwTYmqshO7Kcfro4KAQ+n+d7J9a5GLvMASiS2/wOTx6XaIGe
1LopiXDvAflLq8e9AXUwWkbs7ik/s8p19RDrjkoW46Im6fbj4ow1317+nlYIvWX2jfIWg+EAHj7z
8ENykplPlhbG4D/EhyVpbEcH/kmB+6Qjx7/PMjwq+ai9thS+Zx++nnH7wQrshog1PzGAhqmzFUGZ
ff5RsBIHeeIQLKSVW3cgSZlFeIresg6kZKKslNrDgLQ6nioStp3xQgyoUbgl695xGupbbuLkMgDs
oxoe6CmzBKpFPGAr3s5ikRy9YObAnaOtxYCIrYcENSSC5FxOQBmqanuxnNhYWkOZ+1yaum1tyzsA
0oUO9xHbSV7udXCUw6/FySkLgl1d56xWFr8l2kpobLJa5KJPVsBNE+DKv1xdh2kvrCMQo6AJsN6i
WRAYptNVse/iM2YFam58w/Wk+k3gKC0m1tMI8VUnPkg5arjBFLKR/SMvo+NKbUDEalL9nHr6IkdW
jsovBKC8W/G7c49zeENsLFc0TODCG4Je9lHuLT8ePsyk6PsWqUMGzHA0iogKotZBgDRVkwjRfeX7
kLOGLScI3ovpAWWKZQIf36nApryITrhqyu3Oi16TKsTZG9cj+Ln1uevYuyXgUq2dZW1lCn3N6JU6
Ma5o06OrX8bUjScA/+eZh5goRLKWrKXIH2SApFnn4/1X1vyAcHxVpe6dPvgfVBf9XKXVL/QA7eMU
JPA9rNEXHcgw3puIm4JpKusJT1zOJ5Gr2jhVxwKIA0QYL5LuTBxGCNNJPss+f8FMFUTKAbrfHhyo
ovjElP4DPy/ONqtqLE2Kt37e0iWCy/7FOhVU9DKzRO+qbVrnU8M2gEfEkGvESK+yUkp1xlSz6cFH
1ZHsKClbGrH2Vy2eOMpNnSKjTt6YqYiV4i7OYHESYdnbTgjcMAJLy26sMaSzghAA6h9udpnEmz76
hO9+WPHEjyHK4n/JeBWEfnBizYn8K4K5/eMXoYVb3JXv+zhbbUk5eJwbSypE/VdsRu2IBq0UEZt4
OlpoJU7VItZxHjOIyTBMk5wv3tIrPSR4IMmSIfHAtb2GVlYzJCXZca2N7ZI4GaoV6DLK2AkrAcDK
4IRDUVEbs0BjKK40/tQ5fUoCpImDfLMAQxAxXjqZbGz5eIcYUwOVygq0V2x7/2qFD+EHsP78cRin
PAa5MTTOQx2UNKNuvLOVaQBn9xd4pBiVtStbZIxKMokzWzSiCrgjdCj7z5+C1qslpHr9fMHAKc5r
p8Vaink+evFlLieYLguBxOCufyQwek0fYDiZLsRrJcZ9xNI4cPYuHnJ8f6+hYX2hXGh/czYI4Rp9
u1tdh6g6u7NWJ/K6eAyVt/fxKbB7PXEpiZH28iMMtLbX0HssMxPaYGJ1YS9EMktkETNM56hQBluC
NKv89LU8JLD5107dh2zWqtPxTIdkAA8gWLym1i7X/JCksTzTXUExoP4jjVb5YgQt8FlPIjOqCUrr
mqEjlGOx0l0Ihkz//WLA8OT/cTMFBlWMdLN9x7jIaq38EgNMw6vGJ3fdPRoTUTh4oqoHntB9KaOy
CrDCm0Z394sk+k475wuEU4wrVuLrgESTRROUVhf1G0zykTNVh634ocWn5gvl5Ed5q8Ibyd4z3jK1
fIhBPmyV2RCchyAU0b5Md1v15aqgg479SpUOZ5TCvdhitkFuWJL5CnXV2ctpzU+M8OqK3CdWyACv
N8SOh1cfRoiSYoP0un0onOCrzESGlbZpRi4ejSu5gVP3GEAdZO8Bmz28w3/JY18wUzQfycdBmwJv
IJQXXPm9e2/f8/rID15iu8tKTgPZKZ8BlrlAk/toJqGOQ11pNj2Wg17lXhrMn8cj6UJe39Oe5gJh
SBSKLqpVG5HWGfNIUUGVN0lqdQIlGIyN7SV2FLbaUaDo8hEIxIXugLsh4ruK3b/GBmYWXK5OU1NI
3AAwCltK4fRV2sb4dwg1V3Fxa5L3v4agY4NafQS7GIhcijPC2qvZItf/l779S12mx0D3X6Z2F3Ur
uisiVjse7jv/blQmEnWv6zm7PxK3HP7JcFQCRCcyuivZKb0FZucVvsv4Izuq+wXJrs/VsUMfsnaA
TLeuVdvuotkLcNc3e5ppwIm41tu1SR/Na50AFFI8DcVAw/gf4P5bI7GLOjpCFYJWyTgj86oIq/P7
tcrOF8UTc10dAjeXZUm4HX1rKPmvbLsPege+cg41F/j0OuOZOOPi4XnbSXx7j/ayxUofD/H2h2yd
uv40pU2eV/BbYMMoc+59UxdHkoKwW7T1SdTBdEdebT4EF97dP3L1Q1cGUMA8xzmx6R0XKnz7cgTH
V2Qrbi1YsvP/1WMC6oBjERnC6gNMwkonkdBx4W0wSrPjz9Q+lb1cvLUIvrCk1v3zPNGPSrf6N6p7
Tt22XBxOMQqmwvrQso0+8jGf5HUmptsPQRJLrhUjt6rxkcg8N77Yq2ke09yuq17mStW6+tqpJ5VE
07va15M9SzHU/uu7UmV193tSdY9+9HzyMsELMn1hPlADi6Qz+oSi53jhp8CT7EbiN0K3LYCbdTFl
/Up+XyY3lue+rk6N/aZhThIQxhkUoMIbNyHTMVeyDC0xbI1BPA1pW3DKH6xPHJX2JBR9MoIpRUjn
71qHlKjP9TGlhR+t/241fwHiTnyU93g5sjTglSrvlRo/Dpy4b3eka2q+2AWriC4SRxPGr502/RxS
TzWteG6XZzCNXB6SepsVh3xtmP0qWkbJsrp1FtfjlLqKzOs5XSc1IilN6TDwwneHni+jVCQJk2gZ
eNKrfzWs9s31QEY+ZrvhYZ9Hbu6MHdQW5CVCXM4Ids+FP11VHjfkzyV4hltE7LzSAvMymbDKrc0Z
iRuvcKOetQCAhBQ6+rT73gzQZmElvUCR2xzvzUXvQEVNLnw+2hgvDISA/0fM8sMRyhNyc6QDHO+S
E/P8rJi7bxMs9/jzM902e77bq5S4jlGqk23FZ94YT6ODbII21jLUWhj9BPEQYEijNAyWCYebLdyB
GyyJHTe1WKnCC1J7E8SuO7W3qIsDPWg/YHVTs1g9u2oCtJtDJi/715vO31JkAAQj3+JLE9clrNMQ
+IILmCOuuAiusmdrC+wS+OqsLPYq41VJcYKNYCbe0V4/6sIQfA1Z6zSeS3luFGy3KdU1s+2tLEIT
tfZBOm0A7EpmtV/YAFocf1hvMVNcoE14qZcVQ4dFkbwuCEeF5NI4KMw1MRUhKUPQ98OgF5qvhw6b
YavV18fbmsrxZkWBOYVYpQ3bbaACTF4u0TJzUWzwSF0Hbbh5fZI0P9sMZeAXm5cjCMwMP1s2lhAu
iH+LyXPoremb1DfodsXFWwPd770goJgBHelgNIrTWgCpAHjj+5zs4AAuXRnXVoRGTXacDxtCg2B/
yM+FuvAYRffmKk82kXlgvSRRTlUrk7Tm+pH8W3C+hj5YZ1fd+GzlTKOMQVGFdWKZV76qeg6yDKQM
ZXd9knjrGht+/xu0FtV5AgUaIrYzaayj8Shqx7mh8y+gbxSdOWrxBPuUd0qWu5zqmkZjuk5sFedQ
0N0OTkPZpe7BXSdAqbIUrz5VxnR+FoMBPLKPwsx/RSK7VlI3QxptT05cmKsvd6wrW6SQB84h31aN
ivqttCobEu5sqlG8mfJgGi86oM/oKQ2y0vX2VBQsrvm/IIHY9O/9hnQKpLerP5fZXU0mknw3PgJA
/21mDYwJJc3S8vECVjmh4+JFYDYMHcSI5x2xXZpS7nYpahFFrtLntSbEaMyB1pMqPggDLciPp3HR
BObtas5WCcpxpqZRqOE/OI8FRzWasiXX7YYOsQJsgQJO2RzWcKHSWW93XE9W2DGWZxelL6cw+F0L
lGC6JCQSeVQtOJ/RZ6WRyvxc3vHaQAr5eZEEvPOb1YIRn7W7HqJLL8Tglv/2PKmVeXj7jCtI0p4e
qmtT4TzLLO4Ed8eWtrLmm4zZemCXMR6rOI1xETGdFrr8rUuYT90Ae2L3LKVG6syvxjPd/njJjl3+
n4skbJ6bOZD+fwbnU1JCfJE3lVtkNvNpUU41g7H5NegzWLghGuL22PW48A+t+zu1elfDzMvKpazK
SS1i4RLCu4YJawEq80JjGHUk5zGWZGVbQOo7iRH1AZoMB6JWwR7KX88wTaU8tQbGypxGPbvjNPVg
zxL54Ba2pUJrGfxzYybJnq5RLl4msJTLjUjHvi79B8WIWg4Yr38gY+h6aH+6b47P/QpnqOOHZ3X9
EMnV02vRf8kTbx5eUJj1IYIZ95KzW99/9ond5nu6Glj7p95hhG1To7dBjxjGRIBXs3VZDKU9KA+T
50BSbsiTCnBK/UOoGBwdz1dAs+P1Yg6QWYiygJyn6z15hStYGHS/S6hrqaEAA56l57YC20zASRMQ
J3Q59qAJTBqup4nWra+i4esrl5BJWBJ+kjAneTkFoNblcFg8z2TJw0E8Xrp7B7PkQoBVMmV+5MIg
i5x5BFnibatryHDT+XH9f2yaTU2vR0hv6ZqCq7sU8AgY5auAPhca73S29Cyu3UksSDadJXcHlUiA
IZACFGQmoxXP0GzE/iTHQYN7kN/VvEAK3fmCc1xBkSc85qS2SGyGGdOGAfc+nUphGbL47pd/7y1n
SlWlMXGs92A3i5nQwAyYl6aRWafZz4wzfLbvOd6sPj5v8goWoa1zxnt1OE2DaWYxSFJ8p8WLLdKV
Sxmcqt2HwlfISdlByMCjxvjXheujhY/HODVtIeaattFBoa4oKWI0DxTTLZsw8EL5Yw8vieFao9ni
WyF5e9Xad+1BW/iLo8WgslZTVY2IsI2CnG0YAOJy0gtvbpDHQb7FktIdYjz2UYP/2QPYi+wII+HG
gAoy5vJD6AYSxWaPz7SCr42faCJDlzXX2fO3hE/0nZ1bz8Lym4P0LAac8DBS3tozsl3gauD2NEfr
MiHRpsquEXQalIPbEDlBZ1m+Qt+Q+82AGt/+L/9IEm7JYYGeBz23VvrdeKK0+gY7UWIWBF3N6P5D
PAiCGdnwyspxq4P/1lqZuLJyStuWnS366qkzbr9pzZ0YZpES4sw0MQjD8JTGalDqsarcRQ8mliXj
3Jw5PReBKQj87aKm9Tguih6gw+IxEvaJqTwkQtWzhpwJLgP5cR7EPnlSjsqmagyX9LRXIwOemtpc
qWSYwZo50yWqA7kyE+8oL8h9LI+FhgwWjD5MhitNjGdnNe3ftLFSwbbZPM9qZ+IP79KZLTqNSZ+g
hhJaI5vfqcJyHn4qnS/ChMvOPheztDjx7OBDT8719OVK6TGetf7wvhqbym0Ffzb3Edvq/oOoPqQL
JOlvh8ashARD57DI1tEtT25OkLLxrRPAso0HCyJ8zR561jJln4T6YO/q+aWkg+44Z5kkqx8btq1K
bMEg1v536P6PK2s2Yd3FIxmwuB9h11NquTQ+Eho58EREGebSzh4UamkW6E/h7bNWYYHM/mZPasZz
8NZvPXhF18M8HkopcV+62OZoh7J4mxAJNN/HOnOG2fMUcChBoJOj2TqrEccSf1z4xgaWxTKTLCep
ezV2c9LWkHPFuDiW775HemHERKWx8dnndUrVVlZqd8DOdvYOYsX/JhshgEpIxhLzx1A2V8LTWILA
CrwnY2n2u5h77Upf9yxPsJpywha4VXYTblzFebathj5W45x81vQNQBCtYrBnqZk8KhtevTgssNru
4rDdmNjZMxWDTxwKKAGRrLtkLn4oGHGlynxcnl25hTy8GZmn3Su9EG+odEpVf3RAFadUAUnCk8h2
/YMeYIUzpWTrmuQd1OG+vEqyx/DhUef9RneEP5Bmyb0gsbm4V1ErnJUovTp9zzT7Wn4zfSrEImRR
4qRzxIIqD/fleb19JGleLMsG/POit0HYhz0QrHjK8Wv1uUQYCKOPeTUszPGcu9ItwUA/0+XNNDGj
FcjU9/iMpL9ejlQjIN/d6fyqaaI1AG8G59TCBD31zgkfidbi0eX1aOPt4JnLJ5mxPzUMMzrQ+aw8
Mrnue3DSiGr+Mrli6kRDiPMrsamwBzoDT9fLR0YQ/WoqnRz8sf9cJbAoqrGAlYcY/dbdNWrbj65w
RrXkj4AW9ik+BfaeGirSJYbj5leXoDKxVtiEUDFvOca/kSMDvXRIvDMmfBrBxHR2Q9ekrBBHE5RU
guU3+aKVyuCUNnXBhbzHULu82x7LSeY5l0oxGcwCkADL0zc7yg/KQ4GTwxaKXSwrLgKNxmJRpJYC
yGdtJ5wlojqzL4zWX/J2qjlBSclfIFW1m3j797e7JOxM5HPCd2hmJDT3W716gATnhgWXD6ez6XAq
f9+TI4ybYaZnZJBMJ1m/QstRTmZp8Sxeio9MWzZMfGw/pQwrOpEYNQHVjimFyOpNvAfZHi9G3b5L
fmhp/MAgvXm/7u6dGDxTCKplvF1XFgdMGGtU6XqrazDD1p/hP62CCu7eaITwR1dyf8dnB0+yInlu
eYNHpqY1oIKe309kSgI/AGsIWAnIOiNDVknoyyz7Ol4srsOOD6tBUPzvQTGV45NP743dHOVpad6D
+qnJ+ZNe2VfKynFYsqPbHvidnxMvS8yruxmRGvj+bXMTCMOIRnINgC8ubMDe1Hd9OckJ2iS8Dq1O
8h6sYpZUNaTd5uFzXRBRTEYBxZGamLGtD9kv5tY7aofErZEXnNPkatiYTe2F0Wl4I53v3V9Dr89N
+jZEaVz5zC4E/vUdHfzMyNqajcopY20OA5fmakgbGD0PvaTdXKFitPMx2hhSl3/kklrPtHComJQB
U7Oaqd3OuldELug6xAPdujakITzkESQGERYC2MgAYEGY8xcr2CtCUbcFnRQzNC8wKNFb373UVCaI
UVkAwHk4pBNkL+ZM7B/7s5pcKGcEzb5TpSzMRY21Y2zugY+qPSSZc9HsSvOXm45TmoUL/hxT4UAM
GcvV0ul3tIc9DJ5jLuXB2v7g6LbQaAY6sUpoCoz/f5AF6n7xb5Tc4B1hOnvf6mTFb4dPqnysSyAi
GJy3CsEdY/g2AzKn4oFdvBn+dVJ+tDUjmIxWloSBX27V4MiBi1l/EGTplY2wjshQHxPRxC9nFYwN
sGpdLkjOjvqah7PpFx3amaySBejufs8QMLzE8F+PrxVE7c3ZF8W4o6jbxtLdxM6dDe6KoPKBZsxj
vag8W7c630IRA+UcJfpbb6WXHLzsntMuY4T9A4q66M80GtdpgVkCJL0V+9Qfgpbq+Z62nVkkIw23
hmB19jxsG3nvpYtuUDHOKfxXt+aSxYPkWs9NW1VZtTWwtX+U7/hbT5YdCpX80B/ZKXfSqV8DDi6h
NSItE0yBrc9pKXTA/z734e3QEQPlIQAgrW7BYrrbKX/7YGAVpzO/yjknowARtcAv3N5PhvWDzoL1
EXbe9kZOrqqQ7cg+uZH2XyIuqb42SiQ5i9aHXozfqqHiTM6Y08OJV3Llt3Em/RuU+djpQPiQf+rx
T+l54hZZQ0sQvzLNa1jEXqnzH5O4ep/IGO2zJ5/uKVDA6wldU/vwEDT+UWqwlvt5Yy/rKTk9KUts
ff4Wv0NHOzRUTG2aTh2W8cMVo82WTx/q/wYbAEiv66kUv1YbOcYLBDjk4Z9IZQE6jWOXeNiNKR+2
FhrkXfRPGJrV9099gzSVSycZ0udegexR2NwyCce4Alfra1vy6wLBBeVFdx8oBc3Y+FBLf1q+hPkK
wTjxDHho0yrbZOC0IKjZx5dP/d8o2XMmFZCO94lIxDoAjkmy4TiAW3ujRP+9QxZcdorykP6h+fgp
XwDYI+sJn697dRhxzsoDynXU29FJ3FlSetmCy7QzEbS1Qx2W/ZNBY+5S2Rp2zlbn7q2cV3lCvdBP
5Xn/9qx7+X7o3w8519U/BqK5P8cBJwd8UrVzmHxB4cgdxgOAOEC2lUOXm7zrWzQyz1uauxM9oLza
KuVQl3yUBWrRf04SW5iXiJvuPYU9g/5zsqdBNitYR/sYZz9CuMgybfNY4254wlSyK2mzXqaMgJOL
7TRigtB1ZbJC+7NfjgEnIEYODjaKOnTbj7v9Cub7F6S4vSAg7DOjbSQz0JxdZUKNQjGZGcJr+y42
cOXETR9l6RYhWuM+I4FQflxmnC598Sbx9YZ22aiHKK1HN1PlIMjk8L7QmCEDhWsrYLbL2fy/eSIH
S7CQIramV/QZmTs6ZXAQUsBz2JSW55gool5EbF30VRtAPyXLpa7yS/efCdltTxdTvZDlUHsx5gXc
rZ373h3SWETW4AR+CItffOaOKh3l6xy/em4tgOVsLmxUlxMlN6ShM4OFGny++RLDNwiJSETrI6B/
x32wq8CoDy75npJAUyUIQR4LXr3Rk/aHbGUIrWmFmNFzScs+YK9iYqYdbt8rCWPMq5dlrxXSjaWb
iRfs+vRIIu3bOsn8fi811DGG9ZUOxjJn8G/3rD/z+oy9WyQDoBbrqWGCLgE+NuFxGnN9u44pOoEQ
9GouVqo2WP2VOtoJRlpXeon3hH2MhMPL9hX8OAu12cU7loYN8ZMe624BWijKdOAAxSGXn917x2N3
/5gzSleU5c+HwKoZaKepFzBV56cD7lOO+eWCZSA9ML7vWMCQamea1xhSr01NVkg0BiN2w5fJJ8ov
O8aWkbzZFzq5v6fYM4FmBcJRcgiMW7eQ1HpcDt9hsZg+KzWhHeCOutQmTIbvy3MnJw+ZkDkg4NJ7
saP3ZEMo5rFwyStEyTiOzjVuD2j7SIZdkrk/t7sfaTneJrNUhbwEEEs8deOivlq6iDTFXF//73d6
KXvEuG3po9IKBQqbh3C0rgPKnitoX1XTonZ0+9i5p/tmQIx1aMvRzUExLg1II756d2MxvWbbhPFQ
pXIHD+udFF20GlUIDyCcLyPT1OXGuS56IllwpYyvgCPxTP/udhwG9HM+RnxIlDahjpNW0klzv4MU
uhPO+51NoUNHZyWbx0sX6HLCt4Sj/llQ0FMQBQ3wIPJyzF+tvnDe8smo0hGC59foeEpAmrDoMJo5
s4V5F+qZ3SkLF2o2R4fyfc95v9hmCMc2BA10xI0F54K02fIQ7ajBKTYND/IFH7hKwTDUEQW4W5rV
XFw40D1PZYWhBxqyxZ23ndlp+dcuNGFHuz/7MyLkpv0urmY33aJKzpWdgL51QdA1quGdoC5gS5eH
7LPIam4ww3jBBvE4s4dyTulaiOH5YcylvrrAuZOBXhnp24PhnWyTHOvjP/vD+EGzbEHzVthD8bZU
a3lcofsvH8mdpx6dJxW+pYDrVC3iHsou9bpUmWGPuofQ2Xxihl+CMAWqbHjvBQqMa92ALGsvEror
vWZe90w5UiERmYkd29a3BxvRy4MC0cTNoyNDpUb/H9OMTF5nPzaGvQonDDboxjDHwdrbNmdyurfx
01hN3qmIKkdh6v0k+yoZbJ2B5+mDtdk7YmSShimE2abYrdBy4PcIL7I2i58aGWp/suXCWSvQAS+x
sG1PNM/W2GbiUWKlnZVk0FSvRSl3wtlNOWvJvrXmcRaacv3PV53Rz+qTJDHbmLoIoc5azo9QkA7v
jAp90YXtv6bAUUV38lH1kPwes60bC11IELsdAme9h3GdSSEl4LKjv6oyuZCRXdWq1L2/CxG6Hd6E
xus8VkrdYUYTApAsiLcG18fLiasBdhZ5hTE1f+eC1C3UcJ79YBhUY7y9wQIWxX2jfVsO1vkQ01VF
nUFu/qsYOLwEseOOZ7IcZ0ePgkPNBzmhR8xJl0sPPlVp/y7pBZNLLAeEBm370sdSDZCruXFN2fiW
Nl328+8QZt5FAnd8yaS5ncU6kLQ6JVw2BHpwelJbqhzBibpP/GNn9jZt/dWlCpUowU2G4VhP8363
eBIvzMD8hcv9pDfb8/aq8YL/3FbbaWE1K281yRaDxcyQmVF4pG9L5pXCGlOcz/LVrbKFLsKVqmst
ZPEASXcSVfGHiVvPSr9VwJsV1vOOTJe/7Y7IzjwqpyuaelH5PXZ4IeHsdD5fh4caHtv3yHY37NqR
7MS+egf7lAZXjdaKJkQBZ6hHahSsjTAZCXjKUeQURw/vTpVkovCysLYO4SmPHYX7sCrRkwfjobd1
gQgbzm5zpzmz+uepGCGomNzrCDVjPK7x0DNQT3RTymC0jBUJwIbWqbbEx4wbI5iQT1H3ZbXSUTNt
YyEZrunOSyXq5yvRjyD3FUU+N9xLI5vY8jNUq038aNpwQnRvGdXiTvMTpxZ8wRXZYwiE8X5eJQuR
ZmrYN8hZIR1smYV9EUg077HPe/shiy47KjP6bsQeBuw4FMcVGplYyfpyy/Y3+eBjOENaSRWVefut
MIHN96JBdhJGownJRCt0ZY3b3FwIIYU+F4LkNMgXzLD6LgADIUx33gR/RnDsnedo1fYmCczZmYNy
nnaM4kVknVI3b8TYTm4dweUzM6JPp8gtKnlfbYFt1bbUhFDOLSlg7S8/uj3ishZMfl12UCADMZNm
PA1pNYl/3+rsYQyVzJK8cfVsVPfbvYBQMQu38d2bHZwKcD1EW7LS/22qXl1B6dz7dLO5NVPONKNq
z4JFNtzbS4XgaZNXotiayJiroPGIl+ZHNsxhqet3aH/2INy2YaKhpdN0So7Mfd2Dj/ALi8dbnbV6
ppvkZfc+w2cWrD+pnobvQYoqJLuT16wAzEobVkEC9T2w+ZoCPBuxeFbRoZGLsLS83VirAee2KZUw
k93SrQUrNgpeRyDMzs2+hoFBWIHzfncxoBZjyReLZVpu1RMEnQxkAd/yD/fZcDfsrQXR25Zl97BU
IkHnKRVX7HRlo+TH8bv1egENMFCoD43/FrB2boh6B1LY45tARkehrN267gDpEOOQeoKwXJKB+Jzq
phuaER0QpLCTBKBNe9I+gX2SLYKegAQnESRhV9Dk2ti0IK676bMA6zKc+V+L1bKBWoM2yfOXW1Zr
1mp1HWdlLNvfButMNQVh/KnX9DDzHORmL5zbtf54NVT0X1mAvQxUbF/IyNLYNxoslGOr7yE2q7PQ
8EBjg9m7weN+K2UAm0F5TRdxxnfu2BjJDMoHhIoAyjI6lqy1uu4yR2t8sIfVIZCV69bG+niF5U+k
1ChqBSRlg2NOMwllODdLNUjVh/NKTFjGnGp+fnoD49S6SnLjWyaWjSO1WPnv5OXFZpSjKXQknIYX
VaLpzbqH1e+wMoaLaXIX57GgpxT8eTUVaVbBs4HtnKfVihtscSwsaudOOVNe/Yz7rp6vLz1cSi8I
kDbuViexpNGyN3PpaPtc2oyrkLFIa0xt25Kc7r9bni4/LmfYrui+j+F0XraxgvNpNX5DUO+ANhmr
eSqpdUVgl4qN+/d7jkD3EGjD8SVbeRM6LFvWZd9xLsS+LmyNT75peYV7LWNo/MyMVPZIJKgsDIO5
lUUZGwzN927mItzAHPpeJM2MNYPGmvj6MTB67CW/84dAuMyU2hfb/8QYQedGoOha6RSr+Do7prJx
dqQmwQBY535dR+uhry2iJHLnU87i893MnT7ikJHdqeAot5PSaovrrg1S2naK7LbGVK2XvxvDoDVy
995mDbwr8IZ/rCkViN58U+0+o1Lke803csjPPeL6Bxjk3kwhK5XCOR+1rK49b/fPTsTtNBhjQ/Yi
k3WGNxgVpZPYNe+l6YDogAzl3olYg9XuuSCSL93VB0zqVuENGgePIMZ7SaAsgk2qCqKjVuDVJooA
5ef1z9vnq15nOiEZbo342eCpFOqT/28vXLO+mJh0UBV2R6Fs1AeJZX+5oHK/OAY6Lz9DTkwr7uo1
oGfOzrVUCMqgzNsERfxM1YRhX2Q/t0ZiCOCszFye6Dixq7qu6tqaDM12S/FjI3munI0+fK4bpAW0
SFa5fOMsGzFw5vhsiUSjKW4RtiW1C+8vabO2FGdC1+IHquGiiJGAV3YoORB3SaT3FC6BAvxc0upf
VqmOigAp1PzTmysgMz4uQBh+AOOaZTxh+YVviPJEUTKdoeyAVs2HgNuIOBqEAtSw8bNVPs4z/nGM
tdHKJ1WGZaeOcsY6af12LmFwfUllQKjVoP5achsEXRd12ZSle2rcg3nxLD+jLiklSTQYGmAljyWm
46l7+1XmX7317BOzxVGEb5hxgvGRAWddO8QGLJf6rTup2Hco/EWuT35FITpHAq4tRBh1E/ocsCYk
kQv/OGoWDkB7v0TRCwzNLNUSfAMpBgBlhMGTugFhxQ3eVlS95b9RXdKaMwQjBun01fTgM6HAdzn8
vPEHgvSC+SBnkVjlNO4dAUSQhA52Y3t8JV9m1Ul+Tq8B7eNBXjoqt1m0p5Zc1EmOr/But6zDyeiL
WEFPaaiH9JejEa0CgkFYkGRweJMthRrGjLfmBjacFvPzGo9nuHN9BdLDZuFZDPWRbWDrLY84Bwah
Ys3jLdgGtUfHjoonBGxS+3nFblfrWP3VxgIEwok+augCgFVFlc9fpfa2rljEFHaKt4GLejPegTZ+
bS8Cw/l+nOeps+NC9aa0Sib+/ZzQEOBlsoJYmPRpQMoVcB9qzAVoDjsUGbd0Wp3AT4t9bbCtHB6M
0TYpEiZGtHjqM4fNaI4Sx5SvM0UWrAJLkNnIKOGDowwf3sWaI+GMSMwG0bQLnVUur0aD8p8+5KMm
WlYEQduwVc17oKuFcoRx+ITB+se0+Ig+ZRxy035KNTOxi15T07BWws8bJ37MdZTz+jNvx8XixwUO
chajw6iQdeBVpbz/dE9s8SVHdd7+R+oUTgrm1z2zGwaTKc5lcmSxfsiJa+v10VJRhoza8D5IVzcW
oLzQYU0zSbvw9HC1fmZ16P17+yEuayQB90jY0+adj7B1G3ScEK3Pz7Xd/G26c9PTU9eU3mwTTL2R
diu4YHlmjCUJ79dTB/d25uaqD9VUz9ngbWjbFN0RrwQwbwLmtU7b/lz7TMtP9QssTwT5zLS9LXlP
QIC87hXXBtyWqwbncOfvgTIbd93FSN3BU+qZ/p7PDu/HXmdCDZHgskodK9iS8cGCXiz8EybJZc64
0NbZeHEokkFxiiG1g7W3zL1cVLHEB4Al04J13r2T54Sbyzv7mypuoIaehMogNYugbQIDWZ7m5Fmd
D7ehWmU0fiHL96A4mrQgTpw7LrpoQnHZ2omTdfRa/RYUbocuXeWErM878Usej6j5CO/BzI/QGPjB
KSE2Jr63Fqm3O2npChyhMRK0NdzCiMVUqhsPhrJ4B6bNmOXa8AtSDkqicKavVXKMj7Vo/aUx6Jce
cG3dnSWxo+vpTmMVzA6Q3MhYWcibCtoGlflHyYNdIS8r7onixUuXYp9/Nxtizs0pWxSZ8phXrN4d
OamQM5RNwRcB0gujTT4T9WL6iy2n+zlvYJwtEu+ELpmQVs6SJjpPrzbyoHNBiCXTh7a3PzXwrx3x
XLFvipxW2EpAoxYUUgpYbiHzwy7mFMDbHheXXD5Xk5DhiTDe+UeqQi5Jb3D8zJC/l6XMa4jO4ksG
4+52QRnKJJDIQY9PhiyWadn+q/+5xJ7kg7HD262JpLOCSwAC/cKvnBTe2yyd3qtrLnJoxA+PhprB
nnRyZBHaqWXHWeBCDzfEI67CIWGNG4kmYPgjiOZVaeDsFWGF9lUhsWjbsivyu8AdXghNkk5wJpsB
AbkSBX3gPp1mekduT7llEPzk9Mx8IHyQ0G5gU/y2h1YNbPq3DJOMWr2Ivdy8UC/K5JgyhXlf8HxY
MSgYeMBc2ahm29mBPMkVbiWYrYr5ayrQjs+jT7jLFYt1XUv3efjqWKnjx9hBFkBa/jDM+6lxQaLa
hogLd1XyG978ovekpL+N/p56NtNdlvzesn65Jrwzi4h2vh5mL7lV/mReVGp8tjI1ShrBfglaAb75
VJMwl1B1J/1mqmBJVScS8wDxhirqVdIMQAEeV1a+V1N2TjAGhlkhuWE/HK57Oxy3Y683Hd9zCvVf
Wu1i2yIgYmBNAcN4qjVmB2EhbgOqJ2vn2gazuwB/Hb7KK+QoDrlMnMGWk8VJi4y06rigNJjgS9Jg
/fGckeZBAsCtd87/9AVhlmbiT2HITXKrCjUOjmXDAjxMcOoELRzinjL2Bh5LF/lGXhK8M/6s+yRI
1AF4R8Im0RYjJ2WfA0ptC439yZtoLaHW/9WaTe4SJgoxz0mBxS36TDcRigeX+my4XfQSSZnS+/1p
/7Gilz0sqmHyLXvty3rm+3RhPo1eWsb66hZrtAcIjAXMhP4z/CSAvah52F7xQ8SONDC3kDmrCPmD
eu5eDgkJjH0c+c1Mwzhe1rn2idm06BG1zKNM794KjIschHNXM63YTjbm4h453+xnMZ+jpKhtP4xO
/EUJSd+/lFkI006kC4GPRpE8eaFI+CRx50rTYDnqVIqKher6dOvL7cv4iNC0k50zt64iHnX4tGXX
4Qh4TEX8H1f/t0AhB/pBDuBHLM6CkFEp5XEZHDcNI1epfemRGZbx8UuBuaDH5dlS6EZzv80SPdNk
2UIke7/vNwOH3gl8mqGj/e1Q6mwbYSVU4VqHa8YwnnMOcUMgy+K0KQzxAx8EX8OgP0UY9YJR/v+y
YVkm1M+AyeJbx6lKbwsU9cfa9EJ0XE+BJytsQ4EbMnMRQYrSYgK1gJqdTG3U7Lezmoa0RRF2W6Ug
a96jr5+1ytPDFYNQxavSN1+Pisa3ousBK9fhpUkYBT2AELnBKuaQ4TTCppLEAWJojX7TvGEbcndZ
4izkaS0vokyaPN8fKrachfeWxOpKCrOSGDl9gAL2BNVyQAKtzn10PqjDsUWVV2bqqWYDXcadfsFD
zDu2zX3FLfPRdpMlOgsJJYGnBX9Yw1FG9Us6SfDhTSz/1ATw3ctWNwR3SnF1WAY723gHLYwlmC1+
QU+ov+akP5mu+cG78FvTrlansEN7L6aGmSyJ5pE4I/HS4rQ3c3dbkndRZHr6iVV/fZDVPAWz9JGG
3+uz34EAvYroQITH61eMdbOJn8dggHqXo+q8yop6Tppw0ngol7pH5H01+0h31a9u03OeAJB6Kndb
bZtiOENk2L7D7rVzzvrt5xFeL6YJdZunABpxCsS2OAKkp7unimEo8xYTy5p+XFYZ3DfwxY2WF4V6
bgtLp6tLs4qxnrSgE7+/+2g8v2hlPeT/RbSZNpzHdpzvn8ol7PsZDqbxcgQFBythZHniYYXyaQoC
Uh9kacF44zm08pBcbjJ96AwDdIrbqbyiLOZ9PO/mO8jQM7EpvMhkBfCRrs8QioVEQqstUaecDH8P
kzOlJoHXA12S1V82LVhqN/BwDEMxO8Dz77w7Y2F/VMo8EOJaC/63Ainq5oGOfORMZUXgwJ6zgu1J
CUrbgH4NMmUqA7JcS9pPCaG4ojZMhlEUP26HX9jGgFRlvtSaD9xoXQEnHhxlamGVc5/nE8jHq8WS
Tn8Cd8TattjSYXTQC08ysEry5kWNHQRuHot2YMbynXyWqF52enxqH7KpRpaEZ75Gm3wtrDtCmv5O
R0c8QVhjNi7xlFG01hga66TKStaSW0ckJT83mmSSJ5Ao8zeKNoj4JBZU2vijG0bk/zkT3Zc87Dn3
SA0VdetjhuYXoimEXjMmdu+Y9RJu+pARnPebLUJOA5woSYEGn9vqzgOLhvxlO6uuYe/qkxz5R8cm
tP/iFMK8Qsd3U5fIZT6YvRiaaKudzWGdtBM9ymyWVwBtb+Zo3KSaeCCiEdBVw+0MMPsd97ob8flL
aooSStWK/N9vPhX14y2Y8rB/Y3/kbiqGSrcbmsiKDdk2VajLjgZlTMUw/zVj6LKlrlzxKB5TID0h
HzPWrwoUh58+P6IGE3Vg9fCy41kFmmmvn8fPC2ZPSeUYvgJzW1i9rLhHcRAN7SIJfmwgXTLAzqOr
/8Eho/H2JnrmslprfUQsarQoFZhhQv6A7Y6RHoe/iReDF6KLoDhFQAPByucvaFQKkF2pbnKanjY1
lOXoC8EClKlVZyHWHxdhOL0eqZBBY88ISs4Rt+MXWuzIHYkPwdbLzQrXqo9bdTkzMr85zEF3JlVp
14EBb4X0f6NC9hpEB057WiYy8JKWbuWgT+qLG88E0rjFTfvCZ1tP/Jk1JWvcljxRjdTVM0Qlr1fd
geVqRjpaTks2SY0IuNSCw8+2UyjSnWfWl8cADESViy537qoZ7ih9VuPm6VikkZ36tL4t+s1xGCNZ
sdvG/Q8rhmaLi9YfysLlob9XrcXpq2u2+qkYb/l8NPYs2deb3g5BZULuRPE5pndS93dMs8wX/o/r
kLl/pIOl6dRn9Uuvi3pLK//fxTNT3xXmnBUVOMn8KxVWEZeEX+mzmGx5GTgR+2ZQrOIuXqqTPqYh
QPKE2JVCHHdQ3MYUSzbjOPeen8JcDldeLSc+m9O49/M0Y/K73AC5JjjWwQWC/y9eqDHBFV7yhjEH
pqZMzkUm5TRBzPv32DhgJOBzjG75dTONkv9WtTv9Zyr1pGCSRgjSegu/rFjbi/y9Y7nCxR5wW6NV
DywmldrnQpP+0DlOSBndyj0Z4lCs9G3geZY5IpJDaARp/gfcNaU+Rbmpq2cOstG/8CZRwznbAPEY
BEn5JvFW6rN/pnsnj77ang1DJePiPsCHIvxrBxUANADkub0w/asINm81XMx2kMzvtEXCGXci4arN
6faB5eIM9niSivJIJyaJHNxX7B5y8iIBqumTLRrV3GfB4UMadClWHMsRJxfvz+wvq8AdRKnzaWtL
Np52qzhG/ICeYs7+zIkMIf1+BNH88gyuRjAgCSFw1DXSuWsICXnnb8N6vMnCce9wExnB8ljMIBh0
Yi2tEr6NYBQqyFHJkDFckmfBYvVOSlsk1BZ8xABBlfpvrDf7diHio7Npb6ZWQoljDyRr+BXYnppi
4Ln1sKXCfbcbaoYs+D4cJgYhmr+5aaWZVk7Z9Gfr4MXUhQXg6SCgNqgm924lrI5LhR4YKAkYSu8N
AEFGA2f1x7dHNLTAH3kIR3bs/ERHHe0HvuO1XYndraf/zvC/yjxXJ8olaoRNUC2nW9eX9cdjdn+g
OkysWitmw1RNM+aVyoxO1lnBlwRgbrMajlVSnjdib6JhR3uhtOKVCo4PbGJVGDdVS7z+tFTXY4fT
199la5Qalnsxb6fD1CVZO4Fy9CrzIC7nIeqMe8pNXLzrqILC3yNjqr0RvmlB+sQ74xSmrKUZCMvb
CaO88QMHHcAxWS/F4ZewQ/kSLKCtuo75kHdelNm5vDSemRSpc+Dfzww+CzM5g7fNmu2H43Y33f2M
OHDhsXfBnmrEwq+8s8OM43lqzXKlZe1DI80DceJMSejDvRHwuEoCrNtQNRQ1O7X/tuQ6503IdTbX
xWYv+2ObIxTpsK9dVcKEi9AOG04XEqyGhNPR0NMrIWYUqA6RKu978P+WT47CxXO23Sdl4jQtxvLK
Hz7ExZrCE5qKSK+LeYNpQuvEhCun4/AMR7xQCk2IaWX+PXQQ0Z1Aw0s4FidKYaUBOdFVWMqw79dG
mylXNCMd9FK5rr8TRHFc8lhcru44c4999fvbdjfnLDu+uRBhVSlhVUI1j5Sp/gNU852ctBCJS0SS
ZCFNUtFWn0UOsng2vK9agddC8lscGNZKU5nGLaLsDsD075DBWuQ4Z/CnrxqkKzjeeGZYMNfUMV/J
8HF1WtdKQnoxLNLiAFbtW0qevGkco/6DVtFvendhuJYUrrmPAsbSGA7D+huuAGCQgEwLGmHl8LZa
5XtJtFr26COZ0i259wLozwMHARZyZQXBqNT7pqwCz+VN7VGSIHz5a3ng1bmtf5uTZgTtLaGgFTve
hb2h8fedpnBnB6tHleZtg1qlj5NoI2y5nsE1I5GuanBkbRIMCYrc42HrCRREqYiP4aUbwOHZIZSE
HurCNFhCwDqLEIQIVtpS+CWZ1/WqSbWruvdUG5j40NzZxwAcOoBeU3wP1hBJ4Qmvw3fZ3z/hegyK
A8ouLwkzUuuXX9yewgQgzQNiD6hUriXU49sW/TeeggsjBqKcTs8vYopNjKGv89EPyCAogJmYTDI6
xsdtJhzT6s9DG7uoQ27NqvevAFBoQ2gT/gTw8PuO0zumxxHtrA7lMjt7cB6ZUn+fnojmKPXNcmOS
tT6Li91xpGiAZGD6x6WUwhBGfPDNcWH/cbHT3olndb57QUWxmFEwdnxurWdMtogGy3V3muNHdEWR
SJn4tsSX40sfqS+m+uS1g2EIlL7Hlr2CK8UKjYXWc24JKw/PEs3MORhrzkl+dpbejOVt7SM2He2R
KuTaZ+KlPKvJePDVz9GPxvxAuX5WJnbDIiLHKCdGEFtYi0Y2QCbtRNgx7VeltuGEt0os+hpLvftO
JYlXOg1QF0wIZ1KguW/gyr0PPa1L8jiBq1UvhXOrK5052IHQ8h7S4PM59Gn5V9r9a9varP+aJTXG
2bJfE7V7QYOcxjPMRD/kFAmWv5z8ublu0k9Bopar+MvO2WMUZkyRRjSIXQ8lUH6300uD6BSowa02
NHKlNtG3sZqKbuC2ZMMpFcfN0/+EKCj+l09w+nbuhTAWWCayJge3c+PsKMH6TvtbP7alifkk6b+a
qJ4IdgHH0VZcI7bgHjOl8rXwKxgS1WDnU7uqOeNtoPLUb8DwNBvuf0hCJrxArI2hFWDs7k7jcEeR
mITkbF62N4+4JRvXNm1yLZdumh6ENOYDGjL3ySNyFKRFbMEo7oy2rAbfFUnNQPTi3H4sFPR6RJTp
YAK2rDau/CuHy90UsYnVTOnffWVS6iqCAYOvWm2h9afBirXac4JYq8QPflSFc4esvHbYk9S6HKZp
mpBJsWLyjPoMAcre0Cg3jlVfFJo7bIlzgf+AG8KUYkbMQvV5zwQzjlONvX/GUEAza+4Vb+DreD8+
F6x5igUeh7/ZMACXZds1sDy/D59aXLs5uhRQ8keDyNLvXgJXxrxA4ukCOjl42qp6IymNLirX1Kom
GGkBGrFi/ZnwLpeWc8LoIqxstw/dqCkFaTONauBG/hbI7+4Ie8W48Lkt+L+RinD2Vds2Xx87w3Y6
VsQwl0aheCNhciL5zujenz3RJOn8XfufDc0MaYaqKb/JMY9NcHsQH8gWoUHX0shMHM50uPClGXv6
H6h6F+1GFcytS07ZVOMbYwfzBW2y0eEr8KkKP54kUcDvLmcElvz58ZDnt3VsXetbId6iOoqekD6+
Sw23CCh1fsEw/RfkI8iCbjmfNoBAQTcwAPaBIoeu/tllPWXBLKuuvIlhjA7Vmj8Fe9Zi4+idg1vv
apN57L1V7PXp8iVCvBp18kcgy0I3/vzXED01jrKA8NXZFC8mC0/N9Nk7GJMbBLMxCjQA6EufpAJK
kkjEZKSlI3mQmQPYKrGKrhHB5A5ffYNcFv9dsiIQieYCkf7Y6udghgaxJ/5g6cKGbJYq4HTh29cz
c4k20S0LG8qhBGHqUysUPRTHcFZtCVEYp+7TTlXXJZXD/RM2M20heJVFMl92gmuPKnGySHtde8PO
EDrxSKsJlDe3ivbGbqJd+k3bh8JPnUAr6aD8cBl81SuRWHktIqp+Ku9pWZexkKIEByB3UW1luJZV
8+xZE2Au3qqUn4Sd8J8zQ5jNr+d1TNHjVyZ4uVbGTqZgiyswp6QBM+wMDPmwrjWfdSI0zNP7C8p8
izJoFtGss+g8BefNBHD3uzsIEmNulq76timG6ZrE7ZaJZV2fPg3geAveM/C7FNsK0Bw6t94KeYa7
K/rjwynF62L8qWF521ens20TGmbhOV8CZ3I1hwvzVXdwFLrN21aIm/rvCmxj8impgiYUb0ZzTaem
qgtQuWROJKdVTKKoRosw1GSz8rByiBY6qQvQD8XxP6t4keShf5Li+oVZMJJtVfnGl6KtwoPudFew
SVZSrQLx+1pJXrDxOpCCbxH5uKd4Uo2QlAz6OF0UPLRUtUw20M27RJaAX1rEMXBRsTZP1l7MbQv3
/zKcjsQ5AY0Ws+OGqF4kBlzrg9nDozno6f8dkMCF5eLIt0pF5nk+OZe72ZusbnCEAWTs6PZTEb5T
GspzYlfws7kdDKl3+B7cGj+Gv0wHBH+CPvJhO64JPF+P4VyzHVZpZ1YHIlYhC6JwFwDk5IUwN0Bl
pcASUuarjThUcNJwKdtVv1pCEB774+AgMOQv9zWgoxW0HhoWfTA7og7Pd9EWUeE3cFhmjxbE+dp1
/ioEBaHoueBLr4UJIqWW0RetUNlDkMAa0Ucb2dYav2inrFXY5xQBGYVzW2fbjyZhaLR/ptpvFkFU
o2HeITtaLNqXLWje3L751zsP21lTx8+v0ANZ5U//zWSDwVVSOOiGdj1bn5KyQOu9TbLdmhfvNuOq
5eBf2InD2k/iuupgrOI40fYc3VvcpaouFAQxYpVBzi/8I4rE96xx9m4/wGVB3G2DypuSv4w6lQhV
dJOmRqHNRShFA3KoVwV3zMJYFUUgyGNFe/aBAWrTCfkOeJAcFXe5uG3IgLRBDCPcIecA3YYsV2DG
ao6ThBaABNOhY6dnpwC+1TjHtoThS14qN94WK7h0wMzyH76mOMawynbK2ottqzKzO6EhRguTtb4r
cfZ/AjteCrzRteFXIxkQoHsrw1FIPkFcm+4EhgoWL0xRpQelcRAe/Ol8ksFzIvmisDZJC0h42Ck8
ZN1neonOAIBsodV7eeZRoXr1l73EAByS4gW3aM66FZWJHmX1ehjMZw/2+UJAwpAJ6lo0zmc0Ju0u
GSy0Ja3WcEXYlGy6sKyHwNme3d+hNYhIsohAtddSKiw8IoYScWbBqBQBgyF5847/QZSWJtxcxmcq
lBTaF97YL1v52xey6+HO/1uHxK0nnTcjPnJqID/bde62RKiDzFHr+aprwndmdoQDhHjdw6UwNupq
7BdPdxEE49wRiTiNWRZTxf21ymj/CPN3R/vr+fe+gsOimXaMHUa2ys/RJ7hnJjKRni2yASV6vQqG
lvt4AILhlMf6ktZdRksvv1OTpPVlxY+4ps+UT+RSoXgprHGXoVwmWlO45RMPh669v9ksHNt56uKo
GWJBQl6SAfq1j73y0jb4tTyKbkb3kyFZDMvQAfY8LvE+zM3kV4N98kGKpUKiD1icAHUmapTG5Cbx
IiyYvT9tx48LGW12+a/BTbZkLG31JoCu27ZqebL52jZJkHmiphxnwHf5/6N3FtYFL/2RLZ3jBAtN
W32OU+eaa4SpCrwgq5gDEd7/0d8DMaGtKVr4++rZXYTuXgw2CUPxfK/XFKbvDRs9T/wni8p7kihh
Btw4XUC0H16Z/fUo/n3G9QlyXJIJbbXYU1DgOZNm4hPIBCo6Sjy1zjP116nDKcTVaNRYhMvvknW2
rdAAuEx8Y63xwC4CSLhFeD2xnMfIOxBb198j0e2MLtRmsyeUmmRECUjXfMgY6QUnpNsYQDNLf4sc
mJfYJ4EAjHlD1EyJUDkl7BhH99M204NoGrduWZFfliYru45EpGC0XgolQ16F1GxpWKQf5ws1aNvm
76vqP5hTaJJgI1flguG50OXz6X6IculVUyfKf0HJNvHUIsFr5qE9Kmo+I0AXwemQlJQapXSj8s9h
JeXX5YznMQGLGfMbUHKokzXUBurt33CwQR3cBmaW0ryLxcBb4X/d04P1tDOE8qTN8wPnLIWcWHGm
5X3+BaEghFfFGyb8YPKLiCD+v/CRbv6qMdkr1vl9LbK5t6aCHSfnudD2uExwCt4Z47WWnYMK5Md6
aeTq4vUdYa46/bx3bDMiI5oa/WBEg779jWALiWNPTEy0XGvL1jcRzCECjLOeS/vweuOjnJ38mR0A
+XUiKe/2eQRy7J/RypxA3FZGBwMQLLbfeh4JWGGYQ91di3UGO90paFFc4LXRKU4jC4/6adFzAyWB
zglHi1sFTrmykM9ZSnx646OxSGp6BE1H1OVIt7CGIpdk5ahjWGCw3C1b2g3eE5RoP0u55AYXIKcK
qKqRasRCUBYPqey7u9YvAucE0K4bwKtwh1XqrvCxA3Wt7G7aiUNuIzLVavoQJP6xzKpp0enuj/HY
5pWIR6lQUZiSiXFl1JTxpmmccU+KBWHIn3VSv9J40stH3CeoLG6PL6vlLeBA1D39MBjGDQJ+UMth
oQFnE9bgUQW1f0ASGnzKPUhuBC0yfHeBBuY2itW9lqm7TAorQZ+bl9J143MylrEJq9QUN7OJaIA1
i6DPSmDg6QvE4Qv+ON9hSq1Kb+Zpaap7+7+M5I/tLKE52PP3oz1KvtxFktvxVU08tmQ9LVDO6Blm
7h84SOZuTe/QzZT/d+fx8f5bcBWpk0RknNc9cmRocDslQTUkgB/P8jGOxT8GVL2IoAfC6InUhSiS
mYBmoIaam6DV75RXddk3vPExDVMqgUTsPmSujHv0S4TZy+t5ruiPy9/EL+ARFnwvJBMsvZl7AJp7
N6Cq4bKahR9MEGSaRwRIlGlSd+pxv1RcB5v65S40bXw6JIp0EWPsi/BAYMtkki1MWoDgkehQzI+R
U96P2atoRix2QaUAxz8Z6DxOcbuUMkedTnNX1pby09DPGzA3DqvBlzU27SGWesY7htrqPu6sDQlF
7fbGT+GvvWGsC+IorrUA8fOHrqrRahklC9yeg4tIdLOYy3ObGxmdnkekgT7jhl8CO7GCr7+ZthIH
M4JrfkztKoHiAIjz1z5okC6PlJ0Vc43Y9GL2uWjk5qM6T74KZjzE1yyGQU89jMFdiphz5hScCiN6
4+u/aVBqQHU1xcnF7kXbwS5jHIXz7qr7Khb0A8gBwphcFGY3svSx3sPI543zTfKec5moH/wYA+Qs
4q/QsdiHtUNcq0cOqbkuCYKILDwLWVzBlwGA+TXcJmn0d6zVw7wOrHJ4hTBwjpzX47ibrszEsJ2n
YnHRTktNk2u6M+Dq5g0y23EcWYwGKawGfdXLPZILBHL/8rSfD7yZNxVItGhJHSC9P0tpYjIGU24Y
mHRTHagbgAk0+QDy0DlvEKPRx7s1EgEsXIEIlZ+p+Dc/KBYgD/JC1xaoiG47InrEt9yo2KehP+WO
AlIdGK8+LqXx4bjBcptxPedRL1JGzocLBVK1nP0eD5cEn2riKt6ZKb4zI50FNaEXdAbQalmAtr9h
Q2vTrqgy+lKWmuQSqKcGWBILEQ0DEQe4Q/jHZnTdEJM7YQniDMM4rDwvKv5sKZoKoRWqcILEirFP
y0inz3vw6mtpCCN5fHCuO9pijY6hC0Vatk+vMskXH+lHkEWNiRQwiEcerlsdn2+GloUMzrzbjfVs
MZFyAHkRUtUtA7niZLurGV/TSFlke/7cjKXOC7jNtlEhXM6HQmO6KCNvJBe+eO74Kfc5UNvWaKGQ
VxCbsSlHdj6F7JW5uF4yXpGbI8SrZc1PLVVjOk2+dn6+i9W4Ss2lvUtKsM6CQ9lRSOJUqNDBjQGT
C9NrIKJ6Tf8DkZmCqcG3zCYkzbyl6Ta001AEhfaBCgoQZ/zwScAx0KPbErb4E0aVgNBO6Kg8Ixv4
JWz0nLNysE3ndyz0I9BPpcbV6WiMO9e5Ra/6ULozVtyKW8URBuMo+D9Qv51YL+dHZRa0i4om+6BH
Fi5a7Z1QfLFkoR1s5K0HLf8x/t92BLYiwT8sKMWoSXU6FZxh2Yd9uDHpPFl3x2rgLilRJv8Dsr60
2g0T275AnYR5Env6hzCxhlGtyPJ/30ns9sMFP+AYcDF3N3seEztLfu1VKV/TqDh2dIS1wj2Bs76G
r2zQyLE6PAIKn10p1j2qBlCIVIKISbiKzW3qiA8VHi2kv1DOX01BlD1DFmFoc+tRAllgL7tGtozH
6ke5SUorxV25UbPDZGED39bWLsSyKJNaCB0jT5KjmQ9DiYZW6mGSNuuyirRNniFdfmQjzZQpUxom
kgKrkXhv/CFCRNtG1L13fr6iOT49lo9oLbIRaPHnPKUSyFGPFnAqWh8AeN4CQO28nBpS5Yj1Ng/H
+OCblhSO73Pp4QA0NgyR59Wg4fuKXG0xhPSAs2ASQLWob2yAj/DFNFsDCtV80jtjHXvofyuJLE76
7Y65AiY/G4cjR3RV9jVCChWwT7xHWy2T4RlRVqU7d/MPU4ce2MdzpA74cXfGbgRGJo+MeQffsuIU
VJt0X/V8qT9lts5+ZCpwVG5RqxjU/ZtKjREEfrnOJHp33jMtAxa+BlJ6hC0m2tT/Saj/sJGUg4r5
ROpQUhX02FM+CaACvTf2tRTmcK2Do34ORsFmbrAR4HJvgnwxIqtCw7Ab/uUgCMErZG2dHzYfPBND
AmBzcLUXOdLd8lr4COEjlnN3r2kvqjd7LTOwAoetIzz6ZhXSBWU4StCv5u2/oS2R15f7juNIv6KO
ROWog2VELHvzeXJfMLfEuwBbwQpTDMRxJW8Gx00YICs0RJjJxnOa8eMCUivgU9IM2XCTPXae/2Pc
mb7gmzn797L8rgZpmiUX5yBOy2nT2pXxR6TxPwVnhgZV28EKJun4qp34st3nd7xn8RR/nhlOkIzu
GY0UuM+VJNxnRWuWuYqJJrwdEo3rj7J4YwHjCWYZ1vjKPjJUn4RORRVtHd3PIO3McY6JZrSJfxBb
DkZk9sdl2jqQY/9WF7LXU1g/23h7hrbgahdcoic8It7lve3SkJezlxIk2oUr3MNk0RohvIM53QpA
pnH8ZD1ZbxyG/vFrlYHwFfX3W4YKLa7REqFOEtmFo2Xd4zZ5T021E+a4VSsR6AZ3es4H1zsbtjlj
qVxEwQPSloLw7BfB7ujGtxpRxIRCpDw5WtgZ0D2bULFNCyoZeBV0PYhfyiyGoggJGy7eBU4Qv+LS
5MduiBN24wPmKrQPOL14Jo5pnT3m5vnC1kQ5erfKiCiy37yfyoe8mw4Bhztvpl21lsQ+FdbvFtz6
cFORWiFTdanFmTyA53Lcgjgp64I5C8QEtudxEpG8B49ps1H3Xv7oHswW6W2j9FR2RKfbjqNVcACF
LN6U8noqEfd6WpLDfxIvOJpWs1bPxuRvycoyDWfDXOmuQPqgHmn343Ioe51VssLTQGzDy+XJL6Pa
q10x5E4QNI5kjeTRiYpVrorp4QK77xaEH9jXD6UQdrAGb6NxDWECL8JVupA+AccSftZUBc5uSakU
deZTGD7KVo21uAdBQWBzVbwuYkIz2rGTv7itTrDssUCKR3Dkqd1iubk246WO7xbyTmXdT2L5cXwt
SgvCxTEiEm6btOgfAwJhWQcxzCNvkw0UZNV1lfPBMWObCbOxYX0q4/bpbnFCy0H7k7qy3nr4zfSP
kVSBg5nVSKSKEVjkG8uxhQoY7Q0chBADedMBDvnpcdqtek2dLJ3Trhdx/Xt+YvPVIHGoB9H+U+iz
dl658SxfQ0L7LanPnqdFNapn4Jf64vQ2XL5ks3Il3+3JvoRiYQ7ubSkagoSsOA4WTV5sY1xnp9wJ
PkiTIiYRj33eZvP3OS7oTQOw97ZvVbJZidWpMarbLKekkmSZnZF8HYVMsGhrzOdtbh0Lz+yFqN7g
I7pzJA36VaJHRtuymatASO6ECUndCPJIng3R8Djpi7qUWKVErfDhmjavnI7BcCusA5+Sk+MYOzMe
mMbQ7Sw1ly9ygeAt8WGbcHrQPL/YDnRTVYRJlHrNo2p3fD+7MsEIpWKJqJmzH4ApTsns7mBaUeP4
hrNTnghbweVPGLUJNi4hWS4/t3h6nRQVxwEZL11dmDPnDwFWaX9X77PS47QlgT0GF2eN8vDKPYgU
SvhEFvS9J2HCmhQQo/i2JdeXnnqeQI094tnsmha039YQOCPLU3uopEEf2Mte5yCjpYkLqXO8prFm
bdnmMXIIWyBTjUFtEAou0EL0UuL6unakJLICTWBFDq+e3iQcFVYIYFUckqbUVwqVAejkiHgoXwSA
0UkBMbTI2IlKAfpZUPjIrAjArXSHCYk9Kvqb1beZ1LqjvXiS4g1eExRnvTrtFzwXUnsj9KGJmiRy
w9qltaYPulXEliDXamta6r8v4MPniXcyWbznv9079F+OgNiAGqfb25j/VAI76EMh74zE617RA9w6
MAZLEjL/H2RpfR5Itn9IOdY7q3jmuBWbPq4We/Rt7t7+Kk0/ILmzVGwXWRoJEDpF9hOjMvScvAxu
q0fLxGndpAtJ2JSC8PCDuR2DikgbvV5kKXRLEvW6h9ke9WTYgukIqGwg1LoIeayqgmAUWCdWtXX8
anD0ffvTLmWbls8sF0Uza2a72FdVUpTT4DB7Ox/h3+qGzLhTpIRgLJf7umWeNGe+NuIbfOa/yhrv
MbUMf9GCimo1u6b7tP6i6r96BmuumT9Jz40zKvg85dTRnl7qMjtWhit5czADL1LT71btFxccv/JQ
uH3JjdENNSQDonbhACJofso9s/rV5s02DMY3gHQcvymd46hO++SRtIwijfqKkFL4AzSDGX6/iWif
N5i5+BpnvRZBKC1tvS68cP8SazBUvFZw8AuNJY7t/J8Xvq+oQohyMp9ERa+nSGwmMibUxLakbLeX
aiMQAEMjYKHsoc2bBEQBy3oK81zGsjPqxPulm/PKk6KH+xevgKErMS+heEOMaHHDAV68mH3g8pY8
P3dB8lDLzzz41N+3UWTTmzo19oGZ7bWnrj4YDlPV08KN9Wta5/dy6yiiPiLXiOrfUv+XIxdCJdSB
jtombbFHJHiVjfiYFcotoZE15zCrcXJkb++snVfOU3BE5Xti/DNHglI1o0fuUjsik/1ZWqAmFvL2
AEdaV+P9A+WHDzwnc+I83KEhxuTdm3yUP+OORymnYvWxTOgIcmMWZW+DFxfLY6h5LK7aiAizfue6
xvdz7Pwh7JeZlmLMcsKJ+mFN6ws68BV8qG9l60x/b2xIy5qpPexIfrvld1QVIAgBAUxBupSb+cX9
NIiv9D2PRMfY32w76n0WKBZJ9TewuQdWpBQizVtB+k4ZdFVAPZwRtfs3cPDS4x30jz4F0Rhmh/mE
HL4kjspeFD04unEgS2HhUE0oFh0x2vRkvak5HE+8Y72yJWQmr2LMqQCvhotvUUxmm302TJQNzCey
BHano1tBDduGrxeVx7BUuZTLekkPb0j/538wywsIDnr7M87eHpzCq3n3b1qhTf7KUHkJKMXTtKMq
7Rg4b2knJfEalRQRH8qFxud4pnRRLA7zlA26lmYF1Fp3jLSkS/wfV2ZD5MFEQNz/4D+umueoCt5U
LbiNyPwkPjbJZQSrhcQK8hnwlpXRJGvK1Y5e/BBeGgNRXbl7xnrTIIPtDot1qvrXA0J3Tr0yIoI7
gKLo2MIA8xE4zJb4tpdgMpYUMUljEKlwrxk3xTaiv9EjT4djJIJCyaRAdVEo6bDS1BSzEzMg1yY/
m+ll2DmLnAupVXSucJWBPionXeXTBj3bEEOU4O7OMG8SBWZuLr3PmJ9h94NMNIGJZHrj6jfc8vFq
wXKSyqvG3AiP9t444JcQtl/I/AmfRm0pfm0W9NmergoRL+X2Xy03ES4ZmhTGsnY61Bpgpz1CiE6k
6PUoX5UyXWD/GRfdcNHPTvgnquCdm6TPRgO1pxt+fBPZ5U72iRYv8sUeLve3a9xJgmKDADDnRU9v
ilCa+lfDbn8X9mBRDZ7NzndOfxvNyGKU1RNVk7dxTgdKZfTO08zFDDLZGmKnTt7H+KjZhh/MP60/
eKYeY4JG+1CierHN9zgZwb73d2GvJ2UFwq+te/0UHh77JlvS+KkVd1MOmfa0SeTlj4nOHvTEPX4+
6YcRddif6qW3O7Kq03a4pfirixPz8XnITgtB+WqGIDp5qPDO/oerNEasSDJzw7lFn8uZBEgq5S5I
ksVSrNJsHOonLgRxX0D5sicQdXUKxhlLvz6VdjjI15LHfNuADFUgZB2lnIo1iLiKCPCcpNtmjq2t
4KkbffK8oU5ydEhIoC39wEKbUqGhwee/j0eiy8k+7YjAmeYP3s+FHxQFj3SascHCcZ52dEbp654C
BmVzzm1AlV0d/4uEJ1POIiGIE++zbyGGlvnrUbLzi6A/B4Cd1y6DO/yHAw+1qGuqlfLuvPDf83fy
AsYgDyOwmtPw/vxzk4w9tp2KO2Cv1XO+D3owd4/aM/KldQwq7V+YRXtoeXzd7Lol4TO6ipPkXArV
fRlMxl1VQHUIr+fKMJlcr7cV91szt/XDs8hoxEBHeCpklItAcncl3UnO8ZAYFg7Okx8waJDj0Jxg
vSA/efRVAfid5rmbY+ZhipWgFx3TpJBeeVJfspnv4NVtdLAT1mGr4ZSZbjf/EGmQ0i4DuBa19gGC
x4gBDgZzPZInqML1y7yc78o9XnMv7D8O6UBOdxHvIFdUpLMaC4PpVj0p0V0bN8JgWtrNJyaWE7jp
bAbzsiJ8ylee5umjKuPqf1aMlyDfFT5RL8qLXsiVJ4/gpbSuDwQz4zouq1H3DbCyAYbXHakrOy2c
bcFTw3iKxInCN3x+E14D3XWO8PIAeeEi9BV1Tx/GD3WJ/HJEs3RE2VVnpCln9LMIQEjwwx9MVwFL
dfs2ZNN9QGI0sVGlFSqA4IkHtqY2tvHm+DFX70u55j1GLMlRJUyjzUhIL+GGgiIz7B9VqfU5rWSE
kp//H2OnxdO+b3A0/F0mSQ4DrCY+ve/VKEX0coD8U/Uc74NHcNwsN4DSb0fMbjRTME31aUbnUDaD
0B5ETnUWerKkW4orNF03A7ftpPmJ6PA9FltYuV8nG5EWH6c4RcAog750WbHTkJgdJjw/DAmfFHGj
ILfjwYJurAQTTBcM4DakVS8KJILOWb82S/weCyF3QI7+4BLJwQrkzSyj709TC2//jOqoA57Bp3AS
56gHJ3zrAKRIU4j4Rqqp+rav98/sLH4p3HLmymgX7dwBy7GefFcGfvzXpDFhB2mwGFS8D+WL39r4
Dav+/94kjh5QZaKpxSWQYidI6OiwDdru/KHB9Ey746DDi2HXLl9XXswzPScNXFjKAS10jfChyLuE
tfxmX3uko32YrZE/1pXo0HbxEL8qa44l85Vg4KdSQYY5k/PUw1nv4vOV7O3aajxpZ0w6D57B20JB
0MYw/NC9JXyw8uk7r26h4E/dmzAUR8LjrpOBsXwpAy8wHBc1umbLUMIt6frWB3SkZdGV+U4znZX2
pNg17ZKFEswL9V+dxiF5/KloUdDbChZw4h+kmT2JBJMs24l7kB60PCq82/6qbEHS/LX4/CojBn1n
PLQg5da5odCfTjcsSuPNYtHnPri7tqOSho6jYM5YXqYOPxsy/e8TgFE1dGYJQL2+Uuzbpd9ZyzVu
PFcTOK9Xv6y9WwYf18YHcXDKZavFtaTMWUwtte37HTH9+GHrPuEQHhFU0gr3QeP93+CqSbBLMQWL
IUB+PLJ2KDONmcTuzXEyaEiXAFMuUYkT66JMRWqTFjQ+yYtKS8pNBU56wQAPiqCGB1WuN+higX09
V2xMap8enADwPSHWUQd+K6NOjlokjPCfNsrgLema66Gp66Eay6sCK4d2VPILC6yWjGoSzYCH6vx8
N+a3gSLNNHcZlQOdpEXRBs0qzUqOqN3TSiKtfh1pry6OjPYQXXJPWslm4cf+ZgPRGUsOMSeDYj1d
ZzYAByJ14kkdL6ykI/gZxPnhC3TzKitfiUPmgpjRzOrchjq6akUTlwnuABg/Rcl7ld3ndYZaIzi2
w9BxJjU6w3L7B9ndyNprGZ1/4R5U4xWFcH7bEMK6/dtk1SUpo/F5b6eNh+LteKAfQRf0SLfknm90
6q8s1O4bA/Ge65MQSi7AWAtEO73Yiysfu9paafU3vq+ziU/Up5JCyB6OAalhiJfhzI5OANGyc921
qWBzwfdOKpk2fijk/aqOyUKgtF34fTQ2W1Z55R51pr9vygK4QzeqdkhCFM65r/6YRLRTf0Q4bfac
dffsjpDlJGq+XloV+C9zEc5r/eKNFo3jF9e0NeiEeg4d8yv1WaRVRO6S/9BEvTJN0YPuFXs+vlaa
q6cxqxNu21uWTeuVgTmlI6CKkYa4S4fdq11eXLp4syscz4334p/rFhDeCz3VwD2DBr1cgOCdDpXG
IWOWG9wyVRh/HYgcnfUVxGHJFTv4+jmH6HxACRmK1hkxbbBQg3zfYSKoqlqXF9CIbcekKAmPrg3t
BWoN3DE8NmR97nYbI+xvKFbAu/JIpehG5uM0+IAhn2eZ4c5WeEkiOzVExh+yetQAtBNdLV+mlOmp
AmdwnfF0nrXJKvCmxJLkQaUPyZxKTWVk88MKMck5U20s44HMVgq8tYQ4IEShScCEYF0tdz1LSQSh
uQtwGcpbRywVhL1NAlZkD2ncJScJP1tlrwjORQ3SeWvC7RhJg4FJCt3kHtI119X0KrZukVq1H8xU
8XlQY0gj7z2QnZmFPVsdvh5dWhzFeZdh6C13b969HdXLGAncgXLMvt+fo36qjNie6g/+C6Da1b7G
t1bDWGPi2/kPCZbW9FHe9GSvhAbKVNc4Rpeq9CjkY4hTaTDJtVpyLxcSE0sfRZyd37c09sLZMTKf
+d1YbaGaIbzMnNjvgOqIN+3j6n9z2QKCAu2j6THkSmn3a55vkXolzzSY6uaQ5zOwQ9pRUlpHlR4b
rzdUW6eJy6rBLQLQm7bmmVU79lQcoEoF0lTIGyylOZH0qq2aAof2WpnTVLHn2sZ4Zj1vcTj2e5py
ZyRo540vyxcRYyVbuE/Mr2tP3BX3Nb912uWCK0gmsHAd8hsCQ2mVrVKDntJK6uP9UbDnxmzkmRCa
IvTXe7dZAryBUkQmDlpfncKUzPUKXt9dI5ST7zR2SJFZTby18n03Px913+qpnuZ/mDwHtduFsQQY
yvAMtw+X7iadtFPHkwpZtfKs5cfFyxZRJvLUIvCZZ5sqkf2kHs54gWK635Eafq7udqSxkwGUMVSn
Tt3aZz7lzqj+lUb8WVCYOgr7VK24tCD7KxTRS9RL0wTECbNtGdHwrCoNpdAaJvvyjif3iz/fiFuG
1KzjWJUNL3fgJnBXgMf1RDntaOooZMfYDxG8RnRgHnyMMXngRlVysJib8WXioWG/sHuOYBrZzC+/
OTfZNEgEqd53JjonFobJN4bDBYRagYGHQ+O78Sgjnm33c5oa2Nuxkd25OQVwz2oZWZ1ZVzP4R5BR
RkOKF5J/UaKYS/UhJZgGxVeTXbGWTCn51sdA5gooTzWsoaN5OdDHnHstRPSiBugquT5gQ0LKWguR
PVBCF8QNZlm+giQJ5j+SlAy/ddExWE2GO1K/WBP4N3Ez1A8uF/DMDGh1EapRk1CaBh5lvcZER2ie
a+4yUXKWBiWlG9iB+p5dtWN55nvHGi2mb4VD+0PykU9WqqvuvHEQx3HvXszk0aIWPln5p7vuD5mq
lpHINr0H38YfX0e6vK4l6PsLBZs2yGSPckdSWWZ8ps6utvetaeHeiUyrFbdv+H6H8sBNDffO1xnw
17v6UODdWzmtfvhJKYxZcq0cA9MxdMOZYnjQmTWkOqlVjn5VyeuLBlMD3lhVbINSkUE/Py+x3JhP
tXhVuSQKJTkRizoZugl5ieZXtLFFb6fMUL7hPl1nH+VxxvvFPOYVw0hM7Z3jt0Wmi3wJyaBnlTE6
liSL74eB02u3rw0O69ia8MrjzCdumkzGIYAW6Wouj2HMNo7B3qSDDS3UCUvJObYPxX3vO38q6f1f
0zvv6fw22ctuWbjx56VaiCE/yBHPBH/66Cus7sdynzZ6E+8wBBqtAg1QjHI1TPMSGaPYpCjUnKGp
ThbdOJVKC1SC7MT5FOKJF57PzCH5x1hDb2Hf2VciFMqHUvuYC7BqoQLKgsHQyva2T7aV9FrtiG3A
atBv2PYdvBXJxOg5o7O3Wc7es2cIRmSejFlzV0qR+KzqegcwVoBMhQtZyRyovNJ97IbQxk/d5PyJ
u/jUJAPI4yfEaedJcB+8ADO3z9qDP2eO8CYxZVnZB5tlQDdeNmWpGc9o2SgdgyX+m7SKrFwaKVtY
ildFd6DLlgYm/Vo6iAfoDJfKCE7MMNhc8iCOuIDxKFnaHvE+DPIKwxcRqRVLV5q2UaZJZPb56Cic
HnQJLD8lWxrTzaZfI6KYmj0mtobh66Zfm9n8DiZ2nRKyHH7nSvBE1sMCikFQU9lrJu2tPN7ObgH1
aLzf7YCWQoq2e+Zq76Bniv4wWl6eqyD1fn0RJcoqZbJpvb3Sg6txKorAWcTtv2NvWbnO6E2xIoeS
YCr/JidINbEb3IFqyKxi7KlYaVRsic9vra6HDNDz7Q2TrzSkVGf6COFFnNR8d00fWpkor+0dBi+S
m7LG82sSvq7PNPWxmw0f6D4MevyuG/dIJuycz7eAQ8POzL/fDSnQbiTohfLPU0XUwUBRtFDlJnHs
JmZp40QkZzpGG8JbsMpwkHE6PJI7lID0Pbb+Li4SL0iDudxxaJgFW2sWcf2MMJnrKo3Lh8MThFN1
U3kdEd/sTXOEAUVilrUDcvmxdm56sxiTI8YQ7B2MIioPjBBmxXi1klEZ+S1qlz8SzfQ6m9rS/LO7
Vy7U7EYWosfaWmZUvy8n1fQvOiCK+xRsTq7SQg+RkSfKISUCoRpytmv84KyVs0E0gpELnrQPMQyN
+EVc3wCZQCvVzW2Qo7A8J1ccm7xEFd8pM5CYBWCAtPlJWVjn5M8GLmEa9TGSgDRB81hI4Kfz8VW2
NakDzsTXCq3TEhOX4ZcTqmXefdCgqeZWQE2eCv7XzWyKuFVjvTixlk7I6eAmryEix8+fAQV7R2EQ
TH9zuKozEp/u/aVqmYEdj9aEy1eNcJf6DFWbpjNsaLTIqALIOL48cBYFm83ZAA8PJS6tfW9ojr7c
GWFAuFbEpQJ3IU8cmfU8Vm14ccmTznK6g/JoDC9IzyTW739vpwu4I2ZYtBoShnanIFyB5tyDLvFY
VlyvUHRZi9e6ag2smJRtYczu8jvgFjx8Fn4pvrkZasFi9Bx0lH96gxdgl3vFe1vXScDWiD4pYLdQ
VOOfwRWSJq/kXuE42ZtaeGe7XMiYtXdLLkx0FVtU3K/EsuiuUpXHOgkUolQNcEyY8//AIdNpG5PW
NAi2vnMIWs8zCl4IPRL5/LH1l+ld1O1MyaV1FqxspzF2LvyZhAdK2yViTMMZgxBykAgVztO+LA6n
Wy6nEUuWgXxzb1ltFcbyffDHmtOIyS5HrvRdulLfPDzJCw98UIitiqA+a1dhUg6F1YdHCyvHafQE
pLj5EPUUpaMUvzVq6MTUIU2/40pBqCcz2DNNVBUsfvMk2YrbK5gm24zf5u9QI+/bWK8n4/8G7o1C
dg8b1/VepLuGJvQWqzv3MsQt/2KJ8BmHwq57tWMAVbY0H+HyXIs8ka8njQFYcCzY+r8L7G3sxlkw
HfoIDmQlM1sgSKF738D+PggIAcmYut7WIZzG9K4rmPZe5vf5gYLLGw9Af0KZJhEBfv4bxwMpTR2T
PCtfv0kWSmc+DrQjU0wmcXxGemj3qHUM+tiVmD+tHi9h5VpotLfebaLJVH+cJ5ftKWkb9ELstGI/
ajAijW+TBFswTA932b6VHwX3zffNNL7osKljMzIkMHYzolXDh3EDSih5yvZZufqzDyHQ/BaS2QaZ
moDk4vBvNXK/xQ/11AuU5HV8qUUdH8QACJQbv4KvlnKmOQ8MyD4ipygu4sSdq2Z7U9Qhb4IA+rCw
g20Im+zk5fskNhS2CIsBwkuu79JwEV6Ns0+DxuMtcXa2MsbbM+vCalSzibcccKaP+UOcOrB+L+rG
lGVzHCqn0IIw08fHsO60+bzUltFee+wQGe9xtaFAj0Hq29JbAXYro0VZiWFfJGhdhsvFIaDaZh+5
Vi1AId1iEHR+L0ZhTmM2X56Ft0MfV6ojWziEYkDJLPZpbW7UI10TcV9mk+lN6XjzIufcqTfpBpaT
4mW/UcMfaeLYUeBRpdtl5ukkLsdhptoQIFxgPaQ5T8MMZ6ZaZ8aN5A/0NqbuK7dJBXLWFblIgRDs
n24Oc5l9SwQ6pWBS9v8nINeYxt/lL/emJjvcEQNw784WysRDxoKJON2kPDZOJHGRnxCaihc7R3cR
B0IiqiGUuINQIeXLsK83vt001fh2GZZbugcD1/WJcSSj9bN2OjtUjTYJXVPrb0NYICioZLf3zsqZ
jAnfVuh2gNmII6DLlChuwe0FgapY5IJUAwckHbqV4vsRtMCuxAf6FjpKwdFo+dMUbK0+fce/sZuJ
nJdTSLpUD4x/XRb5vny425Pb/Y6CUIv/5TPO8/Lib/us/RHGNuT2JRrbjY6HYOmIPqF5+1sP/bKG
3MgCDlXE8KxYr5qpGdIjhJ+EnwL8Aw9U7+z317055On9IsVivLS85v9jxD5MhYys7E+kh2IZDgh9
5o//dRmLyDIjTLQ2y1gWciD2SvWBYWo6o62hXy17i0mWEPamTbUYtWveXqnZIpr/3GqNUmuYOzoC
+Yekn8+kDsmmwNnllMFt8uhqo++mbXPXjquTYL3XLiNBgvnd3mTcOhpSTzHB0qSHb9hAgmh1F5Qx
s6SwEw18SoHfXwtARjIDSwz7s/NW6JDosEKpUb+STF82UyDgW6lQ394iOwA98a4NCNhd6Y3uPCOY
Av09EPY2t+hid7R9J/N9XKXtg5/lPpUeDbGwUHdnDkpaX0AWu0R3p8OZmxSMVHS08C7MyafPLlSx
JlHo37QaeM/EY9F+xDihdGhLpTcgH0c6nlFMDoCqg4js1R5uJCSIeyC4hK0f1j21PgfDFNC/t+fN
iE5ccMF6n5ycRIHM5BF+LeMFDReYLQxM9I4QX+lP+qMBOTshNPkvMAUsgVJxLsUDDZiatJ/ccPVp
bEfycUAQmfdrRLmuli1n2R6Ik29K8JjBqAYzK1D18GWNjmTE6KmBGga3Sf2+MnevY6P9TvDBOc3m
Amamo8cAjcE+0WPNC2NNlkFJUSOYRLOVGU/gW5uq84LLrfacp2vPsBBwfzLsFzHOJAh+rTdw0M+D
s4Qe6gFFPpIpaiqRV1ECJHRQTZZd4TxR3H6HT0LIcOlbie7Q2ZZ8k9MdRD2bT3/vha2usFSOflmQ
DIK2D4elxF7whcjWehqNHlWgKYlGxWjGHwyKBbSbr2lVOVe3Rn2Nx98hpufqVW8P/3Wtwv1B/TK3
ercbjeVvcEXhTZ+jRZRK+RFx07A0HvtN/Mor/+C2Jz3DcxIBYa+EVyIsEolLxRcKKwzPCXcB5YQh
LeKnPjIXp7ISuVKLuJQoOO/ygu1voSFoEaeX7j3j+nR1AODpA8hW1NNajZyEK5BMhJ4BagwBXc5n
yAfgG+YJbhZDUI7rwQELtJJmo6YV+l/jhVVE/khZp9gdiFU2BsRku88w2cJNAG2oOyjr1X2u9CLN
HOUon5JvqOrLjxOxIZcVJNBzF+ZFr2qwXIRjRk0KvMKIKR7gmrTFJ253bGJiVqq++RTiXTer3QTk
mgb1+VJB+p9BgudaRBwPJnbUn50HmBpVfs9FgIXCC+s23wVkWFu6dzwkqaQAxMIh5H30hG+l4xgA
J7DLFfUh33Yl6AH7JqdmhI8TbzlLDlFpvAnXFQXMDEg7FrOASDuEhV3bX7SYwxaSZWLjMOJBJDJm
ncx4ygSF/3JDtqZHwb/5hPWadLwqHjCC9VJUNadrfj/2Y3eNP7pVyyn1bWatjcReLzDg0sRhVlV6
qbXieyURKyg9JYtW9ouc1Hhv0MEPxN1GOwBi4djOZ+ZXalT30dmPmkhuqc7qEOaokJ3g+j+EOfTV
QjM7X4eET6WoydedXqXBXPIK/keADc5kMju2uYIBfy+UduwGSyHfl3ENDDFfrx4ZnjN2s7tk2JUF
J3wXb+f0Q4MJkljzZloxNYbd50WqTLrQEIKJ9Xw2bmZv7cw6PamNzHLUomg94gWyslCK91gScbI3
3WP783obMHHHFGVR/FCfZRscnELnuvlpNgyZBw0dQxyQtVaSNdXMnAXWOQ5fZ7VA4s0eCcvHJnbt
9I6R6JblwOl/jv2J4LhCIUCgyNO9J9f72q6Q8hCq/cHI7fZinzSePYjcsIdIO0XvzBcq5iXb0yoG
tOfKJJcU1yoEb6TvIMu8buDm/OMlJuJFNH3KhxSzxgbKggpqZtFedYBA5M/i5xYo9KFeCb7pop0f
MXflaQlfA5pSm5XQ8fw3iOorwaB0Ua/W0N+HdsjEsKuW35Tq5kdDjAFA0V4Wq0jCgrxK0Y4H0QY7
BXOj7LILuf594IW/EG3rBwgC/VyfZaZaH9gnyIz2SBoIVVZwpStM9uFj3Dy0SYxeYg9iTYBXwS49
mjDm6gkN/2hxlSq8qjm8vLyENEHKfSKp057rzzB3JzxeCJFUiS+eVgETwosJyLsA0tWq8S7Glaxd
AsXz9n+v6jnxMKlXbRAPCqGIZcmbhZmbrBcBGotKvxnjyskGj5MvFPwoidEMQJisFASHg9vAEfMp
16bBcMvFp4+B64O+WQVywYzmzqET594gN5GzOZij/QnHjEIHIC4ay131zcBw4mZlZu+76mBnq/+a
dbH05JxdSn6iCprQhqu+/HaoxAkPTwXOyIxHscvGZVCjZn25SVmp52tYYg2Qu5F/jlsjiz1ISTOG
XCTF9AjMGl8FO0aW0Eq/GVXIV6a4sK+chBcCpNcOanz8Sk5ly9pQqJ2ml8VPv+mlDtnEyD+sHR3T
S//g7NcumbuR7MPQp9GprwJ5mbwwxqZA+1bBvs9ZlhpSqOiY+9/KoFDyYGn/RF8TTVz2tN5OXE6R
R7AiDuPCBQ4la97P+73AFQ3SHRFg8h/lSjn+qforlCqdRXLc1k1OSw5icaaj81HUMFnyuJRlMvvP
3rm8gzzclgKOBGGDyt5YKnL0pZXKCCCeh1eb5DSLtXJcZVOzfIdFbFnC4twPC9fhlVvkvpzQXGLV
r+p3v3NQgDff9dn6mBjCnkAxZfEbVjXaE+ONdAlFHa8B3QxWDuFF7Gi6cKnWP/5ZENHG7hdWzRYu
ZjVtvWOeU2zXpTR5WiqsAR2G8MJ3gviUkCfjMBPZv7yMpLUp2nGwMSc/U7aKoQ26nHhv4vXD4ahX
iOqZ4MfiwoNmgqAjERohRrAj5ckRD4+pwqF1CrRLB5KucP0idpe9FiO1H1RcoV45F6OCuoQkGPJ0
4PWpTB0rdto8J+qOpR48XtgI655/5VXBO+oSOk3FlGACUh9yHg59VtLaNxbfSbFGBQbDDbvBvja8
CnxiaQnu00l4tew1XfJbY/tPCNEp/RvM8pvsEwCjG9X6gMjQ19u8P2/xakBFkq1TOLymQNiKiGQa
+HvsmFTdQxRPq/0HwO0JdGo5JDsW4vcjLv89s1mwDlQL1XqeQLNZoKwHY/JGBGouffnCIDuhVEoj
QU+aWkAChWs30U9+4lggQtDcu7vGYr2WMotnD+qn+WOT/opl9pC7N/GvkvcC0DKGyov8TEd3O1l3
92A0ktwChQJHp3GXfK0ElDJWgW1tRYrDfdq6cx/IoWAYwD6Fn4WGLmRKXZaKE8GOkHq73Y9h52Z7
3YfNP3Drq2fI1YqKIUPn/L6n6emVJhdkK1VLFq9nVB+Cq3FNyipreiuzTO6Uzhs9CoZ4LFwwhZ1Y
jyfHQJEg0MrF032cEmxuH1NpGQu8bizjxjeTUyn7bbrmkWKl0p5g/3Et6JSqAqA1thHEa7CdJ0QO
3z4plcoT1xKH3uDcNmsDNGuXxzMicxPuwy60iHB/9p4doN41FHQ1MUVgNvgx2nl9aj5EeEisKVUN
b4XKVy7Vz4/2WOKZ0MPkETjChoAhyp88TIQmriWSCk3jgMQDpWPKgwPUmIZmVf5BobuZ0Ts870fb
SK/uiUKpusbj3Ym6odFYecyvJjb7UKjj6PnKQYWps77rWcmECKii65VNXHmAqZZB2nyoHciEIXRx
Qmd9JSc7roQC3YyhHR1lwyD6jiFpoRpHBRUEk7r2OFsEYCzCIy9tpvrCVXEjwwDonBxzuG2erU8t
VckkrOi1Uy4nbJrTQun5apazq593ecQQM4Qu9vWbQbXZt3ZnhKc17hWLURvvCyS5mus8v0KVTijd
03iWHzcdg/pvv9/gf5s5HHM08KEKTUAb6PhURUyBbN+bNBGBtY2fZqvbCenIrMBf2JbrGmGW0/F+
990whVEDWELpyp53/C/QbxZjgkdq4BFCgtEeP1CQF4aOxZ0PtMTm2BcbGSMv4y/z2alLyH9hTPEC
F6THxplZEYAvKrqoboydixOh8ovLXG/+Ht94cMuF30Y8yiD7DoPRM4RGs+aumMD3LcLYYObVMYPd
a5nBDLvLvB8u1phTLxdGJ+YzeOVZfKLuHrqaAsBkiWAxTPp9syVuPSu6T69athA5O3SnoKtwe1HZ
HqsKPeRrcrLqPsKSIq1GHv2z+rjovYdUsX1ZdR0svbPH/wh03VXL10+JYyJ3ehOUy7uTqkJYO0Zl
gSW6EunZP92PWq2sZBf5CBsyf/WX0jVN9Xs/3s906y6O0Hy5ZBKMIwh1X2yJRL5PP5xsuFWh1dvZ
V4cZnvg0EzUjubwSI9dYIx2jQRbOhZDZcx+b40OX1SnlXKztVCEblTaYIkia8FCPl48pczwDpwff
8fw81iR87QlGQKMrighZoUsGmz0p866264WIrkkjWxTUJ/IR0qT9zwlcVupSQOFacEq/jRgJmyhS
gzRabzeeECbVD5to1Pr5FZ6wX/Put/bNGzkzwaITJswsGw45hR34JiS1VTu2bNfAMfHLU3p5h40p
cHb2Ainq9gmuNQZxs4AjJtifcMPC6B//kX3w8ZHkRWEetPPpxqGR1S2MHbcDUtk/WLHG28UNicoC
IDP5Rc+fhe0dpofrv8roaUzhf4ifzrSQYGIaD50FriQaXZP/PNS51SN8nD4g88xfCexu4+eRTftd
OjK9N9eBnvmKvLVKFg0xuqF1/PNXZ7UjV3j/A2RXO1qxEdm/hw1ijx7OIN8pJIutxK1MX/7sLWMr
JLiJqe9nZL8F3xTvZFs4KCWlXop+5Pnyw00eSx91H/1L0grN2GwE581FdmJpVYFh9kjMVIk7RUpZ
OrBQEeLbuTWy/GhrmmJM3vgfOwn2Te8EOce/ZD+QuLrBjij0znmbv0syr+rc1ICGKMOO5s6ocm9+
gT7Eo70j784T/uyLTXQuwC2IKKOlpG2TDIN+m/Pu/os5IxDLCKEZmI0/T3/ScJoUzxhpbb9bELaa
f5NPUZg7EUpoCjNn2GKlk236coLVAUmXLlKrhn7CYKkMuxYBIQUwO1wj/H8kJQzkBgPhxW/WfO1O
N2BAZOCuFabAYc3PFsvfkQCHCe7XrUaQ0Iubuda35EerZygC+gUACbexEzQWkaR+twraJ5mobXtn
bV84wfqMkFxUUJFjr04VceYDf003gyACJgSqDTG19W2HXMq9V+CsU0s8rgtEjiIfaX1oYyGkjqvY
Q5cAXl/A03h5JWYAFuSFTjhAA0OeHqZdN3sGZSru8rCWRK3dDtbgFALAsGsFPNxxxrA6APnbQAUE
L3rn3hjOX/aWxBOgwIkEUwW23jWPYYaHaeAJdBFv9oJyEVtHyqVxprqlrOHankFhZzAtYeIKlnB3
pfkhQopmM16pdjUCOIF2/A/G05FeUCEYkHSPkwJRKVhvHViGNs09mzaWZkHhnHJmo364wOB6ojXN
GXGSkprgZ6VS8pz+2NVSUi3f4K15rDyG6UIpiVYWrGX0ADC9WspKjgE2SPCIVK92+udDXElQz+Xd
GHP+m4j+r7pnbzTcwSi9aL8OX+pGxNsko2/TIBdNMOjDWhPeqsN2Q/CjAw2AY/hnsxb+IsA6A53G
uSDYC/F2lCr9vxfUyKRn7IdMQ5GFq4hXdg823fGHn0Yz470PaMI9LJolbbL20J4nWhaWgPqaPaB8
1V8hnRDlyINo5dAvOdENabMihHaHqySbSnU56q5ez8u4BAkQPZdjwoBoVaS2+e01cBdlGqpywP/O
EY0LS0f8Vlu0WAtkyAtCAABNKS71j9LG2pal+nWcZAzX6mzhh7dDAy/1s7m9Fdz8IPcY6JD4bgeJ
eqtRE+PeWIWYjwkL5ChLUxwxlppOhZaY8814BTZBQ5uZjjjWV8V3w8J1xvp1DogHq9sYBpwI+vl1
eYXV6LRm1VnRiw5KuxS11x5GoE9P8OYTRmOPQa+qAV7vEMRrwYEO2mZSl/bcvrvp4wW77z1HfUff
Bh5wGK5yRIiwlmPSe44yEx73K9U8TRzwqEs0bk6zeG1KUvQrt7Me4qQWqA8TICrCmrjFcGy9qONc
0w2QqdqbAs6/tsxymIpt1TQYToNFe/CPXBESKChW2+/2fmIUk9bboG9BakTdETF9NhrbOC9eDl1H
cwD/Uy0c8hAlbB93H69kiw37z2DdPkvZdcZIuq3lHvxpgNdihGP9ZnS2sTOFgKkprupE2o3k0HCk
3uzmrzKEjimiTNARhbtd4hqhOLthWcbsJXNrENqOZT2U36WpjTZ9pjA2Clb5piLHf9pXHScfi06w
EllffsPGIsdrJU+lGZhLHr61UBwkEFpMGaeB3ttwTLNjUdSCfY2gxfl1GGEdBdgpH6mit3uXkAHF
d5shBWaK8OaZ0wNfOqXIJqgw2pBV4sJeQLh1zTAvKUATFgKhrwQELIA0ON3rAkSPPduFiETdVzUU
0XckaojeOJCHF/tXjamEWKXAswyR2inNjyhEm4qeBrT2pWz8DWjWFX8ri7unDR2iQWch7LR9KnXt
boMDpfHSKCpmnhKIcbt2C5cmApkwP6xOvNRueWuchPGJQInjUfCT5anAGzIyVn9CGg8VOjEEemka
hbRikIhnEbbDbne/MBOsa3qRaCwSZvG/Zq5+XymP6HJAfV4kaRmc/v8XjCo3tm9oUHO7rBHIIhh7
prNwWuA672M6TJJQBcTRC6CzMxkY6bjzFs7c4TrX1SAnf/oZzYVhMJSTJUjgnAR+RjjqY/zU0fCh
02z4xNfTHLYiVKyaAWbRgmahxhaEi3gAdH24gV8HZh+1bEFLU/iwZImcj+xQfWMyQ7c8NGnBJeMK
M3ZhyM8wBZMiBD4EHdSZu/08OnWfKftF82B3gQTtkbDmrEiUqlznVE8ua4YRP4saks8FKVS8tFke
qU7i3DhOxzxzCvuKy25rwBhmxyTtAByRARu3RysnE2hHBSeDcb7YDwuAfYo1PfWfLXsV3iJ4D8oL
VslRsTAFYGHZfJezgjnaW5xypdwQ2M0IVyBfcLtA62QWWexty1KlvAt6ypdTBZ0txfcyYcsaSDXb
/2HTgQ52Ny+LQjuT7FUgjJhp+aLAI0IQ7pvYDew9j6+fy0ZafYco/a8x8nJ3gJ3aotqfI+csude8
zBFKbTAvZy1QJJCt5AC5R2N3s1o4yUp9gFQ6+P60idaUAaQmKt4AIhu8EngCtgTzhJcs4z02Ma0R
Vfz/Vtrhp6BO8Qw6GYMoPR27CP15L+3EyAyzfa4W0xy1A0BinGoebLgBLZeQ49Kl/2wWAfF+VUMp
M6Lf6x46z7hOi18Y3rgZB+uDdUMn5I7/6w4iZxFqJlhyjMNZlGAmK2idSlyExjRlzRj/KAfvxmuA
35AD6vksf69BHkOkAJlhGo7bGsHaSvj208KtB/FWSbDDe2h7jc8CB+nby8gGPG7A/P0J01Ks3gl8
DZjNzFcUiS/ESqo2hHvhj2F1kxstKK8/XtVYRwvySgAbMEXmTwZSfizsmA0pI9Y2OA1bnRniO6Ih
yzLOxjO7hl8jbAv73Yk5AzXQcJDfPHgHTATBt5620WWNlZ3Uu//G4w4RhryTvq2AOeZGSaK5wbtt
fKvaNlA9qGr8FlCf1gXmuMqAbePAiiAoEww5MBIcjeKMwT0G4MsQYezGOAvfDbKt/46GolCf6WfA
6SBWAUyqYg5n+x5jBUM5y4PlJBmEEvsIpYxH7sAV68hGXUAo5KDXNWitwyYXd6nDTz+TTd0tXM8R
+9nCdRzZbJ1RLWsiJQitVWy4LVkSj8D91T5r7pIDwbzA2vyZpKPBH5A/5vvMxfVQBmxo/gH8KFpl
QfIKq4gy4UmSzYeb6VYqFNGp3xkzSs8Sw3LJ8QXtxva1j8NmShH0Z9aiahMi53fcJnI6jwty/orp
pAzydL2Pz2bcgLdcJlg2KoAOY+5EYopyU3ZGQB0jWTXCHeE4El/rJxwZgSiRoG59Q8IZI3zxCbVX
+HwXLopDdrZ+xTyvFq3mgSTD3gMTTchNl7ba4cAaOrIrDohVCt+xB1pw7TTj5O1OUd9k+hMOahon
gp8c4z0UqzG0zYEcI0KJyqVVmyOoSGavWt1N6imJLCKg7XAKHXDZlIGoWt/56cGiYXwrV3f30kaA
tFELmaVRltIX7r0jQ13sfzZ9iDb51bcbWZ4kJzdK5abAme01mjjeZHMEmCUaeVkx1qNE3iz3Z6Mb
25055hppCICXMIaKGLbQ0Huzln7owddYmzhRiwlMFydQK+z0nZuw3dS17cPTxlk9GtkaDdP2CB4L
INL7N/ZHm9tEQKunl5m55zH1s08Bu2ZDIAN+n2FGzG7+LZAxwJVYVsqGRQHHk9xcVzxHODkkAPKt
zji7Tx3bumfyXKCmhcwwxx+xQQCeq2NDdUWqldYKw5c1qJkGtVxz1BLM7vIO8qO4ZokWvrxrcqlg
mDkP0xxVeVNQ+RV+o/aiyLhZhtncyfanH7/4z3NEmRitCo6uJ9tHhbXfWg0qqQOevsPg1/HBXFOv
yrbRTzPI7XJSlaSWgSZMoqp42uMVnzIxE1+5LiUHV0cxtG6eD4ENmFx+jmQLQvSm/63S0Jj+Zz1M
ghpMDWaj5oNUjapAJ8gJFBA8S5zNvad1aNw5PwY6KVsElRxe8Ab/gWCj5MWNWeDDR1QD4l/coWij
OxZMuWwbYlqinctbvRFyxEADDfB5XA+qrQP+BX7XkTCGWq4mh0jm3abl0jHx5xRCDhRjgEBzJ0qY
WNve9WHLdP5AbFZcptxCMu20o2O7jwTB7Feq+KbksMOoGUg0jSbmVDJhZ5nmrLimFzNwHVDS/QsY
7y1W0DbkHYychNImitXRQpxJ9loqwFIiLauhH7bIlQ6inv9HGH8hBimf52w2NTQnFBEdM31GVBII
jcvue7MDFOtBovMtVZn6aPq3hoWnCBUQkhBHNhye8BU14T3Zs4+pPRV2Jd8dfsuW6d+TijHnWsXI
PhkAM/sPOZrLKcMxfoddv+EkC9QfKmzt+8mXb/yBeexhSZhmj6wRH8mZd3JojvqKPkoZGL6bPvmh
kf1AP2hRlUjX8wDX6p/r4xQS04J504abV6FVY63pgN9SEdsbxmE7193Pd7IvJImrgd35zZ9V2WvY
3YcQEBQ07xtlOdDydIXuHUGcvpYrRoaA4eY2YuaaCkmRvJPIb54vvmj/y4nip4HqiPO3nuwEPzJ+
wRoJVe+LoDtsSO3lpR9ZEdMxl6stf/m6GqR0B4pIkK0kY/DqHry7ea+KvBP9lbyb0jx7mNPgtNZN
KgpbJlvv2M+S/rXtOaVsGEc6/j9pV1/YcBwf2ZMTvetPsIiib6n0XhKsPwbJ+4myMzsx3u8wEmKL
i2Ry8w/oXCXk3LmEUveKed9a6Z39mn26QxT/qTzcqoDjfQ46MvutjORPO08e6NALXMhZ935XK4tL
pyHfJOj7YQt2OZwBe0jMranhBx8pKJDepVvaSAwCVFrGADk1TiLtxVr7ECD3OsAoEKYbYRAFUiJg
HCaO+WGntzmSDkciWOsVjz54rWYZSjnFFUcD7vyS/dnONCvm3+Uo7EgapVX7DPmiTvsna10IPlox
LrWcExUCxkEd9DbXEmq5YKNapbxbatwADOQB3Jj9XChngqy0r+1O9zCxVN8bkGa9/PpO/cJiZjTl
SaOrBUBtXrz0hp2kWfq9EF690em++rgov5W612lExjNRtH+CW/pwrdSxJ270X3oPOm32h/meUj+X
wuZKj0vFvuHUjtBhTD9/osTBvj+WPXA+O7baIU4ivJRNJG6EAZ50wOb0H+kpgUa4VPewvUYdxrNg
yRN9n+UU/QI5MuC8cB2Y0vX9enwux9puCQ6rpOPd1Urvx6HkbIOjIWyBzpKnjthoJfxJnkRKT54O
MUntyHa3lAJC+z3aFlFhgp3f57XClEs55tENEudwmqIfjwHnOaVP/pr8q82OsomiSjFzxTaYkA5E
jlqQL43OTN2ALtQYdQAdP5Y7jVkEtX/cdDgaG6yvFVwUS//dW01m/cY/4EAJtl/+IF6z6dTVg94n
laUpNBdhfFzsAkjmhNAhxF8KxDGCn0ysQ7EfMNv4wSS7NMvxLO18CbMc6RYLBlATHmVzEnvS9cMf
vaC9rGl8DaStl92GKmuGPcpX5Y8dhlPDGPntM2tSXbA2q+PYKp3sMBZMpVccwg/jJBYpWwNPiv10
85cpEz8XwcWXr27rx2atJpqAhszPemTpUDiTUqhpABCqPnFlbMjMiipgMtsP02V2vNaga+zfEHOT
hf1ZqKl9qZebjmNw5C6PbFyWNHqzEPWo1kW0I0QmWSb+b8J8+y68C8s8zpMBvLVng0V/Wa4lzxCA
VHaX0+R1WOOOZYS3UbZ0K69U73uIrKj+O9PxC2916NwBShanJxd0EZmHKLR0zZAMcdKr4PFNOW7Y
i0y07sYF+YwJoB5XjmP19adjDuuFhOgc3Iq39ceY2x6vVrJLDGqmutRqxttDh644a2CHE+odakxO
9M2qKC3vYwubOMPku2Thff8BpzgrxF9KrAY0YWN8jXcp3tdUhEITUIOHecHNQhDy4m2rP2prNXnt
+M2ZPWyKEdxWLhYKd58rBqJVFuNqvHEaOJAjL5TtH5yrCn1EtGUAYOofLnPxXcanNKy83LcUGRUt
tyhXGAv7+84j3Xsla/mU3DNHCneNJYVE2/8Tlxz+zTiJjjXAEvi3wK1GAdJXh0Ip0PS9fWS3rj6q
zEeWMGT2mZ/txB2VmUQWauZtaPleoV41Vhs0YLpM7auUanInF7HZLZefujLxVu55XiXfogF48Uwh
y2GrzCXildRmLnNJvBS8emb4zq247WbADKL44sinyBhWV25opLMpwE1cnz+88pmuTHiAKqpfWgIl
bKKexBXnu4ka8PSwDUZS3+Jm5AU6E2rxfvF83aoVzMzwqmbY719v6fw290F1FBanl+9TFJK79OXr
uq5T7ZZI4Bmhn2mfOfyYF91EJUMFbNI/sUCi+15NMUhccVeGgSLhOyCBdp8aRZHE288R1hLZQ8nT
SCHfKeYyUhE/853TjfCAuDghUQTqildH0qQfgDeEg2S24iXHvFNtH4inGvqH2jynBjs217/2AiLS
sYBp0lQENuFdDik4XptQ2XMjIQRjm5hbmHwhXd1VbxRnTMXqqfzZINjn9i+STn4oHO3FxVA+JfKU
k5WiT02k0PDsP0izIIeAOxmM0Ji3RVgnIXPKQlTvy+jKox6yIjA/c123hLgTlaJkoHH5Z7+N4Ucg
UW4TlztilSuZCZhxtK5cgQ3yTlygGKO6BKgmV8q2n2TN0un3mT8qnI60ZlZRbiZI7MgQQdeQ5UFU
xbbGGh8jR2G5/PaO5pZFtn6L/VWYGVD1FF2MKe9XJrdDWpONo4QFtNHomOFZe+uuOorm0rM2QVba
egnxalb7Ue4ViZkAO0xQvE3crQsMMBk9aVmrfeRXVSaSYU/Odw6RzDphJJac3/UvJ82zqRq/DwYj
3Nx9U8QkOQCtRjjoKeX5E5OvQJhNzhi54M0bJY3TNFHnyQiqMU3UaUxrJIvBMxn2eiu/zsMU3p1Q
HYpAyYwpdrvGjizf5ec8IciHS23Od11/Mcs90JRtdGgsgaOOgE2bzhtkGRqmz4LNIcQRCkofxKzi
YCJ7giZvQBC6i27YEIWUc1vYunGC4jLIl0rqTNLgiB8KeWQ0UQ16SCKI95x7HVtUhcotEMdxDuEw
PPKEIsaHRiYmBGGyHaprW/VwmBaEZdD6jH0a/u+91tB7pWFOPZKkGxEdf+Ev6BAHN5hTDyp2Vqyp
HB2Cih8iazuaKDVEyVmt60QgIWPxGQYhSIqffRVShk2dDc1HC6vZvSMull4gaOdKRxLRN6hPLV+C
XEEIDaMXvcVzud6iWPO3h4iZGo6wx2wz14dspnc75e9/owlqHSQC0pT87ND6CQeJWnrMuurBP2NZ
JWaJDkeIpCE84JBAq2ESfpeVku8rOTQFeKSP/eMDvAyV+iUdvRY9GPsMToQvH+/itnLUIT5MgAgv
PJ0C81KlnnseCpfG1GeUGitRVWb7mT7aJ6rq28K3jxMrucHQ4+vS/m4a3LpBp6+KUE/3Kerm1Ggy
kzoFj3yyrR7fLK/ddrfQccz4JZfikH+3qtBkkj1Q5jkdHMX82h0qp40kef8nGxAHNztLqHBuUu2v
lN/VMqCo2MQF0u86m0QSLITHSsddi7UJjiiE7cPjU5Phkr0SwB20Ptr6vIoOcS4k+wi5oljfDSZZ
s1xR7sHrnFWeh8uZiZrYn4PBe/g3o8iqCGYzGmxSUuhu0TPfpyK0bfPVnlG/i8FIhe0TZfL30yCQ
89Z8/2oQCjibX0pZoNXob/HMgm5k3UkzBw8/elS8l64r/2C2MQD6a/ix+aGa9JVqa3a+yNN4gqMP
bpqNIFMMux//knBU/WL8PfEpjcmqDt7wgnpBoe4/pJ6dcfQVBREYgsC/8VowZyqZy6nbZaC7aW2L
1TVa0H3+W/N1x1ohTnYiZERWlvOtg95JXoZilXRYdTeni30gDVMMOQbBOIzqjfGo1apV7vzOTFvY
YU+l8/Z5/rkXCJSQ9B22wtVLX/wmpfU/4nipthzqTRxr+q0u5utQmFK1AyLOm9P3+FLVTHa6kXdl
vpdFz1rbs0TxqZK3dUDwNFqA1p5ay/Vtk1QbIfPGTq3F61SDb7C7IvRMl401gODfgHajB2Y/iPVH
GS3MipNBInF5WxYuJXEps/nZnsjZiDNkrXRhQzRDYUlCixwYdwl6sZL89XEyNLyXDa8mla/1E2em
ksjS4+Jm/AM/0KWI1RVCXfada93eopvEb5BILX13U9Zh6cwnsYlaaF5/gfBf572D1iXUoE+CjVU/
v9LXJ6zGAFNM+sHdLanCxzlUpSQ0nXIb4DCPlIi6NJPuGkyLl9MujHogqTwOqxquor4LVD/Jco1r
rmvyT8yiXpX3HmNE7uh3HKFB3NrZNibBcwRnbbJiKrvRqhGojycBaXAcr8uchk98YYq0t3M1qjsj
Bi/qdko3CfSCgBwgufAYGQ1fbolV2Gva1JRCl3qLTUrJMKcEh56fOuL9Leh9KMW8377f+1IltjLo
U+G7kpDMgRnAkcxqnH37aIzm/AXtpzc9LcD99d/9CKWYMTt+1GTU1rfUGZcnFPOmzTVZhWzrOshB
dDwFJNEFMDniiZq9Pxtey+nJ3wE4Aj7B+GTWfs6uRd/vhptAF6PkIF3gc59PYYpR7s/Ls+7Jfbkm
0JmAIyBBHdxulVBWECy09HleGwFGHYLrYeNivBzZkAuyDGQ+OXpE2YgcEDai6Qd3/x6msfkk7PRB
SrusmnytwsbmxVKM1bblE0M4EgA45Yfrsy5Q1SY0i8FwnGv54zXgGtBPDN1kmtqnGebt/Id84uUn
mJBZs2T/49sAQdtNc3al0NyyrF/ylTApgREF25WX1eO3Vw/EgqKIUpAux8vG9dyFljnDmZYZZ064
gb89kxDPycDBAfakMeTA2nKHqe9wBnCW9Hq4fXooOhJqGBv90dQPitKed270xI0I1ENmr4MvARP+
c6Hw9DwwAjxmJ3r5Bg+Fi6GXkvAFBIwQbMP6MOp6y6l9zHQXFA/f5ipiqsRMVP3e+TISKe5wPQD3
iNiRzW/QmFQoUtjfJW0Ge2ZHVGbs/Q42xloWSF6ssqrMl1Vl8w2DvoozfvmMdLhBCV2///7LBDIe
7S/L4HcaweHe9KpCmq8PbLjlObUPi9h5bGzI98MjYBR2r5M2rzOqcoWPKcI128g0dE+f5en6DKbO
fJKmDornYuhFhED9WpnnloOwla+By3Leh8InV7w+W6DauegNa6VGtAoKn8NCi2EjsDJz8ZP17GhB
/F7C3WrAAuSP6ehXJYDuvM2cP1s3iSvEi+SXGsg0SGVKaSfYMGqJw0/3G3lzHvY3qqEexurjzysk
UAsuPGTl1sh/X5kSbpQeekIzcJbenoXDriZ4/lcsFvWHcnjVgaRPTbBFRV6/BHmSkE9T9vWV3EqZ
HOlXSNyViX0KG+GcN9bRDNweBDIOYbPOAWaaiSuUxFomO+u4GeuQbVaEIE4XD0LxfXqR4yminHGJ
N7yECcLvCmfEvpMTcEfyGth8t02NHQrz/WGn6bdWbxx7R7/AysHTt2DQw5yu4p7VV5tXO/dzCnP3
gI4PNe7jXIOda531WOSTOsKqeYHK1tlTdELyt4p13xt6uMhe5NbiROiFTqlWw2VuHyUZef2PSd/H
4KZWlw9sFVy0cZtSRV6ltE0mVgJ5DOdc4qJrjb/Ab+0d9Wybsk2afc+gvVjL5sW2P7QMbALDi4K7
P/vMsuzgjAK4A1Je6+5BBqxO7CKbyz6DEk6aQWR3xPQCrQSGNUHkR5KQJ5HNMdv7NmE4ee/dgfFP
g4Iz/lQOHZBi/B5wHE0GfPLyC6XyjdfuDY6RVaMlx3M8/cISpZoVPQ7c1y6Qx16hSCwg08+QV0WK
JFeQl9JntC1Jq4/gwW2BcnGkyfLmrcXNbu6xf8oTyfqTMxsIKWElnCPbtInY7Ta0AaJN0cTv4ZJT
qrzOe2flk7kItOXz07lnU9G0UrDHJTpvgcVwUdcpgBpJCweszXmTV75ajDQAPfKbatSb/ju/tt8q
x6QUlVt+bWM2JdBtin5KbSfyHuoPgNv1+aPEm5UL9Oi1TKdSvBTSHQGFn9/zcfXPCBzXPwktZsjf
Ys2k0Mt8AY/wGN75wWeelFzHsEA8hv8UyD8CU4GAFK6QVJxN/brm7Wl2gcfjBByE6ZDVP40dsCfV
Lf7ppxhrC1sZMRRi6cLa8yzyPjBp84ezrfaawHp50RRxLEpOH792h6oKcm5N8twCOT1izMNvqxyt
cAWan2WAvnwXWYVtqAKOQ2clP9h5XlPXMvvSnIKhV3xOfntDHDBxWBjoypUhd9dPoFHaOmLYB81N
oAD9C6nKpu4aFEgJu3/rH7KF1Sbcahhjgc8JiRLrIvdRMZAkI8wsYM1U0oeDwnCahQo1kNPLiMaM
/4GnDzFq/L2Iw1ioSVNfopTYIVyLsThFK5Z22+7jkQhtvKDRwPk9cgdmWOvVZ9jvAY5iQdx/APDS
05vsSRbOBTw4jx1unNX0QXsgEZUl01b94kJTTZ1LlN3y80E3rSE1brSEIQ/xPs3Ucp9UDo81QSM0
D19xzdmMB3ntclEdoJETF3x5eqKXS2l05EW4HFa0dKHfr/1Rx6Uog8plUUd8krajLb1qMmgIoe1r
Bta+lpMUYqnPINoQqdCcIBvYCsJ/jD59XfBEuQN0MTRRRs/YHeD6qloaYPqYqDtZYna+rRVwLAj/
kHh39JzPjpckIWJ7F2E2u16BKXNeMmsL4pcqPl2LIkhjMkxdk0Y4uESxAqWYjfxpa2hwfewqDM05
PAtF2mbkqPc14au3gZRJR4xSqHOutZb3st1vzZedG0yv8yGyUm9tUPyAd4Ept/vR3MoVxSq6skO5
z0gxI+Zi8KkG1eF+Dmd6KvYsk/COHzj8TuOC2Q2F1BbIq4Q9bTG11hDFqXULkdtVaCQ/YYqg9bq7
1S08rk6AllBmkMAOsRznfCuS1JoSZXaUgy/Udqk73/a+A/xuvxtnAJXhqT+qpJa//icp8p2V7RMP
u1DgMrYvDZSaF8I6aZ6c9osx7pnQd68MI3aRqE34D0pkmyl4xBF4hi/XaqAf4dt04/SsUQiVh4eZ
3HW9SGS8L1+SPZsKGA/5nxpBbyqFbAuaZKVGO6/0JVbnNGw2+uVBKMTinj4kaRhKCy5PQd+ZN37/
S6+mOdTEDMwXeYKY595uuU8x0iZQ25QEkVFPzIU4IYia9Nm/d/butJIVwVN2g8lRYN7F0FQTUixQ
M7SjtOPCir61ZQrw5a+8D999GNqIiN/icJlIbdaAsPSYKVK/I3NCS1lq8LBjZZiWDSz4Ctueawwg
3aHOadsH2W+161vtmC8um9Ud8bd0UqFK8j71y3dwE+x/H9K3DiBuu96YjMOR2YYEi0W8B8vIDul+
d3b1CzZiPuxSnRfBKa4UV3C5/AaMtt/loeoihDzpIrH+S8LgiRTjShHCLjXB8V9nHcb/m9lJdPvw
REzRiZDiezAhpB5yb5O9sxgVY7tOwvV3bNPp5SiAslte74moUhLTsR+lCjbQIHD8PPHW23jCfHUW
RHz2SNnt4Rk0pUe96u9INC3sEBwmfc/6XicCezeRMeOenJ1KaJW3qJbcxGlyml1rfkJPEevrd9b6
L3uLvo/0h1uFfnBaWiyGGgoe8AJiClTPcQW0e2M8c7/zl0N9iGOTDM+CtzqZqFEcSd0FWM6N+/XZ
9ucb7D0SArbgiOAsD42lreUhjX1XVn/VEUpmIcBXwmAQf9ZQgqSsp5jEqA29UkaO+5XhcsvaOPYU
fXT26f/2PyJEGnoifIg7BSH43jmM7CZRUTEG34zsIB6jik6L3A7XpvquzyXW6atld27x3z58G1BN
+ESlV0cKny7akHYIH22MGOS0LpxRALg0jFw/GWnVw+ZXPH76DBcSzCTAxtXxUQtQBRIUzUU81QGH
V1DnNtLgCyHx5U86nR/MMOFXBta1TLpH4qLh7MWRJGzQpcwV7yUhFdOonHmBIAdzZBJzX7wvm22Q
adC81WHi5SeDaUNdmGERgBnlZoqwYK4dwM2ydmBZX6/CfikldFpxDqN7y82nC7V8czoXLDLzVA+r
4Px7EVHe2YxoKhHuNV1QAjnk47HAgi3kkoVk/XeT9XTkiPlk1vvMpNO3ZMu5VDG9dT0SXCWhOLK2
Tcd35U0HbvK/qugp/EbV/KMxl/9+j5ar9C+ic7/M8pioutGZhmZQTuQgQhY7PU8brWmQjEcDZzP6
kG/47/WLiflUEHFXxb2eAj/NWk9ddeZlzUQsz/nGHmaEUWX8daeqV/KdcYM+q57pnTE6m3F2O67h
bN0dGKs+gt4BhG/PLRZaCvOk+iS5Rea3g0ltM94uOPFRDZ8ngWxng3F/iuEAe9Hw8g8y20qzwlBs
iTgcxvs5bzJeFFUNipTuOBOdR0Q8wKN9zG3r+o1OewboYwwhn82C1ta8nACfSifO8FeUFy/BK2dc
GYrKmDteyQtZ4L3rh3piuB2n7+Xi73YvAFKE0VN3QXEbD7NzkazkgSBtnpROX/9YuD06vzZs3Sog
4jXm36S55IgAdh7A0B7Z5F6RezaQPwj3BkNuyDoX5qLvfZ1HTyZgqb/aaunCZFifd0+bo2VedNwN
ihXdp2lagpsBsxPG3Lb9VoWz7ZMFyrA0ysY3/pKbjawCSBaxFPAgiZ0xDRGogZbq3OpT8uv6+h8V
BeUdHcb7LkCpHyQTyXPn3eAOEUv8SvVAx8C/uY9BX3x5IJyR2ozANBwFoIFJAu5sRHnFWtnLIr5O
S2T14Xw9Fja0diNmOKil16x+dnqZWf81ZGQuRgk6syqL7qA7TvJYwANZ9i49R+/5OkToMlraD/MQ
RHHbD2iK+DEeCkbSe139HWmwzxkhveaGEQ34jp+lh1/XKwo9E/PMMmqm055PZKWUSyxvI9HoQXmx
kp9eQz0yu/FRmS5cMd85x7+ca+SCeFDLnsL0QSGz8fVz8pSUgd+W0LwCs24OfeC9N1SnBycKOkSC
6k0SAEd2O95qTjM6pZ78KqZhkBth510RA9Q0WBlChJNgNicIGVnBmvf8awQODfF9vs96WL2UmG43
ebdzuxF45kHwwcBM5/wlvjj3C/mTdPoSgxB+eXCHAYxbCUM8KEV2MElLj9EUxj/mLM1aIlMfeo0z
kXxlQaggfigrolwCLkzIrMwsK8rSvpDDPYqiS9K5WBVDRNv0AdyFI6TNDhagxuXIUPJe2S6djiWd
SJoBWKZ7BZ7KetRPxhglzzETZxgwl+aHwP2BA1W1cEG/KE8h/Rbz7uO+LMJxb/EBYIfO/fLqeD2E
qEd/02zBcgBs/eb+0pA5J2VuGYTXcqI/fkVSnuuwFyPtsyryVozaR7faeMVaUN/SucHP9YDurQ9r
pS9z0xvobnKVcx9pT1TcE4fd1AL2IC0rsnkeE+J48Dfts5YR1C6Otg6fId+LeSCRMSv61/Ic08UQ
33uvhtXHDoMB4QWH9ZYe/yBkaJNvpB+1OdHJVml4ERH4OhGo/ZPSZhfAerq2ZFf0zvFgnDhyLbh/
EQIRrjJdbyE8gnBnPurAO5AVn47qs+dXyoguVw7mgLF7ZZNvRDt6QrHXMM3LDc2x85Ec9nIeT8zH
+3qJisKy5UD4J4KiFSZEJa2D4cB4JRcveZaz8fcDKICUEboS5Ed4v5j7bgm1swCWXhezSc8Pi3tF
q1oQhmSPalAYLNV+2Zk59F709V80j3P+ebNrtlTyj6gdbt/qoe60sC/uZGjVdsoYcCCwNLDA2+E4
fpG1AWTEyQ9r4HBaFgoNDr6RX2Vs0+OBWucpSYig081u0uqNYyZMtaEz9ps4yRBaCBjdZ17VtRhp
8y0UVlRArAq3J/VOzIfUFfTltLMxjVagUebxmYgBH2U/wGUv+C5rYGVtRBJJR3jZZya/EOU8c2Yp
FvDCvr6sKFW+L0wFbfvsRTOnz06ccvckfVrEJizbCBZaW29Dx/kcTxOUEPCrE1jMbBjy/Sq5KHN1
K20grZUz5QJAef9kPVDxGvhsxSyWsNnvQ9l8q/IktrmdcLJkXehqQqcmwf4j5HI5hK7fsbM4x8N3
zORf6EHWyPkUvxKAWjH6BgaY6JX4Fced4F9QI0y0UxBBUIjp+w5/yEJ6qjReEJ46g3Y0uDwK2UhM
xXAIvE1u3OH1uScpD8ND96aJ4HwJHcvLNpbdpA03pd+SSzkm4em3pTv1ltYNCg0nU1rLuZgWUc3l
cGaEmJ8n1aXCkSGHeu3aRkDYrjLpen2xwVwcFXhjE8aStep5zM9uMfRtI6XZiq+PsDjMiQuF8g3C
Za+yympJpLavUVKW8gPWJc/q7HPhMyBEXvIQ5lkyz73r87wiu77v1L06LfvIlIcND7E8deb5NnXg
ZvMGsGqcAVceCFQkEe80k5JcsUONQmJBbAMdMBrL3ZIHgMvZxgpooI9yHFApqPHrTbasd4n7OjGG
BQPYidap6T6SxClYDk/yp0Sgk4Zj8TVoz7Ukmws/hQYKKEUZcoHwGo6PWoZAc7fp7CmhI86idhcr
LPTJlyAUctbtYSvr9/m35IGveYNzElFcG7jZD/hdA7Ro9Oogcq+Xa2mRFDwq2lCx+X42h1eqewgh
aN7ulmsAudFza1Qx6iWZGSvsgK8RC94GxG4GO+Te11y9VSp9xa06Gv6MIV/HZVXQF2grxt6iO9ee
P409DJezXMa+3HTRbq/k0aF2r/URuL7ZLI4W2bzRF9nWVDP6FdXAn+m+SkafuwFU8mpoAAWq276c
mRdFqdSP1TZ0TyYBv7lj0CLx4uHL+HNDXNVxxJUN6FIF3AruI8is3dyZ+zI7D3r3rSfc7b16Om6S
KC+YZ9FYWlyFrSCZ7Rmc0/8CVGi/SMlOWLe1U8a5YoJGLhDpB/mSXnf8rmhTKzvW6mZmkmACTsKk
UaOv7D3fbbIDagjnIw9NtovYt3iCYVS9S6ZJahw654SpPzxv0QHC12P5tv+R1JlnojPDhOg5emRp
ZqSjEjccxuDpRoGZ5UJXwp08A2hNWG6b7W5ebpeFHezj8pxosM3cobuKGygsyt+XuNNqZwI76WwV
9PTlQRsitkjpwFtOEKo5xceUTIbHAAebKsXyoz1EZRkeHS2T7t95KSuBDWECoGcbBnBNyK6B/zWH
/xaA5X8NdFG0a7MIyLrtY89eNSQyj3Zc3/tBPeEcNF/XcNoz8ClkzpHkrRy5ZI7cX/1GJsIgmtt+
0OeZ66S6LGMjSieRNvd2gPdPKQ4Hpna6wh3Ow6pm9G4g+T8PO0sdnUxfyrWcq9lQitYzEDpW9NWd
IR2DL2sx3nfGdgOcsPAo+lqXmH5wwqUDF2RJUTjGZu4pe+mjlauedl6OMXuUn2CJaZQRDp1RrPD/
bEI3CLV1yt/rJOHbfGLJpYTvpd2RZTzxKrn7nFrvRnoXvddr/i76iCBuikke1EI/46OvSwu67Exp
mfxnMScqHvc1i0T6pdpjRRnpMBej9/CUxsGIxY/7zilPHvqsJ20bijnHp41yz6PKd0193lzwUKFS
JgRp0MM0St4gSxev83KTW/RYzDsHCC9d8vmv7Jl4E8zRzjXOlAp8iaCQw9Gq2i2YrcQU7SfgZRnC
1adQMeY9IX4A9h2gPGD1VRT/7j8LfL2TFVGBLQCt3pewcWPw5WQqaLrPMWwtSyCNCtBllijO4EBU
14B4GQzTP6pNJLEwuueQuvZQ2JmdLdubpXtywEBvjNJy+xNh8eKxt4Roda/iiiu2HeGxu4tUQZDZ
H2aUlCgb7DDeTkXq3m6bTRIy1mbqw8yqu9OFjwLvcQ6S3//ND/ng34Q/DbjhNZBGGqOWA3x0sKfJ
xQw5P1GZwNPNYD9Yx4CEfp3u+QD6p91qJA+9A6YhhGk7dLkIlQ+YQb8Tmlbv8ChYuSSkjo0cIAvN
yefRGvay/yVPxqdGiUqfLWZBUsP7MTf3RJq0+JEhPEvUpTwt/JviFJyzs2md54hN3GwF0Wu+usSQ
OD8Sivd1OkfAixwVgq4XDWpu4q8kdgTOrwvPllftbjQ6mhvsPKfoXX3aa3yNvEpnJjdXqv9BX3ld
t4uxYZnmeo0DkMI077oOPCCDHYMjcg+bfe6+qXlsdS7lCTO60jmikX9OjpaA0KkT24rP286uq2uy
MVebD+7LbjKMgEhCSzbryQLjsMtNWe6UiOWOFfFOJBJukaZnn1+CM4H9OASovBi0LjjwfP5pswu+
tGLQ5ZGoKc6Kz5rJBZgdHZa5WUm9qt5PQeACUMxyRJXk58iaIuWgYGo4hPxaQZgKTJqZepYi0tJl
2nE4hOHWxVRkboz9U4DenzUjzhW3/f92FLZS3m9oNiDoV9snRAFj6hxjlfh5tSo3C3oAGuJJoVx/
qoFMGC3tUW1f7tPsEhftuNwd6kG/buaj43Ub7fF9yfHucXo0VIzV1k7BcC4F3aXcMCsyaWc8l8+D
t/ETpAUnKLSt5z0T8/Cbz+OQUotKhxbbORxJB7/n1sh/TXPMu/rjdJb28HxkuwUJcNScuLbnvuu8
KBfc1gaO7vP4g2EkkUUSrS3w0f3HKg++0rNE1I+TD+TXwUn31SsAs+VFthGWG/ZzSUbaTrpkcMkZ
J9EyefWo/SzFIw58WCdrGPSyeqiYvNOc6UeznRz2E2EauHgTnk/D4tHuWJ1DTn6dyNlSMlgjAM2j
kZzUnpv9SxMGcENOuuEnqah/uCxKiIljPXeFudms64MjkB/flVUHLhZkcHOV1mJ4BSAv86YfYU2C
KMElavU1KRIvrPQ+GPxoWE8Nenwmc5DaXPCyY4oi7wbwSJ0E5E4BsBdIu/KmKK4NQ9WdN3jQJyLd
fl4AzArr/jbH/TwwFqvUroI55FDYWlsgGh9U6LmVLX9hPubcjTZZwznjqn/EED5ewLWP1HyHnoNd
vWFycgGnAw7J4Gqj6d1+uhoMvhJ6c89d7n5rS49lIWRq7z2TZ6YW9di8gw39pZrr0/yH/OL8vFcT
YJX3FYK1F4aqedlxkrlrsjorJYBbfXnL31mGY6daQu9D61XoNK/iHJaL6qMTmFVhO1+vYF31W9ul
qELXFc00KOXdMdsiFrySoSW95o5Hl/4Rut9s7zQQLhXleKcfI+hugwZ3UCZJmeMdcsl7GHywbLOg
qXjAUwqGo9Cg9iyqPMhL8P55bqXuPqR6AcMP5hxL/XW2EKYKGfh2nLbk/AKLydPxGmpF6tTdlWfN
zMz7ndVRhxgek88RXcrs+oYhqNmovO+d6ZWyz/Ewghyt4XEVZQgd3fUh31+G15YOlJ5fos4/1t80
WDBTopVf2XEBcXNyFkJ05hwP7nLC6D7vlULYHaZXDiEhpY4vGaqudmES3W4Fv+2b5nVSHO0onoAX
wowWGtyaGGL9iEryCWWTejhCZPN6aWqgMZ7tUrcl3llImecBZcIUMfbUraxuW3ZiUFk5hKj4il8A
Jatk76V3YgGx3UJgKz8g4tPSm7jAvNJgyG00Ze8ERz747M4YxMaDzx/DLoj7+0eWkwdj70N3tBFI
znEIbPyDYpY2g6uXwsj2iQzP2IAZ6+LnOkfFjz11eMBnV8RSdfXab1Gv6Shy8j9Ivw+HE14e7PN1
65sHVhOfDz+c2w77jcqw3Fk74fwJdfKUYeE3MAFo7uGD7urzUgIYfa/Aa9FOn3T1EHVuU+ZC2Ier
+RHf5QjPzsprN5UbLZM9gXJe77ELRY+dnE++qgvae4tzKDRaoa4dZ/cEMuIZCS4ZXSQG/o8j0kUI
VQ5DVW0mmIpWww/G3NZJJu2fuawANtWrXzGiGavDqprRVE2QG/2MjIE7Nxo9y0vnUxFRIzA5yt+D
h5mTY/PLHN6PeCRxrkknaNhnncleaPC+oNG1H9+QjEPC84AOhkeaMKykXUxurGu6MLnlxaTO2itu
v4nwUamMSAvijhDeC6oLfuqzClVz632mtbGzzWw2XoWdMABSLMAqWUrCrOcWysj4o44L8vEayR55
QMSbuh2VMbRLkY2V0LEk5uoiq65/VYyaz0rKOHcvoRS3c2GWo3EbDPWJKUXt/vdoyE51vhOf/zNn
VibcwPJGbx0mOCguQvSbC0ZwERpcpaC7JsJmiJnFGhdJrSdUFjpby0VdT1z+p5GW3Xn865tS/G5k
mfDu7r1ab/tXyxGKYQla9efrmoYIa/G3GPnA1fY4YGH1FW3DN4jVanOYpk8Q25eJYCKS8bzXeJen
Ilw1ScWpwfrm0CO3gJ2wg+snzI+Di/j9r8fl52dICid4ISF+JaDbwMnBfi9BhwgJsZr7dSa8Q2JQ
jQaIx2XC7+LP3AaMqrQySLAUIy1tRK3CHbUAYLYmBCi6gQFbLmTF4Mhu3vVk1f5qdzFJNk4eeY6i
jE+nhdetFFP7bKjYSrUdJgkEhS9G1vjTFh8KDwVSF1yk+UVtKvqfJdpxbUNUU6iHubwsXlgDX/0W
YN6pLqZZ+1pqB77Kjgzj7A/C7QiOwYk92L7ZBqqQEOv/mRP3dhkMFqb/PUtTOg1WAWvvBTpNT0JP
gIubgV6nJI5D4QbJ0lAO+b82ZJJiCnAhkPEPMOSDfCjGaBeK9WOEsT7qPH0QRYtYm76Nf8x2nzhO
j9tr5R9LJuFfBTpPHBnYC4zYnfNjFz8DHRzl6gf/PQjNmxyYRIRyMwM9+WUshvE+YbUbRog3G/pl
Z7hzi+X+uSUyoCLSiVruDbwH1xlGCa/z960BlbguMrf7OHtfQWJr7oGFTLyXvWN6mQO7c8QlDX1m
7ss0eHIYfhH5QdvgN0ScLGBbulBe7nGf3j1Saac5xB+BFFPILVPgJAF4zef3AlcbeoGMqhkS1s4Q
ARyYTzpa9Lbp6uKAesxjWHi3YDVW0Ms0lOASVWbfdqQR1jFL7ESAZtuAUn/bKDddr3tZFmuQWjLd
9zsRtfzo2ytWizBP43YMXz1L4ZODKp7CBd1X+KgUATEF9JcuJTtt3mBXUfSmHvMKZoE/CiO7A0fJ
DvuCWgv8WIW2uasjqQVp9rdfRhxPF4klQP4a/sJAQKOYsKjsmWZ4UH5Lt02La/ouA3aB3jdGMgTG
mVl4AkMp8kBncdAWnJiBQSa2NKau94/xwpXW3T+MJTHQz0L6RbMcPh3AIlQsQ9VcYItIROhn8btG
Ir0N8aJk+Qs95WbGxkkVmz+qbUU0uSx4SIevbTH4PS5zQfim6KsJ4pR8dDumQYp1BkLfkF29BXxs
JWyS+DjVsrJrbEXgoHRhLxNi4YdFUarJ0oN6A+LxURY2lIO0k6J6yoAo+YcEqtdyrIwWEbfAFXFD
VlKV4oUVfrMq4uoUru3QttyKBpAX68wBEaaOZpYQXk0XIJcJL3zvpTMBgrzR45tjHGiO4p3+wDRM
GKa/GhD1JobsE1o56Q+ENJTH3ogDwjixKKE6rKHUkXzv7NBO3D9OC68gCVcUalG6oaqiNS6KS/hQ
aZnLUvVG3Fmh6RClmCCiPZTGCBFJ33JGXKeQm1rix0p7p5M6aQwuRhMHfN3kNEeQxwSLRSK70MiJ
4MTr2vFOhIDWbfAyx539E6ioKCSfEfss74F85IaJhpb1F/dDJLfwVSn+MJWweoKrGAviH1zH0twa
ge8jEvDqDWpfq8FNHk5Ae4w6o+1xe95z4xjdvRTsALyiBjEta6lHbQnlcVcgWJpEHoLDDpKV+6eh
xm4fXTwabt+CS9sfdIfT98la/VE7vOvOkItcyHZZStvRYfO/PbgfzLXLUUf2iHm/oZLoh4PpfPZG
7ZynepOviPthwBRrwfad/uHEJATbpFdK01o3JJHVVF5TNE6Y6rVVkgs9GAaT+7DQYGqe9gK8Pcgk
9inYu7DaT83+nGBFuKl1thgiOSqlsQM8Lz+9cqsNm8qN8AoOQEyui/66mfaWZFApnTaFOpW38AFw
F7MprglCvxDmUrtVF95k8C9gjQjZcEySN/D5XPnlwvT9NDOIyM5LLN8iXXlCQ0PVTPK5XBbVxsRE
lpIFNkVvlsrggP4vPn22+Ipe7RFokgc0m/1jTqEQKxZlpOhE1kWHhgiKEHmP/6LP7YKo3gHm/h/M
wTe4N8IwBDDbtv5zwc/RCNyAIoJxIc6mnpw1hTkfWfI+Njbzt0QH0mIdzKpWM5sP31Q68Dyk5GaM
aMe+JYMXJwFHmBX2bvFBQsxkTPUGHIIxg9LxU7s3bGH4ouYN2/z2eCy65ggR3J3VPTuIewssIIub
UCrEQKQoQOD+b9Ca+mi5WtMH9aGwOzI4GWvCVGJahXrVpp1g4mDYvVoUNGKuWFBkgf5qmPiMN7kp
s3Hmmd5p4B15dFYndIZLU6GubjkvaKef42SHOp2PZfE/QY08EeJ5FoDnjrZOVI0V3TWk9nPAzioA
o/9iyjBOJaU67HxbXBZBRUfVQnBbwf16TI+AibttiPJZWVbYsEmb7g+jPkB9AFZa3st7PLPPFDdH
g8BVid7PecnymOW0wpGkEUKmZGMZOpBr+lQOBC3ow/mawTtTdKmpI7xYh3Eee09uXNo+JkFek2zC
LLHBieoxeNEUGRYeuNa57Py9NXhMvq0O+0rgc4XcHPwO1sTu/B5qKdFNwEtb9dtowDFRhm/FR+BL
1wEzdVomvo+j5XIuXI+UupUmtlo5e2FYReIxpH3n9t+OK/avAahXHPFBkEEJIMaHPTnaqQ/N+hV+
ICfJ6KjIBlByotqdK09Q5kxdobfUV/3my/dsZftI0BZRPsLeKvkWT73j4CN8uYhuqb4Knx2neMIY
D4VRFC80hgqYfXfNJUrNzdXABb10kd+jLxujD2gSVOaYDTS6grjWTjcdqgoAp92jeupKacDn7IRA
rAFJJVTj5xr5yhoytdDlrMNEi2w7LcTYji+OaJ84FLa0zsCuGhIQ4I138Wf1HSQH4752I8+o2NbL
a2PW8c0SEPkHEArq5mB0/yr5etRSqtOQD98dy+o5DR14d1GNgcPD7FM/06hp1pp8LTZCEXqjqTaR
o1YWa8V1ki9vcCp27yqw/rDBEfbnpT1HeVBWmrDzSHDJU1vNqaNY3ctvnMu7RwxWerjsDd/tzM8G
oOkoX6oyIrvSHo06MO546VjApt4gA5BJYyJj7YKg3dsTDm4KI6ZLR4xsvvHhAiAVsD1vEKoQasRo
nsnjgpZHJlA/zIisXSKRaJdcIxi99zzdCnqA05W/RiV1DSf8eM6+8XjAarospShv0dnqLHezr9xa
hc3IintYe1X51wyHgDvjwvRsPfTqZfeFdFZddkwqGHmrl+XCmFXQ8Of0PgQnb2YI8rJ1RhIFDGCa
ZaCAIQecZQ0tFmCiMXHlg623wB83DiEZiXfqVCk1DXIWEsUSOSLhbtH30meTxctw3FJw0ltZ8EEo
onDNKd8g9UDRqOPhzdwgD18r91N84lN2nARw2BqPvDHDFO2p9cOIVBiAK3e7ZspoISELmLRSAFMh
u4WO1/zSgPFf2IzJGqXUJvMoMW2MJRzQTb/eO9Ww8vu1E5rkUAPZm6YuohMC6pSLE1JDAopYhmNW
1a6VbrDz940ed1ktcwEIOYYkHYFIAWQTRQYwNclNmdaGmjzdzfRs5r3i65mCmgbIcY2g3n7iTi66
9tl+LrcojVqcYE18iIiVhiueIZOEglogEufAtK4MlYuOiOW9cuXYe8E9d1LI0xZFk2vD+685xnZk
nNchV4CA3sksHagsVNMDT+soCDG0ijNYVKi3U5r7P3soklZN3Refk0Hto7CQfTIgOPCfZtt2lZM8
UcL0DureGrbufAk+1dflDAuzFlGD8cX4rijkasHxA+nTpwVqW8HsZMRCtwAthKBQEhZo9noptK9i
GPpt5P7wgfcI5wOVL4Cgn3gj092sFiwFNckzCRi5dinwU1DgEHP9X2E1V7wOkMkJxxD/NodXFwRt
A/VLxkvwSRF0TR3BSO0IbMzsh9V8H7XnOW3A5Hu3goBe66g9Jm/91Yskz7K/dsJamNPEeEtbH8HG
X4/oHla28rTfwAJeD/WJfkDs1yZQA1I/fsnZ0NVCTSQ57j7E1NR2+gF4o2XQH72U6lFcrNXtQZ6x
uxQ9ndY3cG2QsKDF3d5iNWcdcM9EsCPQqED9K9AzSFgAPl1TjdE+3eZ0bR1yijGF6XUVmNKiYTtD
Waf0bMy/3IIzG4GS5JeksmS7gkqBPni4IvYInqLA94B+3K2JujenZEwoyxV4nZxBernItXYurHtE
De7g/dTgDIZ6vbzM+F6F+GpoTKXsE/mEC5CI6FB8AbgUl97mkXXNngSc85i3VzkVXiJ/Yli9AlMy
wQKrQmN7+yQ2Sarw3b/so9QsUeLMMFHfrzgAxKyweTSK4wMaf1DiwIpFo2DPurkF+CmNVCeqK/Og
x4qMiQYV1M43t7P3HRBi+JYVnmGj+Y/3vLgFeD/w+1U2h37GxWOgd001PgBFEE1PV7UsyveIdq+k
nDlioP/lylvoEsIL3LGHWHAMnt18DvxYUbYzYcpXbxbxZdnmTIIW56bZE+Vr8fJxdWbqmAuiDbez
6/oukYCcjf49A0OyRqrfmDGpy2jDdJ4mcoyeVsvEPziIkULpao8n8uLp4VheONYlCdud+DLlrkgq
j2+BvxBbnvH9yndyp8nFOC6pRSkNQc0GHz7WWxMTbUY+IuOD34Um8HZM+zon4IEo46HK5LreTlU5
43fQ5hzvQL2Tglr38f90fmr4JOolCHjt6vFLldluBfcuWbwX1ZAdMtOYVNDtUfYAzYLfM2oi6txl
fgS707WtbJ3NtvLPUoeqSqVHrPVmfB08eriHC0FK+VTn40WR7MD/QdQlI8AebONDT56Ziw0CT2Px
txoAZMNFDRzP4jol+NFB9pNXvtWWpKius2vPg4u3zJH+pxBv2Gsnr7PhEUQs+fa91zTIfjI/LeCJ
9tI3wBK8+i+D444I0KEB25atAxrx5eh00jJAcPdXL3mvQDEI9JyXqUafsIEVEnAULzvxvID/k8XN
qsEY8n9LtM1JOmx9g9Wu3g0MjnWh8fpeDEoDMjWp3ie+igwbFiNPpYF7xDODl+p6lT//NTBPdZ3o
Wg4142f1/mA0iHLsWQIovy7R2PNtV7ykT63v00rUO+aHOSORA6OxI0vE595GjxXWkhbWVFfMr8so
lFUsLUS4eZElvRi2Vre7HR/GMrG6eqe/CZgDm5DjMqSXrhbMxKMSUII0GC3oH/Fe31YVLhvqUitU
B/GgxJ3JX9El3GuoJQWanA5KnCNNdD6WyIHvXlhnD35FuEFXf6I/VB2ovn7zpN2EXQuoevRDxui5
BfVSebHrQW23OYr2UuOB4l8BOxWai54GSNO9+NPpdXDhBohpSUQyNQ1PBJ6ta0ZESvuSb2w3cAnz
vAbNnRsFmofL+JD3F/2QdvIk7OMLVBPIYwQTeOod8GGVj1F+KqTblwdDmF2Tty5os+SirEe08jPf
W1vIJ+q33KomSdamgC/9vmQrPnDGG6+i4YmkDPDS9nMntC0Jb7yS3+UmHzpr6K0Hz0CzwiWWsHAv
ENR828IZzKZcsB/WDdjJupwO2Y7h/ZyusuEahAta5Vasn+7LVXl6JwxEFvjAlD91aNUEnaunZ3u0
0z92D5CkKUgrqg1ZDuRiE+KH/YyXLAHQ/Bg3+vx3rmhVVDh8NrBfsGWez8RR5blyi1EuKGu3S5W3
g3eel61NC27FpcXK7Q0ltKVzU9uynNPDlmUscYPjg26pbnb3vyTkdGI+ljvSMY/OrCw2RkJbc9ZF
/CTavr+URhOB/hY/M0pMnf6zvfvfLK50gkkwGCQQcq2lHV2c2Du2xFPhnzGjnboaeQ03lCXGb5xn
VpMdNE58IqeVRUFA/Ib/eyf/0q3Bcqe3+eySGiHyDQCwOvgOZeVwyzUKqnPkei5zTNQX8kPuyVOW
Wm7Nh+89N1xqKJWs2LeGvDInETD7mh2ldFBmxeZCEIixjqJxxW9CI1QFsTszreuonF/FxsD+YU/d
kBOztPn3SgJOWbl+LLcGFYc+kqFqAxTWQ52h3subdVkKAvCp6hahncGBAiVsMaLK/m/nVgtN50Ya
MO8wxpFxiT5bP/kIle4KyynajC2+gcWFnR3snTB+J5q5SxEKcdc8os1Lbu5AdSn5V9BItP44zgo1
9psELWXOMtBvUr7kKiWZUC6FZAOQ2UvYzdzyrBeVFkH52ZgzBpvSBjfD7EZUFHBbcKxxZIpFP2gK
sdPReNUNK6s332/YQt7So5qCOl3RoHS3HjD9NNt/AG8CYbhZSZKlnU+2KwANqZK0K9cAndoDSb3D
6nvgOyVIID2jcF0hwKKnOSrxUDl5l025h8uU5DmJT+5zpTRCqse4P2hIbuOFrUjqd2+24hj0T1FE
p5Lobryc6kcsLrKhQixm4rfvjprOe4gf+XTNeK+m40DjpeMjARqgG3yaqtgrpHZzZwwWPMnhXFuH
2UVsHV5I2+9yG4x9Gt8Vh9BbFp2XpeWvqjRISmtp7p5deTNBNWMiZwa6eFr92FoO4KaC1e+eD9CV
MERNowV6FIAYj0wkVoKwcoIwqLKVLh/LOtspSI13XeiRDPcAP2Nh6H+d3HksFwJ0JQwxdx4cyUUm
nAAAtKC2bmp8DIpDgWHtO8vXTYQLwFYkoFcTHO3KARkJRcTi0v9Nqq9ZQ3s40vGZ24k+MxBBGs0L
Vh1hm8ZKP74xgb2DPBCI5D0vJhspui+qaufbql4DrrmFI8bXIdlikTK9TzZc/tHtj3gBxYnGuAIJ
NZNqaHBFnAwkJKV02nPRgAKUHcqdZvegFLhVGJhjAlcXNNeJQjvyxfagpdjQubatJI32nK9A5rZG
lshh40/FwigkATLeZBwH/YsDlUJGUG2jWWPjDLor3XMqnuPpC5LldFnp5Ub4EqKqASRBPYTP/qga
/AF+8D3gfkSZWwzEAwMm76BztBmdALkHsOWLuGs8rJ1uWFlsHVw3xrny+kcl0dU2ucdX2dqs3HHA
1eccmQUP17WueyPRzqMNnBfeOo+UPGhfx/QqteQCdz7TifQ5t4aaDJh6nyvrejqiPEMhGqm8ICbS
hYmTYl3RoFaKcE8rY5becBahgO35WBYWYWkNRi9+/teLzKfPp7QhYZ3HuAJC6CKlnEz3ThZffE8T
CkFRUssvYointSc14IwYIzhi3czkmT36hl4MvFN1sLqw7d7w47ake1CALEhSDeLtu00r7kpgLTQ9
mlR9wJhdRbidUwwAAJyKQZXsdKyc2Btp5iSUtzHCJIygTrhkErIZCAMnS+dr6wkQjTCso47IIvO2
gYEibIn07M4Uaib9p1msNIidJMzxiNSrNin7s1KqkRoY+sq6rtF9xKvwIedQkKTmxVr151njRIdo
2maXKHYILzYuxDcoAXAFJJCAIPMrTs1uQi5r8adjYZGJFaDruuVCUJ+1OjWQrW1qZMowt/QZ/phC
ckKd7fZ4eEQcMRzzSm+xD0otiEHdLE4Cl8fG/i+n0asfzv2wn7/hOMmPpPhmvKj8te3sLJRTlyrt
+XUOdaxV4QerNbiLohv+yqh4MuBKjBXnChw7uI0Q/weSZj49LzDFGVfbv0sNzN4h2Kzl99b+RTqr
XNY6TqKicQa2fL8xLTiza1aCSHngjCmBLSBsfvmfsYjegVnMzNTXROVRafH3iV09mG3lI1IvJYCw
Az9aPcNHo16ZQMxqNT4bgWx7QxW4FXznGrgWu7zdgQpATS4/jinvlnDdvkJw+/elo7juD9DYPW6N
/qjFJtwVQZLhgapc6BZ0ahcH5B+CAd5K064Oh+kkVeZZWSzdnlLo0J+2tAOaNTavSLHKBCDgCI1y
v7+lG9HCs6x3ll41uRc21c2tcL1aJso94dDcmwckYJsTwasGZHSCO6IYXyTR6U99Ba5hiDuZxQHf
eoUUpgX5G4YM5ZUqEdR0tt7xwm0/q2bTSpBUDfabzckiUk0h+nPkjtv6JYgEdCiz07tneA0a7YD/
m6RV5S4f/+ELvGph6F3rBQvB9xsNW0CTmTk8ypdqjrLTrv/irOrYY343olSQ411GjUfF8daALSE3
oKzx52sN6CQ1YKzc5Bo7Sxripk5ZQyJ1Yn4TVTBkh9o1Kt+S3IEiQOsJEou5MBbMCfuoUZRv50NW
NK5sG/Z/hAHs4OfWfAAIi8eSvrxht7PQoDEzOMxyptBcbJfwA1W3+7ft1LNNrGBVNzGfAssNObn1
nFLfQ+8cgfIwU6AxbBDI8DWhU9xWoL6LBLff6M9idOibfVU3697zMk6U5J7GGuSfPsd5puA3uwEI
+LXLeen8dPQC0RYtSHo5TYuyICtgEFNzsHBoqaFj1jxcg2Y/XFBYEQ2SJT/0ozyh42+kxxVsI2xE
eraxbDAjrAMK93RE2w2r+MLVnvZPQUzJTWnckXd9iqlkSiMjD5XB6HBhednfByQ7TP2q6wLuqwHR
ul1hXMLngxcJZzaJhsd9HU/OoqC/sEUn0DJf0qXMakro1BVmASH2IxkjeeHBgtPQ8IKLEyYvWGT9
E+VY0BrgT/fJBKDJx/3bqAcbKzi9z0SZkd6CTCQ/L+gmvN+6V1rNJAXcwARBnWqwDtdacEfsypnx
t+WZWOBU81bOgQk7aIzo5DHjo8c+zOEq0TCI2xX1dQwEGmIlDYGDq/EIUQkgfkMeM247dydNrKIQ
bnwXhfqO1eBxyhorWUw3gCUYd+IMf12a6zWvAYuSJrXVUR2apoD9xxAPtFBO6Yq9E1H4V+fEGhwt
TjwHKER7BnCfx/mx4IawaDxCoU0sSE/WDyQ/MYNljkDhPuGfYP/CC5GV9kMUwYQaGfyOy2GBJSyU
JxZNxNz1TrlF7ncyETG2DzNmKr3g7ef/USqDKnRU/VCzk8Jhq69Mg8SSnH/yfaTJG+S1K5iaPJug
z8NKF2rUahtBk7Ad/2LQvFAKZlrY9WcGDCvDItDOcZSSxNvm86ZvYMrF3NP0+i/hbBeRbhk1Ypa7
45fQ+4/2qrKE0ZejdrII6dUf5bX6sDmKPhOuchb4ifTPBauolEWk7rLPustaQn6Z+sU9lXhDnQce
5GIcRcUUjEzf7uLcTBvTDF9Wgt8saisDsA1c6K+z8PxYcmXa1XvSvNKohjlukz3lcjiEwCGwVH4R
Ilm0oPKg0kIJOPmXsEXXHv3Wqmt35xo+i08JGJdNHvCiMN/nP1bZLGWAA9aHNAv+1WjyP4ratAIL
2e941ZgI2jk4q2M9fQV8XRPqeyxL8P5jL0rs/l5ncjHqo+/ubpm/q11If/b5/Os9E1JWYi1SloSH
Y4VRkiVF/2IThDbIl53CUC7JtBiemUhbeLh46gBISKWBUwLEa2tMXuaCo30Kzu/UX0U4eVQ5txyg
BSjVMpXINnbG5Nhgg+7P+HDNIvpmFEPgOQy1R5IogjvjoR3nYTqCfYIiI8IC6LDC2ltCuvwWst65
HWvzwfeMEBj7hQ9hMN5qfE+IYOFkRw7nE2eJNw7dgAzG8BgxpouO00FDS6iDBuR2C8jonTyC3PbY
zfkybRETdRpq6WHlsf5KGhQbWEcHf9cEb7d6FS4NQk2DvbpPgCeflBSnLQpMN41plhmLd6Rlpndy
/kwg2ZCtVUhoOzPRcM2bzFSegcD1CM6NVdBvz4LJDcaMCgSy0JbKf3yeNsbx7LNs662wyTBbyLro
E6bmzM+8MwNUECVQ+M6POrFfeU0wFEafflPPgvuddM3CB7ZwQUXeBwuipjzjhXosxKr2Y5hZIa33
2ZuxSsZXL15giDuMawDdl3GjIShZfQaVtHDnoAJzdFrQS3DQ0UMOpOlefqqaQpWq/ew8vaUHl0U8
gbr7pjah0tPDqA8kxdONUmJEGRVOvjAVjYDLD9EFIPu2BYHUOJiyvyf2BSjf38VgBVcmcVNVwVSA
4+Hl6NGyBd55cu5D6gafBgzaQOKRXaezx16YsHGJn38QoZ0R98iuDfHtNRbN0lwxB+QO8J6EcEuz
9FeLYYXuZ5ojGARV5HGo60wqSLBKeGELNUeVoCuegvfbJS2wtFbeefrDmsi/fI8EXKlZcZocPJ0s
HrmDYt8wyHRJi2OsBmJXR2x6wlGJ3n+USSzWU89hDUHtdK8U5z58Z57JT3GmVr9gUTw0k9P61yJt
k290V3vRMHFBjX9oDSUbVXHLdfbUTyRpM2793HbUVRwa/TwJFQmCbHn4J3ju7gEniDdBkiFmOW41
Lczh3sbDqizQQjtQc4jJGnp1QdgU8A/ejqvWkAEQBvwF+camWKV6AOUxcKVHmnxJ55oUv3oAJ6Lb
oXXBWh/jD+KKe7Dr4dXT/iRuqn7HIgbPnX/igWqOHlGvC8R3ZosrpekV72mmOkJmZV+7ca30+bM5
WxgMnX7cdWr7Vdvvr3qe+qO9JaA5YtQ4wqgafx8WTQGvFiWMbnZ570EQdjFLe73yqlNlTWu93EJU
clBuo0WA4YcyoDE/DwsgG1Yry9pcFgQF0Q4rLpgMYXPoZ7wPXpPzPjegxrSNPH4YFmtVpI0e7CyZ
d+Gg/ETgPJC9FvqtT8PujYsIuZwxnsW8Z22nWLcqItfXn25WBZLUfM/GTh/zt0zb842LTiv0WC/T
7dfUW0LkB8SIgAqVKH/TjDD9LkOtUx1lOzmLLW7MTxPA3OHsdBubwzygAswSq16lsEhtHySGDpY0
fQuiwwF7A5+LmZmL1JX8tPYghrHslYS5LhUt/eTvdikY+2v9UytduOXW1cX5QM4c/b6HzW6FKMRm
f62j5xjKvJyjlqBtCtfqinuyFpJrJ3gCcagDbsO4pHC/o1I7yBrXJWkhzQZ8l/P62NkyG2DhsrwZ
sk8S3P6k+OqXqiVs3agtSh1htqUpghmWhzNAZgo/TilaLsdrpfufpUYaql18eMPG6MBI2+ylxxkg
frkOPhkHrFN2jsIkeBT5uEgxIBltlmiKr+gDOhysnKUY0xtuKBIiL50nbIT3phvZlWNdHhrWAtif
Tivz7d9fn+ZZMqgj0nMZd0z+perLuuVVBZuqY2YskHWMAtl8g0hXU0e8DdXB329E7LUDfLaoRQtA
QiUHPz/v/11gkSGcU1baYu3ovF18Zm+DgDMv472dH0c6dfEomhDRa2HEgTjhxoOtZnnruUz/+hFW
ZK+b+0vE7XZHuq3QyKnUGMXiPzXC2oioXRY878tkhSe7o8RMf8UN3TYV2vvm8hLEtYqIFaz7rVRm
CpaxDG2NnSAt8g5r3tXHC23ojdjaJSr7lAkZy9p8XpKxCmIPtA9Tuf724uNvYu/OJMoUHPnyfhH2
aul6GDUHWy3Jzij4maVN1zIsuzT5bmV4K2mMxJdJlPW706BPSEVhvP4snag0QgWrBVJ6WWmxsM0q
LcNfwJ0WMojaU7khaoFrGYmZ7VFrS7xvlnaDWYZzmsGoMyz2aB4JhIdS9obQ+g6pgDX3SXV5YIsL
NvRRk+FJVySKciURVU35MYiH68++Gcr1jqHtVZ0Nqh2c739Q1Wiqfd511t6BfdPeJyZaYmBGjTgS
EnnEZt94Suq8SQN3u3QpYKnqbYt30fUV+YpykycUxdYRycp/FrFYkBSWCpHx2qQbA5oOk5U+nlqs
AvTd5qipG5CUlUT12MbIzLtTQb/+NnkBMe+gFm180rD1d4nW+A83KdZWKpWGLAvZifQRS8blA8xE
1U0MWj05bpjaUIRILHGWDeGTNbLZe8332yjvADJoK1kbFNeb+ZCCr9LnNr9Si/MWWA+pX4AttdoL
RZm/09kAwKyxTRiEJV8hrBTRmx7sFUGOk+E5tCU7GEvAdXHW8vWv/kjKk8l1hPxJ0UOMes9yL1rB
rA1Qv0YQJkRatoo679DUSqBanCxCfYITIRtIXLL6LUsTfVWjre3gLG5yCLzEBWas6dpByaLdLvix
/2S0u0Xn0fyJAG1JkvcTUIFZk+5oR6zMELrZ3bv4v2t2K++UcufPLOplMq7+0J0gha2b/HfM5soB
fdPjU6l9QtljgexmQyGyUO6W1kgEou/vhSU103S4+PENi4QKaHGneWnuRCsxrgLJRfDkS4/+hetC
lPlLKnclLlkVV5mfyr4tG+9DPgLRMOli4KnaAF4pIkt6y0MrIiPcLD1RNeQyWcrkIxMPP+CjWJlJ
NYPnEF5D2/K6EYoXf054CmE33Qm7wxmpohv+J++nzaf4BkbezIzKa7V9zxv3SmgYkdhk6f7/p554
D30l8KzYGi3PcXy0B2SCNUl0SHlFJzWMlzNRR82CHAHtM1mcPGT+8geASVwdfglkFQd5c2MYUOMB
cMBZnc+ed0xdjhQtdWmM0lhfufq2/nAlKXDk9b8CzBlrYrwqR9+Dn8S0BkKmDdvIm2+csJYQKx8u
GVTGYMxA8gys/v2OCyyM7nrNG/Tm1EGbw6r72SHoJEV+q7kYkmrV/3c0nBbN6sIGkf6J1VaCmVYL
0vUCbmY6MABoin7orElovhZjM55pGnsdDsIs1JtrvHHjTocV5qlvIs2rFmJZPjexwOIQba17AFmq
9f7qXZt83CGp4v+OZYkjpvoDzhUugxzhSRGdaWyeCSdFlwWcUzg99yK9xdG+e7kLHs6JiiVu69W0
Rd5VZ9HsR6F8bxv34F8LTMMGid/f3HQ/w8ZpKgT7lCdDuw1kLzoCuAc4aQhE5/mVAw0FqtN6Hzp9
nuqZKQGhR2UzEh3rqIDTIh1Um56rFTjqnsWKkxJQWaTQwoB/98lx84Dx05mBX1CobHH9b+sWwBwm
sQxTLI51xa5n4T5oU/7lcT/1u6EBoCBIv/AcKhZdBt79qTxC6/irIhp8uRf/9Fow6EbmjWfF8qi0
OR81OqJ26OXr+7CZbW5OdXok0iFkIcF8suD/s8r35i6XxUXtDN/AhrgMbU+LeycXoa7zJ57Yx7jA
uKWaa6oAp/1cO17F776vwhNiefCfhApxFE8E6OzH3QIr64sTHOaHIkR1bE9CxxP2I438gor/OT+5
LOpWxzeYo7NiOqvdcqgg9XDh0qcCufc3QDEC08IDJR1fRaWcLQMXscLYg5x+3MU/ceJcIGx7MD4D
K/Q51yIpa6nErM8sxxFdo5SpfVLmsRRBc3bFujM7x4sUWCx5etdq8AMSon00MkwgqbyOTdKmAYE3
aVGlZBKeiAo5GM+CdG8P0EV0fYvxWtYWPdQNAv52mLIyVnpMH3nE1oP/rj5wfLjLfCZAxSgNqWAp
V8QZ+K9ML5JsoMHbfJZgmKZE/jGOdXgmdqitUpDdsTjFWYQwysFWee+6OD4+l0JS8rvR3oyn6wnS
tFnWW+SjiAkf9KJmtKeQhmukceS+AudVuBr/SrayoYfwT2QfG5VPXoUqBrqDFyrAKKc9vwFBglfg
0iidtiaqGTRWHclR1WgO1VMCQwhX/NkY/xO06M/m+eQDNUM5AuieGj+FtHfMDQrMhwk/mRc/914j
LtONcxIVIpAxrmi/b8GFm+X5LwcDPIpOvKi/QT8R6GN+MrZ4Q3oa+8I6xc4GpIdbh62knwuKnLxJ
aOk97/HQ4AfxhyKGJ61yhoUcTQUy10maTITB5vX1EKwc/HHRKfyoFiWVgv8rYG2LAixUKnqdTskV
ZeFiuAhs/eOspHfAffX+B9e40py+qqhsTPfPacudYk/cTCH1jttwku/c4PHbNxlirlU3CJjCh54d
D9pcfFUbcuw7YJN3m7uex5kAYMtF3WV/p7tr26+VSlhcqC5OWjxJzRagJeSI+WWBQ5mvpUo+jz1X
JmMaRrMYnedLF5T6NGSzQYWMGX3HLEC0mCQ1uKU0XBrkDkUmFs3IGAkQw7GNB7Z0vdgS+opFhMbf
YUFeWc4sCD7kAL7lANNBjX6DIOBm6nzltMo5pSlwinIE1pc3LSUysHZ1L9O2NTRucz5hWaDjJeeS
yPZuJJ8kENpu9ex/Bk32JPmRXG0tlAGk9+JkukmABog8vmPLBs9kkqMkD7EtHvtFUhGO7EgFcEP6
jD0nhle0IK48i4EmhPa+vN9cLRfMfSF6OZu5nXeAAKwONNlSpU78CMwPvkfhcUTZxv63/Sg+VqoV
qI8xcWSNZULitxp0eZb1lB1wZ6NQsOE6mASpmDeErOB7yi2N/iEdSZ+aj1XEqqWAoea0QYTLwYL3
IiBlNgwdI6c1BU35aKzglKzpCBt7JibCN9Ha7iNLlUvfm53uuKRlSolMufMAXYzbBkbgIlYOefKe
w2amWSFATp2D07uJ2Y3raumnloszedamTgF6LhIxHLA782qqDkmi7IrL1Z9uZm0Ecr/jEPL99iKA
HVGd89mP4nffcvEEcqoIxd95wuk4MtpGT9igTwMnEh4rXGL5zxCKufrlw0ct6Uynyyu1ZH6YAona
pgWJwNhTVq957GpqEePS2pr3JCEfjNCFmvSKrRPqKrD8ceIaEMGOygmner74Wm4qTcAJW71tbxqr
tINUBcG4RJ7pCxcX8kpUpK6ygaIBWAQCJbC9qrqkonSQgBWRWcJf2d+yO9nEbH4AHqQvbvXpWo9W
rXXpurMlarK9RRdOCieFgmRSeZ80nQ7/0QzO844t8tG0kd+K6wYmTna+OpwcZSJ1BuiYqRIkl5qN
G6hbvz3HBvLRH+92IKZYZQr/XC7ArsMv1rzofDN1dyiOyMSv1tvzjWlHgKUFWCHhrtdQt2WN/W8S
28BvIQcy4eRKwIKF4tH0YWJnyOxgaBSkc4eWiXiygJjnp56Us+o9Rf9m6T+r/U4d91wiUSwJmkYH
QgGvA04QDmJ8Bz6+w4DywEquLblWlUi2czMRCrTuOmC2fdpuA6bJNMIj58BhymE2Ku27HdE3H6IN
f0rHJBMqNJWNC9rz35quwvEovPjcIzuome3NoiV0N9jEXwTkhheRYDxV20244vRNDPZC7pM0YezZ
HVnro4ufsMFNGTZ1EZwOcN5OQNe8OdVih9/UnbZCEjmZEccwwgFMrL1o4Wl90fuxs7KuaBF1tWnA
Va2nvill++xMkW1A6Q6txfQplVrTMV92zIhiIq1KODmov9khONx5yXa+vIdYZRlxz7DIj47Bf1Ou
/cwdOtLRgXE+tMRWzQl9fg0iVHUaB79IomdcviU5fLVvmzGznbIb0c4M2NduYs4Kw1nzTyvlvRRI
e0LOL1auRWRVhf/aN6ce6yTnwPKjfyZ2z/sAwEyrnjBUYGvI4i++o+9hPzb1NW8IJNocScJ7Brvn
+q4QNvQmkk8emfuE+SIFcT6E9DVwrYRh78q0V92QZzL0O9M+aN20KUTGlLr813XCUfAGJpX+ASQe
iKbvWbI50sf4KDCFzZn6RH32cc/RH1CbTuKa8vigZ6CtUqdZMF6wA71luyI+eUl7jslz347AuOJ8
ngMPdl64unfsrxHMBWKX7LX9zOZJ+dZEBbFCja3F0DTtboqqlc+Eeu9nx5qDH9MuhD/N//Tjw8ww
RRicb2fZ7XPGSnsIOXbSKhCyf+wNnxA99sua5XFj5IlHnUTdbxT4rZfta4IL4guoKTr9+A7Vzqdq
+pVoUCOo1OO3tszd+UIsJPYZUNL4r2HQJQkwOg/jMkBu/pX/9D6nImda5/7DvRXaOjr4mtkSPuCc
vqwKKPxvPDWNnP/gEmjG1GKpnR8qhcM+oT3tmVPmyYknQg2aqxQXUVKF6+QaJ9OK3VlqlVHN8WYh
w+JFgyCTJkKvRlXt/u+3fSYwSYhjWyMPTOJCdWcRzPSQLNdTsJrp/raf4A4Vv0P9a3jV8/mYE1R/
ngLi8X4iUhip7Z55LCmLp76e+dsF2QwkctncoMmiInLOQHw7/XN559Clb6q72hA8zKFxZRc9ttXu
7RvXQH9K/YLIsM9V9ssaQRm1oJPLUT9hWlp1r9BN0KISYY26/5fPdcRrdm6H5DMrwIQSbgj4FUP1
79Y9BaN02Kl3fmFGegZ905bt/0ijVNXznCvwVRKqEFpCawxZBbZOqDG0Q5fLrwG9cCnM/a+FxxpI
RHp6oUl4bD+A2C/iSh3pIU7CFuI6lvL5394L3EmiA7tH3Lf+tUodwSM750z2DUB8VWAUsInsPkbW
JoEy8vsUYEjzd4/gRC5BoP0CBEixVazt/Avsv2nClONujA793Yt9wA1qQqt2Ax+N5G+Gg7XoCTxI
5y0WW+rdbJlDHCqf7OGzXi59W9uNfRjfE2rtHEzsKYqy6za3G9Df8aMIvxm/ktgZv6w5JAlwmAgC
8SiLBgH3KsEqc9uDiFz385fsTp0ygQWKp4KiQHAZ1CMlY1jzpw4gB1GNreeIqs7tWj9IDyFhn8ER
kaD9h7y7Bi7SmpSjwhvLtLiyyPLLdbNve/4lGEaELNjl1g4diJ2RiIh6Dpt5/l/B1PQMUgYEWMEZ
H3wKtMLu+odrRd/wtgZNBRD+dvMJ8tQ1DtyjPCGsxHbr4i5LCk8aHIf8mUBYEm7jfYXGG9Wto6Wm
eYgGpaNk/clB++cy4DQ8cCt/TV51h2JVtqmSoclWuyhqKQPAuUwJ7SZBqKrgHMFT8h5hlNBUeOf+
f0H4VmVKfEZMliBsXsvl3CtizszI7F0sER/RsbRYMzucSuAe0ENyTUwR9V3Av98oz0Y27gj34sK4
BDmzFg/dGW1FdolaxnR8YfcSPMIOKNr2YUym2gvAD2rrKULu/5cwbGtlEkxq5f2mJwymUcjS4PX8
cdETrbfm6qpOzIbNLytRifxMO0hkF7SbUIijNf3iWGINrE33xHU6A9i8S+1qXkilkZDJQXHJ8hCq
6xtg7QQoIFYkzHkPnHs5H0RqLx04M1SECuPT+R0BUwXqUAaWtYh20VAbyH6CqN57c/bKhZm7OSBP
Cl2LlbBuV/aFgH62vC/6WchmPcy/3dvbvsm3uAtW5+oJCRPKp9u0kRlzCmhLjBiW0d0X4mzBBk20
YcpA9zZezf0e4y44hmNcgC1KD3Y9l4sR8q5KJXSfBfhT0fwt+pE9DNVA0H08Q/Sut00+P6lxEjTj
X0BHqHUKCaODurkvwF7psEaU0BNI146grS+4237bikh1dRiglftgE16na98d4Z1/X+We8wYVPg4g
D9EqeglG0rwLSal4F+0IIkox8v0QF5uhRq4uuQn9DAokAq8pWsARMWE17AQT/tPrF0TPKP5DH+1b
AKQq/tdE6/Lk7dWCAHNXNK557iKN7rXq0Ns2U85vt2J2VAhOPXc2tDTsZh38z5ty1tv3WONnErGU
OamRpih8sz5Xe9NkK7VrtR4xofJ4UBZHUsLfWjMUR9wgEJ0hxneEE93RD3FvxFiXZwwq8tR5AmvH
dlUu1JK8P+i8OVJ/3HpoXbjKS9YL4zBsWk9V31pFqBbLPNZMxnFRXMme17kS03iHSkKjgM+ZCGO6
I41ZyLNFqAz6eI/KEnWF43jZTjUjx6E4gTau4/dQZ+0dgRUCKfqoJZTj4xQlS35h2G0DLSzEdxeZ
JKcEFXxzhqUtJeJBhKQ/cbreQyguhswQrycCF7vpeZc9uQgSNzRWhl04nxTgM8ZaL/EaHK5Gd99I
U4r8MPqVpQCk2APZaNHvqbIuFtNMb+X1WIIdGfl0hyxtlT8/f6ilofEdmIVoN/PzvQdIIMFJ7q5x
iilk4d8CVWc4uKUFBao/t5YpNzHInDztLS+Oq4I9Uh69PbCu6qZBrmznIEyaPg6GQk1M9tecQv2F
p0evSu0zSY6lZ3CcwYTUAjkJI8J4w2/34DLuz3jIOMaTYUrHZy87nnXp30b687ekMZKr5QYcdBjn
gFjHxkZNeNrI1QbwGEIS6icZvcBJjDX+TSvVAqBTpnwMDIfypc9qR7rh5yBJausBC7P3E5KjIBqd
/ulzaxsrmB+FGbazsnjPTOClLA3mY/Od22dvmf+oVIkdRYBmOPq4i51MR0KCuVu7O7KK2k4y/30e
rQmiNLEq0uqrL9OgQGjOpTsyQDONwzsAEuctL96GC/fWulEtnXbiustPcOGbzmw3tJ22b88qDLBq
gPYUnVsw+OLdm12RwleeSqOEeOv70MAWSHwxmqWLtkmheUs4dDg0l9O/gh6RkUQ7CmqLQQChdCt+
VQwtVZLro9QatLuBLWl/a7CVfE3/Rai1pqtsXWaXwFQYiDXfKxszyKJb6U2HiD9qYKB/clE4lXAz
y6rRgeK8SOaaZSDFJ0djplXn5yJgWdU4zLSl5Jgxfqg/l4wTDfSS1I777SVTTm9o+mQJznCEqkXm
FcoA+V7k/ImXZNqSh6gs2K3vR+5FMhYFAZon0BWv+rVPl/RD6b2huc/OFYWCPgMU/fN9a/YwRODj
FFR5mNXZbWxGR0xHASfpzrUST2yo1Aqc5WfBGMnFsm4keXw3YNCXXwhdkOXIK1nr0TGxrnm/iLMX
tW4uQaD/MpMN++D8N9n6VpF1Md90NJ2O7zzby+p1eEDB04t7lyaaxbF8KiR7yE6LRsLuPPZIerH5
wvPghD7Y8VnRbvxHBE6XbfAHvfdOUrvPg91t32zggmzfn8x/focApRBGEIUeB37ipB2P+Y++Uqy9
SHNpelczf4auuPLhZr8TQpZSqSquI7wq3aVQ/jkVSWCubTJbIc5pKNOuNuKqE+j1SmCQBUYM9e0a
0Mln5FZoSKw7VBZNtDWObeJEDy52ADdkqWfiHELvSVhskkJFmDn/FIaMKbMaecg67fRnGvWRe1KB
+1wzYCNAsD69/V/KYhUFZjMMZjia2BBINeDinioU50GSYSLGDPiUzZrk3BMdczCht6+OZD0x56p5
fxxChfz771Hn81B9tCuWXMKsG794DadU3gzD43I8E2vcIbKHCGdkhSJSxFxeqVcJGqI5ehRwNQPT
VnDR0vLzcoaZDc/3GRMinaSUsi8NtsjuJIY7p0zbIFX+3WTyXb08E/bIrrhxWeXu+aArt+j4Yfmw
kd9OOkVTKBf285rtFIh1qVJMhmSm4bel+uiG4cra2fnj2dd1R+Nbx2HAs6917nPNXUa7sJXKiT/d
z3FHTxA4BU9IFTHW+Ib45KqMqeszoO/e7WHglwbi8vAWfetPSgzqRwwrjADEiv+WuH1marXyhGAC
VSzVgE2jBs3H86ueSlDnW6s605I2bvASsgr4p1EOctkRnOwfuHt2v/tiaCZc+DG4HjQggx4Bv9vI
7Z0a26JkzPxOH2Mt+lksXR7DZlNSb42C1jLC5pK2N7xph194GsuQUv3eKNWW+G5oeXT6XALCtlc3
1TPnJOfzVL8YibtdfzYKxIL/OH7at+l6AK8zBUYF01svtt+M6KCOUb297c15bZdnxJevc70yk1qr
68LrXvN0nq6At4stLtEgEgQblSgLKkSu5HFs/lXy2J+fedoSZ3hb9X4lKN0MYw2N/eb5MeihUt9u
fOaQt7ae7OTerrEBDZuhBpzK0yJhpzj5Nel3a8l7yaWKVXvpM0Vm3NChFY1GyhhS/+EsE1Z+6Hit
T9a5usyrOoVJok2SmiQ8S14KI+1Hmlt4QZIw88uIYnraFSknDO3CgW6bFcPQiG452L4QYKHopA8j
ec3DAzqssVhHWjt1eqMELgLzwQq3zpKkEKte+n5DyoF/hb2+YUGB1fq1zmypCfAzQpKh1FLxlHu9
vjxPFcyAj34KTUvcpzAYHrLz9Q041cQy3VH94GhrdludO+iTxtVzJ8Y8LNlGVrXoOhBqXBrFCFBF
W+x4nx6cTnJZKvB5WWyeZl1VSPVWKb5oHc3yhxnp7UIpuxLbj1zIg3Hu1XKdzeDID+syTOn6tBx9
PhE3IiCbiaetDMPeB0i75CmUQNravoBAEmN+2BrOo6ePVrJV8TyNZXcZDKKhMnHymWA8jLnWIXLe
6JZ0Z5uzj67yxKtSWca+pB3yKIf3x7mkW+3v7C3GJgNfR/gHdxGUT6nBMPCtYmIof4cfWGtMxl2k
6kL+PJAszrBssLyiGCthpCXwripOvHcDe12FlPpv+7Scfn1hkttRtma4g70wpS13grwXJzT0NV8H
ZEByiooBc0hPqZW/G6Pk07BX+MCeofgXKJ7dSVV+oqKHpHZnkZU5yLDvDPWT0/dlDVU5Pblgyr8I
xGMuj2Z7oyq2L0KlT7riq9fFsESGxhldL/in3qf7TrNCYmATAUTUw6SKB5yZg5RCtvtJ3eM8BZ89
Ak9NEbI2OAfaDZjFvqLoRkAwdbRgM+RIEWogQr/cZwqIYlLm4GW2zNuDAkKMpWRAdKZl79hqp0We
+bta4YeIbvo44Ym6cAEkiXcRwoisneYA38u18Dw/KaLJb+2QkdL+GLxdD4aPEIx3tPkHO3PIVden
WjxgpfC27/Y3q6XkQyIk/B+kHzs97+a0GyxjxFWtDXXBTQGxoJR3ogZ5BiLKjuZavvUS3t15vP+q
90b6qhGOVDtkUvry5Bp9NJ2Ird83RV/tjgXUbe2+OEKE53VajYh5iXqnESO1tJgszCC73Mgfyebs
lds1ZTgAADmZo+XoLQ5WcBUqY1m+/gBASpoN40k9Mg4pcMj78fjnI1mI9xg8XYny0wkmlOQTs6SX
glFZKsiXyOsHUPdHIBCf81PE9KoioEypdreoe6WkzH/y62AuZCwZg2YCh1YV4Zu6iUFyk8Zg2J/i
/c+W2y6A2yY51qQ9xyjYAicjdV5m50VCKRO5ZFC1myNaT44w9ZwlV5yz5RDh6HvP48nAfdIHeV+G
kCzuFxGsJUI9LRb3slmh2xGVG9tOqC6aVUALIWcxLyrlSDnVFbP0wVOISxpUoWoL+87ksPFLqs+w
4oln5OINk6HZ5vAekQomX+4+7M+WM1aBCwiYDuZFk27NziZKLQyKcLU0E7pL/kJEKBeMp+YX1k50
x9ykh42wna5xgqKl+biE773SfP70b/wSwvfaTf8uXmBLpbMZ0GtbboIBL6kEnudUWPkJqlbAIsF9
Gh+fbwZE42TBRnXoQryylgcFa/fa8nkYmJDrDXdbJSPXlRyfVwOPS10rIadBvEuzlSDlGxf+Et88
vGf4Qk/hFRKzX4nwV9RpJozSp9H+h9ACBSvINBRT7Kceo9lOIFBKTUVU9bmthJPrOrjx1lQCBHC0
ApuyWGN3qHS/aGOWyWIBf8qZ2tkRqpjtqgrF7VeBOIpLp9WYQNzdrr75dwavv8RFX2XgEOcK7TOl
9DoDQ0BkQilJSDtCbtpfPNJ42FDDeASAFAzCGKmX+OafQigC9ku8GD5quNOtZG1i6K2UzIPsRztu
TLbfuqBMnnoYLmQ8UVYvkDWrkTEPVL/6MlLGIvYrhvl71dzAftAA55AQp3CHmF1e+8On8jJI1IO4
ae5BhDzq3DLYxcD2ozWcz1Yc8X4Spg7hVDfgaCuzJQ7TVdtZp8MpoTcqGLJGH+aEk7Q6tRWIQMB7
yhzZFWxQSWdyR81wAnh1ngC85puoTdtzVP63ec42FdGjZeM0W9McKCxCcYtTEHRE9NC2IR9EW4IW
KlaWXeQVRMURcP+pj0sPy6V514Lc2H5qqTywIxy0LT1CtAsglagbwBoxlHtY0xJL67j0ICqbTgVd
NxW/uxsJKyi+lJuxKauFbB+lvPAeYdIYhio9dfynfkqUk6WLwD6RKSQ9AYj3poICNI7SwSB9CeDg
ue0e/iQKfH5lNbdDdakcZJzzEt/Adyb3yEgSEAciaDN4535QAD6mrOArlAhf+qqiI5mic9S2OhbU
JoajoqlIbt1on/ToLOorNrzQUHt5HVEN5zFxHiivDeBGhXEVceAWJJz95AT8nBEIRm1ZBBVNzbd7
fqmE2CAEjL4sIgCIbY1I9AG+57qQzWilTnTRWuHvfo+4T6iGlFbqntAErMVXxwn3dWit5yzzn1ik
I28gXDtIyyXhbWnVzxMCt8SEUi6ZoPBEpOp1mRd6XKsIw+ik8kGvlseU6Gl1w/onse66opyGv9M3
Ra1PeWJM6RUEVg/O7/VzEH5QpR3BU3S9HPnQS73WWiyua2Cj6/bknpQDM50xpALBgU2tbpo+HjYA
OXKJr/N3B0TbL65lX9u/oDFU4FSWINe+ILEiWDQ4VjQl5j+EvLHHYA0GlfMyC6T6YGWtTHMDh9fZ
09q1yrbeY9hDFRao0UKw7ylzSLKZkUvpMBaoDFxIZEqY8t6/uOB7ISkw8sEGn9uRNCwCgUQgQci6
l2HxIO09hIerm49pbyes4k2h2t3qXWyk/VhlruJ1Pmd1i2hd6KNgmVzxpwBZLcPRPR6fwD11QZ6W
KEbevH7brDNb7zLRiZqK6ej67hEQxCfyafezS0IdAlXB7oszsJu9o9zznJkSmjdVINfzSfa7OzfU
4TfosD14zX4CiUPyVaVrTVf8cfPbkHG5eiOpBs8m4vC+dXeLI72ND+Tm7FbrdLaKnalE+sh8s8fc
P6JVnFk4KD7S/ILke8WgeOnUp1ZD0l0DXIg6uxkD8DcFSHRWN+LKC45YsZI+3UykM7sjjpYWiD3o
b3KLDXVGNQjqYTInS6l2gOYbbCX6T9NLT8RcwsHjpgrP59QBxI6UYlHvT+UMf/Xjor9l6tmjnwV9
cZL3tIbpYumsLK3enP6yOXVqY78GCVKjKiwH8iTq6eUfMHhCYTiotPU9ryiN3FM5+FmQ4YOgbomJ
eepOJzqfSdFFdrmPaqnjW6MiIFR/oVLTNr5tSOCpdXYji0xr+1HX1WPCj52IG6EqI1jjRbVZZ6Vz
WuzRTtDYBryUgH6uKxtQNnJ4OBb7DnK4wV+d9lr6toLFSnA40BtLy1ginEsCH2d2QvpYLOJJblT9
drFGyN9MwFI2+Iw8PMx3TQ4nHf9Su3/+Ri7C6m3d12y9M/0GJ2B9w/JPjhfqRlWo9NOt/MmL+oTM
nbpyVUOvZm2em67vEa5uY96qME/cwmT14d0cisQ5QHvI2l61gyy5e50u4M1Y2+zoio2fz92RMHxr
lbJRawvjYzD29um1sywNAyXCwSazG9GZySWrxtj6xyyQfgsnlwqf6SBxLRwjMZkLhMpf8a5rd+lS
7t5xapnqFR3vFkgGv7Cv9spXDeAfhDO0OkDIkyAN2y9QAeUvL8Mx+gYPqaGzR0dlaKb6S7IqVdWt
Qkn+cZnVrjJdDtdVKZ1ifi/oR+Fxw86UMDP6jFW0ZhZAO/Z9gmv34b4ZAMn0/Hr/gAfnY0FLNic1
gHVt9l5UX+R9upty5jOW5W7CXQV+OH611Cow5QNkwQXZobOF3rI1lVSdjYhQwDXCYoA7U5fKo6BW
rd75VGnPPNqnKG3I3nRg3lhcnEX4pSAAfMIZe4WYA9r1FSXDqWQGE0QRsOYMcc6CTS2FPEUEe9b0
KAawOvmIe16Uu9jLomapIWcqALLqnRA1JGgv2XVDN1TiW2CjmX0+GTaAgXzRQijaT57us0BZbBbI
jYaK1EDeDWizzHASWMA6utu0WPkySbeexzk3dlYP33UohiAXjeOcSLH1NTcKsUfHUVIUEV47dNPo
b4aM6fHUSHmNMw+p6BHei0335nERaEt3WU4gVShQre3ag64uD1ig+h//xw6RawR5tavSeU3lzKzF
0JvwN09UM7yo9fkmVDHObeiPOy8p+tRwtdblRfiqGEF6poeN+kvnLPcwQFsr27BxJmKkA4IZTLvJ
GpKrO+NsTyWfON6i0j4aWZ8VnP4S9mpRsDOWCqK+KIr59gX5a4bUSo8w3Cz4DeOJ6IpWWXH2EcDG
tk7iZJvDXQT0K29COdDvYoQ55fLSZV+RTyEXHKZJhkkUP654vMzvllvu2tS77EOqBcN37UFG9bm1
7rPk5h+rgL3WWnaVG8ey83CBQPgxyYv6YX945g72rWuQkIZ1fsEHJiEWF19BMtc5nus4ZR75i2n+
H27nozwCwn14CTJMYaqL1GvIerKSNMaebqSl+iIg8x3SpnvoEKnhVMkBB9JsrAD555KaVZb7Dg7/
fhaIO6V5QSAcBV+vOTBHPEE2UA73wWtwUnuY13xP2Tsg80i61Q0h1syms9FDYtvIZdQO0A3bpYDP
ali8yfukC7Zn3TTI+1uZSvYsgqCj9/hIOvneEay1QVMNpA8cfGJ8HGLsvm0its2Veb2syBewy/Yn
vW0ZvcqjRX7uRgbj6yLgTetyS0S5BADlcj+yykL1hyhp+e+HhJejlZnC2XZY1LFv//QB1k+6gHyp
KueAPbTmnnB/3gOfD5/TXt6YYnwfnwVgi/OXYGRWlU36hCB2yLjj3v72BSt0diJxSU/KTOpqnT07
dN2vSIm2jpeHRvpgYuIkUkkQuSdWjQX5miTzTYYd6zNo6omN1eh/j2R7HwrgWrtNfKVsEoTU98dm
z1hbDir8CwrzJ2yK5vwKydwEm8ZsW4KvmpD73LPKBXqpxkxXO6WV3l4Jl+qYOrab8dkcx+y+3uli
5et+bLdhv6+cuPx/FPaVj3ZcAyF++3lAUiejY65ChuaoUvcefMEN8MqmhNHLYkTZBxJZ7kCtGELS
rRgW9Wd/dc9SlaTct88qo/Bc0Xu5Pd+PjeW5y8hhcu4D/PZNYIVWb6euws7RBhqj0tlrjkxtDNB/
5zHC0NfytPI7cuehY9yDlsB9GomXN71ff0LskJeID10pPff51NcQlzytT9irnnk7bgEBpcjxBa3z
vRuImV8x7c3gOLBT2TwmEG5H8SvMm0QNojWAzpZ/mVCsbtw+w8kO1lU98DP7337A882lgDs0Pist
62YOBq8rJ4f0/yhEGTvk7GVJqtkHa93vjlwTPwff0wOPVZIrCG8C7o/K39nqkiy/Sl2sKl5gfnfB
R+CvaIQwz6Dfpevua1wYXmzXTC7a85VkeZiKvterqnjBc3IPxYrVHImqDWxIOzX54HuW0Y10PDhh
lo6UqTdTApnlEDpRNL3wpQd81UPlKlgYmbFR/nlLJaisvVWGLl/ZEgKDNZo8afIZQbDIR7goB8hs
cC9Ypxm7OzTEoA6sKQzEBYLShnr9zTaQVtMMzm3Uxpu5FFq6VzY47WYF0wMyBdA+tbTmYFAIqIR1
g5LjerBRJ/a9XUoZl3spW3QBx4FCpxwc8720iFAtyH1iKw+Qg5YEj8Ll84BOATy+gGrxDme8lO/p
TEh3xzgaVFtyxtayNC3JadOfNsb+pcZTM2P6XCkHWTOOfhTqstucDxQsdyj2KK7zSWyIHjbhjGt5
sJPiC0f+DO20ibtYwrG5g2jZQ6ao3/f06B/2JRo+Gprr6VCD0qGE8diwn5UF6RwsrD/jCjAoDgRx
XVA2RuSfGLc/Hw7duPgkZGnez76dj2qz3ePU5t4ddCOZNE8k6bWt6U0+/wKfNk09cU0x6y3oRUvO
y2TA6XPGCRqBIV4rQZU2rlXXn61LREOhZd/g+vG7i5LNP/WNBZjQs0gizhdMzBeAkHRTXU8L2iAo
94Om/dZ7j8wvuQLEdUIUtzPQokwjj7wHeXvC/TGSUklzQyXBtcMKXoz6m9EDHKreBQd7jKf8cXuJ
/SCPeo56tdc/PMeHU3AoLYzvgjgfiIXMWhR+AL9LnR0Fn9rBDI4w2DGdXowg+ZLkoyS+Kb+72nw/
iNdcEYpmtXfzVHfeVPI/seyk1++B5g14oX3UZKYxKlRbM2dpQCaUpi5bqxMCLdTKSYA1aCJx4i1f
1iiUQFROblr0D2+s1ZtqHem3J5lpzSmjZjJMjN4wYc3pJdWJp7aveZEp+t0aJOaUgthyYXIa0PuH
qUlPuG0zOIxwh8RSx3cKwNpiijnwRrYf+tIkgwspxIuN4VCANQAhU3UQktd6dQYoavuT66vFt8Hv
5gSQX5h5IBD4c1zIr6UlAKkUzbwZW0R4AnZRIxiQEn/7s5N0/+3yDXekbM7ZLE2NIqgQls4pQSXY
6QiOAVAMWzoiFpQDpgBMTfVmOWeRMVKDhTolv+P5uiFPwkTqWFUy349CLQJeChdMyCjSxpa9fguM
MtakzyY3p/nOgAZUxnhyI+wx5/5BIh+7IzDYTj1k7djNV9Oi76O51Uc3b3VANiN/Swryo43Br4wm
bBe/AGcVSA/Wios3RNjeZcFDu8imwcbSRw38H4ZrCHm7PhAerchSBa2YSb/gY7bWYIhQdJoFRg6s
TdrhPxvl0GD9HXtged66WhkybpznAbEyukUBXyVJgpCCNnfo5V29sWp09wZ8+rUt7x6kfSRZGVws
Y1WeDXAQ+PKFaiHtAZPIDCnuu11DSXZuj4DUleQ2/IDBRvUIZjW/4KGQShpj0NntPEXK4OVX9GJc
KroQy/q0kblrZPOuJMsmgqqBzlei8uw5DYYxDoQkQIdX7YKtcxfipCJc7SYOyxRvUEt4qFjxFowp
I/ufY9YFoEYV2yjesBXLCgMOs3cHPnV26HzcM4TpsbBp1MLfNSJ8wdhzW/4QYniGzdaZ9DCH4xeY
PJBKzXMTsQVIu+IbOIOObMPpe6S+LtUdOk0FDRDRKTRDadkYOyWBq4cw2/T5je7OySALXEzvc/RT
PQZ1MG4BX23AqFN5tv5miiGWLHOQyrU0RMjr8Qk1wCEM9z2FQrml0rb/aTKH074YXUQ7CyFwsK1V
3cOk7Y3w8mnDmIaB5aAbwCvzijaH4cuW400BxoEgp5bf+FZFcRFTnynddleiIeGXcQiHPkj/q84V
sn2hzzxZgq/LHxgXwajQNgKgjB/q+y6xAUG1MBI8+qgGFfeTVMH9zMStr29Pl5Q3TmlX58FNhO2Q
FrE8iZyEdIy7CjaNfQHR90zCK1s6dV9zKrGeXMlA5AIpGXOP1rkSc6dbyi4Lf3H3o5oQBPTKFHgm
CCfz/DEO57NDOLhnMMKeB/6AGuRIAY8UmfvoZwfhne5HGBS9phf+GTi0LvvS35e6gBHysq4HJcOz
AXqDLio8I/QpXxWZvdMJx1UsrZZq788rvtfgHv/OM4liAwHj9H96jcU73VHZM4Douavc3jpc0/18
MQlOBPKjC9zs1DKdvNfzccQ1gN7NdzgI6Z+Oj+XN1s3jaBab0d5Iz+X9NhE/rzFPt65NGVN21Ci3
ldliJlkQu8U/naVDmt/u/AjpicwCptm0kbf32RCmzG+7y5acSqcC+QWdNOwWWiIp4J8GVR+lwhx9
+DDVAcqoxXFri+qiqpBlt1Abfv7mtcd3Uuowkz/Tn6l6i8lq0I0pPMzoh3iEh4rE9E87g1LuvIO2
kgn5NR2QDIy4ITMcl7GvI7gYDKbiGORBFReupAa6ypqupB2o6PY3Ltbdr5bMffib0eyjyhO4hLun
xLpFk4SG1PmGLt8aPQGUkAml4yTOFOfLNNvwa4zTNCpm/+VZXv1NiFpcanJqQAMfamYiwoDDZ1sn
m273ONpWJZV02VD7sQQ7BWfupk07B8IXwZ+mSGaEHdZrblgf2hEFtaU+ZNh1MsQGnCPsGjmbOMy7
CrV6LSjrgGlej654V/IIfmP1EG8NrrHK/fDYs4WKa6xQwFLu7OgwhQq5zg8/jW7VakpaktbWN9X7
emySToEFHT6jTgkHyOmNMqfi2qED40EY5pa19QKfNvSHP2+WDDSdA9AvzWD/PmVYqmn/5u4mEEnt
QwRAMhI0cTOU3e3zEF5w6KYajIVNKRhjF+thadLmz1DjqLG8d3cX3LDSwtV9lhvbKQRDEIZJWl8F
CEev81rYPTioxMXe1E+l8SxSopRcGnMmzPwvuQGHh/IZXTl/EHvr9Qul+9/TUaiq5Ib5XBvRRcrz
5TJpVZqP4u2vbR7UuJNbrr59YsU2MOMNNrBsThVgBmL6mT2x5gp46sYnuGyZ6uw0xRc3elnxNnDl
YaQ+J5Lb8F35f+sW4b52RECW+jPjjJ1ySQ7GpnHxk6+Mzn8cBph88N7Zi83nKa70gPs9g7jjO1ig
908nOZ2dhQ1uszzGaDcBej5/Ens/ULzYQlPfHnTjIf4B2hUKeHnXg44R03uYNJ8GEd1btYEd7ZEk
PBiahnWpvrxSynxe24a5zvcWLDiwAK1GNHfbv/Tnzs3LZJj+TYb9Gt9joDanfFYjvRTe6aOVKY53
vzlX4AOM991BqR5TiKcVgSilR3c2x1SD2NqMLzxPW3y7rLOP1NHOu1cejoBBi18ZFC8ojwR/j0UI
H+JbltYo6U4I+LVMc1bDc8HZwMzAGBBHEoXO4e7kzftouDEFIMb4aXFgifc03DfJolfAW8nGYhTG
CPt4Vfa0IwJSQrNTBrW263vmv5v8+1P7XEkC7FEfTBJW2uzdm81kKA0oJ5kgOBPXe+IUYPEyYU8z
W6PkPx9zTchhLBzQvxmpvYbtrWY+hybnvgNCLiGX2c0Qc4BUaQnYO4D0okznqXVrFTLB8Dvc4wIq
PIII76pTMjEQQooqnIyUjNmt9y4MeIEF+vHx0o2feVdwqrrQ/V+vLA5geXcTvD9KnKsXdZOg/0nK
8q36eiI2hNqu3BY2r6KCavjbz/+sn56vyHw88PSQTXWETK7ZLf3W3AzcGs+qlePZgTp7dAHNO31R
lsVsaDUILkj20PTjnU3qmv6ZQBLzOnYVhwFkg4KrifnIIqD/vvgfX1TUXMvwdOSRaooG9+cL+TCk
7/WK1hsr2GmK0rkl+MtqXe/PG1MBEL2LXWkUyLTe8rvafT5+hBuDqYYmN3Hn9G7modPe41JteU+m
o8lWbZijbJGcCWChfga5XwZHfypB9+oWZAWnMFnrxKtYxKDmC94WdakvW5ajTMruh3Tgx/S/77eC
ZV3AKcivzDn8Ht1+yBj7y6J/Mv8P71hcgbmgZ+J3nKFi2Nq3n144wroJQ332bX8ottRXdGmsR2G8
hXSKgFEIjiIFxx8OKT8bjLWKCAvnBePkiHXtsinhXOrOrCXJDf+79urV7Ya5FPPFSqTgGpGfFZUU
MGlc986cQN1RKtYrVSkVJFFwhQC+hy7ftCCkYjJiHdiSo5V53c+WZKVFfrZHrWsc3OinlEKcxE/F
to3fnkjfAo2Lz+ShJY5UT6YLMCosiPIGxgx0SMAFRY7IJQ2zH1aUGkOGzT6L7T/euNtonPbCXbuJ
07874PlSuzI7DrXiYVu6XUT3erNpMeYbQaMv93MPI+NKHXk3Lc0lYVcUjRMOi2X6aR3KGIUmIO8i
SHZEUD3pH5eAAHAzdaq/zeGZUnPR8W0NJTqLo1D0re50rvuXYNhxPUQfUf+wrtREp3vxGeVMw/su
B90Q3381UEanrTazVRGqioONa+TgJGnfpdaMPoe6+a+QxU9COm9Dcyt4flnsRIUv3NtpA9cjC72L
kTXGqSrcsuPj8qOkX8wNitSwL6Gdf7uR0h6/nMDjEp088AaXD00qUHFobBpRV1En15elEmnOf7jJ
SkZ3eazHLxNP8CQLUZY02xsAc+B8j73zXLYV1ldVd3UDQQ1IqGUD8/HcNKBT0fWk2nVyi9wd+oa8
I/O6BHUQ8T6224Aj69jxRyUTofIZsW6TDU5J3g9CMR3pDTk+KiG+wSyGAK/aOBhsXSkCJhfoBRSZ
ikbSoK2DiKEInfEe0sArgnRHpO1yAWSowQlIxSFY8J14U4dsvDddoHncdJA+nbF246IJzdXi9Zak
hSwKELhhnwogGCisjzfSaruws8fBREqxu9cYDlLTZtJu69FzJHqCvcJo6FjVDmlJZ6b88aKAZK89
lY1X4Jg/oh6+T1B8XJLgtzr43x5krG+B617j+PE25jlkGusG0PGpo7vQ+XPy1cCEUB3BaDbDR9oR
ZH5NO2CdyJMy0xj87Bwfjv9VVWLlS38PFEWWIriZFrLbVG6y++2uPyXxgy3ItXPtbrKUGHjxWfzT
hly8CDSNVfyZ4SFaLdtXp6Cu+wwi7jHJwcu+c3JYPyffNmtocREXeS2+LhrPoSdMrpEakx5KvXHT
8V6/LH+1a+7bhd1u+YeRCTsooVkfffOikPIotjko3L9gUGuFi47CI/TRH88sxn7wgoeGdRKXxLe8
C1xbZyM91Ae8NaWGzP00pDuvKTYYzpVjJ7GWevdKzQbK/QI6e+m9mTiMzWJ136LsT9Gm3Elv/x0l
tJRpOuLxSADfXUQQDMm8dAM4oLeIATZY8ZHANLkwviGhBLHG6z73avQ9GHndLwv2pnTrge+bU2DQ
tKkk28T+GXwU2A79KY4VgJfZC1CHOTh+D0Zhq0xwsO298aaUbS8y3crIyhgT4q51MnhtZ+qELFW/
u+uLqXNHjP8zZUdnLqoIzj5Py4HuJjfnSFTuXtAHvhRR1J7IfJEviRxXkz8WM0HQTZ+Eq1V5Bc4O
XG5Je9ycHrEXJdOPLZSwa8E7aqxYXExwbaPg46MOeZ6TVkudxK4AqrBmnRA6ToJDYeUlqfS5VeI4
eBvGfLwDW5pjFopWGuuDXYdPSfpxSAt5lZp5uhwScYGD9pwh9GXKvZPkg0t25HP6O1RJ19KbdCBP
b8R3FOrEdW25MfsB8ggf/68M9WFuPPHeIy12I8aQ58S1GBmjO3wxvSGSaAH5q9u27HnAAsyxKpE1
zc0TQb7ut0bVJZdpRnaiO8FIYgEO0GATQVY2c2ZltIzouobzS8Cpdt08AmIfKHamj3qGDhyAC4ci
OdVZTnH2wl2+eYLSmfmjIbqFHAfbGJZrgf5fzpyOccro37c8SYou0BhrDF2CUEmYw+tnWKmYNAcT
Khmaz/zgF0RqW2aWonxamAuSxBvunvm87Q+V52aFimAUmNyDYF7+EWcuIUG4f/RZCeWN7qPf3MKN
xRfJIfv8rwt13Mfx/XkB1TVtjdhUgHdDnQ/m7ddwht210tSMh2sWrbmQDTIQDHhL1rCc61zZC0mf
1PLSxRHesmUaCDO2AewmfG4et+YKYHh5FiIfWpKX3RAyGnQrIXQ/dnMws4re4Of0i/xpgmV7KMT7
xA/M1JYwnO3OuS5esOj9yctiYTdUqIGcUfrILIQTN6eAxzT8b8CteX7r4Z5t4YehU0U+nRZY4er9
QJcphzILMDdPbaieqxcHCrA5rgzsEHMdwkoIesfNtR8xZuqYfNTshYGIX3v7JdqVXIkqW3mdVdwo
r4V0jio8XTcxaSPh9VGs+G0JVpCIg0koKWzUXlDRJrJgIMRUuu+GORhKhjHk79PRlQ0xC6amsxEZ
AxAA7dD+SXHG0HX7dWQ4SW5AyODkP/0cCMv6caSM4wwShPR0ynbs1LRE7p7faJ5XjAhSlv/bAADu
dxeJ9oUtlub2QRSU9J8oZ7pM6QrbKpP8+ROcAXGtKpvoyRnubnEq8aXolPQmXwxz/3Yn2eoyPQi1
roen5wxmkHvdkMQ2spYGmquXz+eA88d6wEGHvmyVcYOViMhfhjLNXnlpI6Bpn4dwwOKSbMA6QS9A
H+Qt8TG9BAWJjCIg4CBx+pTfzi5naS4FjwvHrSiTKksSgw7Yywed1mObm79ognryeQQZAtQV74vq
SPsxL9elb/JZMNSCiOgPdCqYJoIMwD4v3h6mXcfBiSjkdmBM/qjPhoS74Ym7Hp+GxosENqRUTE7Z
Ppk9gAVncwkpp/2uPxIfC6f3x/yAvprd3eKqio+bOxh+ehD4Y77MKKYZj8evZ+DyexUYjzJq5RIE
LxgAwSX7zCG7Mhzx8eLNfbLDzQWOq4oKjXiord7OvKxoPcCIxlsd/DiWB+Mn8Kk8ZDQ4407cKoRp
ONe7NOINlmlx6RrDSHtut+LkkCCk6/84RD8bymOm+r0SgEKYBLP2XZbZRn+aUWJp5g7Ej3lR5AmK
v9896l4MciXKceCeLhAOO8WYiWn3NyUy+FaWrFt9PU4xQ7QX/Izbd4ZXxv9T6iBwNiXsMAW9pdSg
HUA305B/aH0Jk9orLDsKGwKb85gq8sDRz4G+7ZNHGeAapHaifUbHdWfIOjSzdR6TcHPJex0N3o+V
lISIIGoF3k0EAy2UB7QIAIe7ObcX8hHVuLRDUwdI+wg9lOOpdpM244QZgYBv24qsp0svwBizpsap
YGI5xE+nOP6nbOyB/xKxwLrvyoNEOm67UdwIXs1oUHhn+rbPWfiDurnwHJa+MfvRi/K7/7pm+zKM
cZw7i26zDuaygNzt21vRNpLlRMmBgjoTnZE1eEAnq2R6LH4jGw/T6DGhJS3U61OVhdLCICZ7jPp4
2MDvap4av2Du6cBldpuZlBF+YiVzdJgGLsjD45MTiz1vODd3fBkxF7+LkYHg3w0yaMl+WnX3HpZ3
yWRrf9bg38zKOcysR9zyId2NpuBhWFHrPtqm0+aOc2eC5MWvXCLEPhBHsGLbcN9hwJJJD42mFj1G
3+tKlBLwxU8Rfc4I2RUviwctKOVzTKIAngdfYBNoAFXUMIQtWl9oRmm76c/K3/xsmT8jltJvuYyP
B8ZRt1ykl3D3fHeUOcR/HJwdP6hsFcfh1bRwtKXNwJPg6g7utsBf8j69NHqTiP23lrle3QSddbRk
5l5hmwom+bz/RggOqV4jAHPCe+YiQmghjtkMQbEkXOOBLai5QzWa2S2NjFkmeTHJgdbcyZLW+9Fv
egWqPYD3bNuADwWN4Jht+HfxXDvgxxedGhS2CGrkg0SBcwUW7/k7twPAXR1BtBhIUq4oRc+HUkzN
xeB7LKWBSAw8sV04GpYuCM1lPnhy4/rUlQPnX1e2M+wSZiJwzg8brOKR2TJYBOZLsOdGDmWymKjQ
/klWR8ZMnvC7v5zIaEjfXsDxRQEW+/yN90Ku63KaS0RhiqW0saY9T9sgN9dgzqWOgt7+siBk8pRi
37IVcLDVRXM7fLuXUNNpcyxXz/KloMM19IMRCGW3ZcwmOKu9qu4ooX/1uzPY8aJtd6YdswL3gB9s
/bMha3L/5jb5ReEi8e1yJlER7MaFolB5Hjr95XtD8QU2AT2wP1hV8Dr5U1cYLF7uQez+foTTzGX9
IU4IC7Tj6yeYkqL+dD2gz5yAeZl3C8rM2k6ODNZuGkbVQ/CUVhsXUiOb37aJR7yp+H5p8iHTsxKx
pYJPj9+Ntc0ILwfZCuQWkMrhAniRs8trstzk4ZnQrXamFXOP4X1kz4vwmoV1EMCFuI+Cbf6gSl4n
Whe3RBbFEv46E/759OMmzbgZs4bcBnp0jX09GWlSNRppBCEJgaeQR8pNPVe9WkoE5sBndnqvWsGM
WxezxYEk0wbKFRpztJ+CZI8F0yj/lzzaNcHwtl7x8YGpmW055S4VvIWh75+kJRp21AmUGOoTqQwX
25iF1ULXRvh+hKXs8F5pVQLMvls1N7fcwK0ACHgOizFFnUSTEhjL6Wm5/GfL3vtMl6O+5jkfZ8OB
X4j0rqSJvCtVsT36Y1BRCV6l4YH4JoJ9amrHBbHMlernSZvooWAnnt5t4jDaB2+pL4OZisfaqVZ5
+6MImwSrShn7fOLkUhk0IV0htqmxghlI1macJAUZYZUetlMQbbdvsmXJq6W8WJHkwUKeso/z5Agl
i+hTq3WGfk0hLO2rUJVY4GzmjdWXO9I1bOxgLuvtBFh7+FfSeel3GRV4b0juKqng/f5YiMHyFbb/
r9iooy675PPKTWQn8g5gZgB3PowUa8IgHBPsHdFCeIk2l69u5ZDZup2u2NToiyYkm8rAlwWpjSsP
5ynt0DCNdR1Qtg9Ahna2bKlhemM1wcHG+cRI8GAxyvH2CAmccA4FU+5LI1kBdNxETlcg7vnhzvQI
9HMomAoLBJxJpE54fCAuQlyg/CKR2BiD3QY7YtEdMaDQzmAGX/o+fhV5O9pvu/oLlNammT1PcVg7
RGx70UzxCNgQvTTeTWyKDLMjpTVAAH84RugCTx80ZkAjHU4n0KkVQDNkXFmDdZNP9RpPLCmjXRnL
RWCY4wOOxqwU+NV2Qa1+4SPmY6LktjKws2uZDjEQQNUF77R+CV2GIz6kisTim9mkhjCCfzFF3nu4
iMfgE6g9fTL92pT4cTwr2XujgaHnA2AVLSACSUjmHeErHnRK/DDMgQoWQ1+LKmUKyxtb80F5rHtN
vWg9zL1lgk9hZsi1EIqk/nVrQK14sQ7x0PAcKYiCCOEimi3RXJm8ZLQi513vjmpeggqcz85Gxv+x
NV82Ki3VbEKbo7fWvny2xPl8vJS4hCicP+XnM5fJw4CP4KC+zxCGfPNk1sWb+gjXYYae21W8Bg7Y
rZ95ls/OK9Po5Wh+S7ysEW9OWZv5vWTgM9ACZUIFYk4oejlphRR8Uyjoa41xTggvMC8UgMxvDK+T
ACQD9S9C93JGR4cTodkWxuHm78SIhFZ7pbxh8YyzEnBwoRup3btxmob6kmSAJA7rbBKbTpQ1+cXe
NTvlhzF/MSpfoy2IxhWCJkdICe+dhfRRBvnwpVd+1b7K+Ee2Sw52wkE0FwlIdOliS5DD6cDVVD1Q
EpOyOsgG+frMpoSSrpobueiPjxoNHolpDsnl3ejvkWXMNgGJP2LkvQSKSdiD/efU8S8y64Zso0H1
0FgJR59+fbY4QAYZg0ekJTRhJMPmZRYTJLMWsupmy1Embdc4hTS4ww50fQY6w2Z+hw25x1Jw2B8B
54Nfr29wmpk1f8/ncQM5v5PJPVL5pC4OiNgpmyA1rwsRBAnWlDvJj4NhEGFgy0i0kknactvtRY31
L2P8YWnOBy75w3LCHk8WEMBM4NZXEeMSrpwFDr+j5OF9Tb/amcDwFM+Ryj9z2eYW0sxy1pYoDtVQ
JZeyjnSKMdOA2gwstekegH0h0USxGTGauFM/7GGew+vMsMVCoxozCvK8gG0g7iI3VPhV8inDFAtl
EUH0A+oY3x+L1rMfp3C6ecEvITKrgjlhFXdTd2D/QmUGbsjqk2RmHTWqo/RJS31RydKcG9oquQfJ
2Fh41PGcg7fqFroD9PuF9ez8TEaWe5Dwz8Y94QqEyg+VGpe8fZQBF7IocovhJnfb/XUNL5FhCMT3
5kW96JfRR9SVCk/hNZ1jHkr7vwXKovFEq7dZsAHQVueNjtFGESOtPEwFT7CswnfNHazkWXDPw9CT
25YT0JWlE+zbr/mcg/Eg2NpxfUcsRvfz2Bca+u/zw1IEULz9PvdCUxu3XudCtecy18Y77k/mUOuZ
vmdtGe/QtbEd+JhMiqp6NVy1e6wildUEoUQXxoOKALJXS9iBAAXi6KGH8SQnpJyWrS90XTNLXEtw
9XRtG8/LfJQwquncj5PhikxKz9YFrV//GbyC+bOO8C4mt1s9XuPnZToPoSajSgLr8vg0UiXgB+Tp
4ktbS9iDSKucJU8PUCDL2tYSfiqWUtYdXfDsBNv04zV+t2ttr5c2/+nZBO0YJBtCXt92VOQSi+X3
pBGZZrSBhQVJaudPnogtsEJWsasWAJ2xJDvngYE15LLinu+OVrqiv/OVaJj8fEXy7ls2PLQy+TAY
w5GM/WwtvdFaehis0S5OZnD8fgBTEcP7qMfCfedlsyygaB3AcezRzcRIbX6DFMljoEBQS0adRkq6
o6csAjd7cVCTK+HfBhx/R3hHFtSPZuR4PnJgLN+9bbr8zs5tkbCA8u6JPGNRnOzFvv7cDkgLOqiq
cV6bWfN5aCISND92UTjg5QeWqY1VJHgol22QS2iKTFVc8kGXCJv2f60ME+Q+gbbY9bL8JK9klAy3
0M7ED+OXL/fgVGmCZJ9wLLcSHPbZKtKYpJTOOaBzf5BSYXSgq99+te4QkQChK7Bi0aNN7I+KhESR
JrranfRj0sm+JBzMEJFouCFfOs9VYGbUCPMXdDiJj3FH7E8fewkox0SnEbXG6qgR8o3breMhYSMY
jn/igQupZopeCMM4MFksG3EbG4EWhQEF0MMrbUuIWXEdOor9I5h2Nbv0VXeCiMDuDnzLQexA0IsA
O0bjfZbOIH9FrOyo0Uqwf8C++Fz2q9vocHZKWfQOj5UYvRxvzI+uag+Aaf//JRRHh50rlcqtmw6M
R+6fQ4MAwtnNoAscfHrX1Nqx+HEmE772c8DQnwtz7T1zz4hvOJ5npmSShEV+1fBAEnNZM27rSfZs
Li/HOoNU4n8zA0XdlUNSj2AGzRaGDuz84evC1o/WjN49sLKZkoSfPz0jcaQgmyZRjFOJoSkTXZD2
CwaeZ7L+Al67cu0FS7gU20ZHcVAak12jv4T4M5Rk+PmUy+XpwqshbQJuZrhyBX88naAml2h2bBJg
8HWfkx4GiEY2HIaTXX6d7UDlGU6LLUoGaxeIav5k1tas79ooj+XyFhBPk+LXqg+AFxn9BlXK6/2i
9GtikUgcFAIC5+C6WKwyyGxoGPLp8Wl5/+6L7lP5adHhvQ4BLkbSjU2b/AwjJT7OtbIpFTfCSzJk
dkBlcOEXcpDj26ol443n3CqrNQrv7MnoL2XkjLWGtq9Z+7lDVfBO2p6oYKc+OBSjHbVTRvDlAht/
8zxmJPah5hHO8dTcvgv07wtaN6vIYgBcZmAXUddaSYRHGnIftkep4ojySntZdM8edU9JgFP9HmVe
+vNTryuBdBmM/MOykxOrUuI7917cDlHskhLM5BCDj7PoBq7KpzSEd5FLtbpwMM4Md7vx8BI+hT0q
ivIAKDnwNHD3tkg08lsWT7A0SWzrgOauGl3TZuLWrDwS3umq+JYEb+Xdz0HT0pwx6TXZKBv3bLA8
93iIsfO0kg600i/3oJ0hVq+AMws1uqQRamcX1kMJF3uCTdSA6w/DCXfu8thxVvY9J4LI0/oU86ed
eNUasMfOU6UsKvnpRP1zfZb4lFVOhYLPjRc4WzAm1H/V03dDF+PmbsbkGTksxcHcZsg7akLrezWw
eFdqAfpSOIb3r7Wx+iy0GYdTw5fpRH9BKJFw4h7ZyGgmfniHbQ4hzlH+fWmN97+FJZ6jLUuo36RK
gmAT4MtMKwXoH450s2SbTUoXsF7dNwmW9+UvXny9KgJOK3VzmR7V67a/H12Tdv/qWVHNfcyKAsyj
mA6Y+6Ijj4K4JC42it7Wfe0aNtYV/YxssWx0HJLnmfk3jkq4KILJ56LH1YUL+Y+tPwbIjMxtn3rH
OBvg7U1H11RWxakt2qdSKGHhnp3yHerxXcxoEUtD0PNQsMNkUyQEuU7G2WdVAxb4btNQlWAbhxZv
HuxIQPmt79Df/cv2aXswzuWsshKUOus0O7gdzS8n0vGZ1IyKHfH/OKv7ziLw7qmmu271P16Eh4nJ
RTaJmenWVfz8vxQVTabHvWe7n/dLZJeb/yjabFMcVQ1hE3qi1IScKfpjN6LF9/uCYMQJgaXYZHJh
kBQFgqBqG+4FxRETi7u5UYWbi+sSsk+GHMqejgYmo5t0gdeq4/89GpkMbgEkD7zVhf1JMQdlDY2/
jEWzNh8hPXJ0FrWwXRw3iOkCAhi73oHvyStY2HJr1CaHYhHcpEPZagrwaGwPUUGANVdPDmg4mLVu
GbuYSSFKT/p8EEDbMIPj6x+CloFYSgrycyR3st+vmA0gdulL7zaqgPjKbkZBGo/KoDVhqN03bvif
duyPwTiKeAwHyXhq66ZtJBR8PVVpjG7Y51OzYb2c63wbdEwFxvhXSkCvCfqfJFyIBzQ1RIHm0fnO
ESLr+pa8gm1LNhvz2lWROzDqU7SJB6CBjaXbqvtAMfvDUGDqKIwv2aMA54ixq2/W2AiMSNNKhg78
4u2W89ahvcBXVkMU7/xIzJ6rswemYErDUgwgPBS3UctH9ls1B/aGc8FCvbQjp8EwYV6zaxQTdQdT
BV32bIKSYZIJc1AwtIvlu2/WO92s+Nvp95053u8RjWvIb7xUFeKUOFB8qkgb6JHFY8BmLIU6m86/
3nfLMP32ZhUIAJKjpb9FHtPN9Vl/aUzZaDGimzXP+nZqx88rv29yTivKQi6cZRACLvTC4q9j9tn3
iNmhxEU1Qibk4Tm2WnoOkQAGRvXAt8uLcGSkYYxGY4kiyOfU+HCn9lf8Jlij/Kxif3VOgYvxxp5F
FbYrNwhT2NkNqoxB9bVppx7Y1a6ellFuNgzaPN6pfdgbYrQcs8J8AdZVYy+ijncS12NGaIoHZGhM
2aXEqFJvuvjZK+r3znot7QNdwNpisx7PiNCaNbTt+F04yhDBgujLPNwq5tCSrwVUu+bQpRm2l1iD
3zSVp22zYrIK30eVHrF4o1aMP2juYAFu6uAkV8CZ0oW+10QjYaWgHWUxmmAB8SFgiNYX3PHzjMxA
YUtEzk5aK5T+7YZ2MaFkIqKurLjGfJek1K4bCdxNAKAi0+u0wZUbCGD1Skt8DejxPOqK1Scp8Psx
1++R/SIgJhZftv8KeeLk2n5u27KwFe46LcIZib+Z+iWxY+LvbUcRIPbAqtCa+8URGatn/o9jpwRj
68NuqZ1ofIsDWe1H2EsGm21OxJlcSkuRvJifCjRpMtL6qigUoE7tjb056wDMhhtAXf4no54iJuY3
xWiSgRVmAIer3+mpNkuRhf6ztixxHqCAn9pSV7c2H1PXAgHf7yd2YR/wPPXE838aAABRDv37uJqZ
O5DLzqGr7GGZg7mKh9ddPWv/O4xcEbe3j7ejdw1Xazef4PPyJGxGVCwCNLvJ+1SFtgfLyMCLQofc
PoBHuj5O5Bj6QaZ5jF5lIwsvUsCG/F45Yo34mxWzMLC1mdlR7OBmOUDLK4qWgkTSQr0PtjwxC6b0
B2UKJutNalbLhz27NUQILAxfmxnhmEPSUHx6YN6EPaOwe0VUH5JJw2FFQlNT0q6N/JRm/yLaOprM
kJXAGHT+5rSej2TUQOmO/3WcrFC/6Q4MEWrqUnLHsdIc5XXfMfv5+05l/xrFnJBKQD4yVLfFEyBU
E0lriw+GBfegjgh2deobpGMAgVXksLy4jOob/q1yQCokk/nxTjDVK766Slg4bdEws+QFzjmkr0dq
IGqNMhOQhBbQ9OAseW40nb0BNtS5ZHx+yiS1d4/eRPLxQs4HgbEEJT/hcuwZ9mscpegkHethPpaS
DsDQRy+9GdR2gnWOE8VOsgbGB08jhvZIzm5Hu5OndnFbpAnl+LDyPLAF3+qN/mVwtaZ/kP4DYySa
9JU8vnFsSoQ16wLOzhIXN+SoT4Fx3nVO+Vyg+y4x6J7AzOtymOk1fDx4Uwn1ViYMF9mhd8WU9Va0
tMlzdNP5MaeQ13ECm0kSlyafqgcwbPX+I8mfWUKtGWG/gx96fyHYRqnPJCvPfo9OPTVIDkjJQSjK
b8eFfCMo3euyrW6W1bZSqbIy7kBhdxDuYYbFal7aiJg8Y4pVRCYN38Bc5KI937tYmqDrBsXy2/Ls
NJ3EG2Vjwwepyp7JPRzHYtdBR1nBhLHfvq5EkXL2pQA1p/P1Hf+mPZHKrHGeAG42SuUKaT4HO0OB
1gduJuM2pisxYtbtBXZRFYFpPow3bWFrugeABfGAorRKrAOseyP8/0fetunChoLUkWU3ShkKL3n1
UipbLxZWytJfOEqjQOr6E7yicrSt0dmxgwCHp11Qm7pz2t1HacajGVRFiLImPzau4VXDGj1syZOa
RwuyNMJQEIRI7E3XThBjl5iW2Qb7UQ7m9yyfL/5aZu6Sk8aYhU4U6Vcue/OpmKFO3cgDD6DUFIXs
yUxWf0IIVd6LTgeVftrDPyKA1YAQ0BqfBrjrL78Zx1RXU7ozofXznDvSpY+oIhSSDmuIbXoQ9FTn
mDvgKAEgOa0IcauG8jW7Pnja6thZ5n9pmQ+IBrD+Tox58aRhUQe7LeV5D/W/3ExLdGW/F3XGTFxD
QIg6TqnS4bT/B2KoDS/3uJFclsO//cRetRj1V/7zLm3qpAv5h2HzjcqUj9mPR8Y9tjSgsqUG+sea
qjPWxolgnoY9IOqsWGZZie/9VmmHWpVlqD8Nrfv5Yjzco+a3zIdXhG4A6MGwj7l++6P4WWazWOWQ
EZUqyd/IAedy71QMtn9VZ1bmW5u5MjVMQD0cO2HzT33Tppuq0iu0SP+6+KJgswJCuhQY4PmB/43p
QkYzRdSpksc3Jb9hhSe+FG0hzx6EBdfVQQDlkhX5E5xzvKlXZDnn+EUqIxc9PdvnnrNILs7KYTDJ
rlPRE0EPo4q8F6e6UB24vQI/7+2rXnk9F6aHKVoCFquLu3bCQrCfCpXmk6z7XAJWpj5Od3wxszDB
GWG8zTVDek6clD0+DyW+FLil51oqpga6FE8IqnVX/7Mqjoa6ad7tXEdYEX3abEMDeJJhLujN0GWa
XeMexs5nofOFq+8kBdqIx/lwpuKDz3YzsvsZ+VPhqGxyKq0CfvNDpJns3t+DZABoku/VUwtcA6rw
avlCulmHqkslbXHBbgf2OGu8+FoXW4iyYB30RTYdM1+/8EdDVfvEH+tnxXMGNHHQdKl5/TzytQuR
WpWTXR66MDraXrVSq/JqHxE5OObHG99ZExL4nZLQ9tOexFYUdbZhrXGSKeIg1q8jpgqpuVpAmwLp
Cv/bcD5TaXPribDSKWJ+ux0agGJJrpRN/e2okkzodivfEFLCHU6YcjMTaVNhlzEwbL2TmxQwENso
C6vYzFpc/p71twsikECBSRNJFX6V4eCiJs23qWmYJaPLH7IPqbwlY9q9IPeiCJK+DZahidcA0VYh
fR3uXM3mI7LAF78C8CDYBkkYLy6wnCkayM2DLby4Dto7itr7Swt7B80KoYZy3tjcPrtfFeN25cxa
brVdu656g47yzojCC6cpAJqVxJgSFWSJbSM/7Wc3mo5FKgvh+naXy98pB2XglcV6tHPefYodSKj4
ealy/vjv2aWN6Y7jFo6Jlt/HEkCKLE+oL3c4LbPwzipwarmtlPH8/1jjCbi5c8bzgdpdWdLiNJWn
ICvB7tVlZy9MLP+cqIkz+IPgHq1KTnT/AeCzTcxREeuz3Z3QOt1yHWeGw6Xb6HBmCVgTUNi0jnHs
OpAqkP6hUdqjhGuuIRpj4QXyLs/lFZKvj8tPdJSM4xrJLpbN3E65kBCmDA0Er3aQnVX0Inub09yA
Ya+vz2XRseQryVWHjcz2qhdhbA3euSbOYR7Lv3w13WVuIaKIzMimNCO1j4ZBhcuyVW3kwPqID4TC
Km0E6KYNwLP1zAEjBfiIxKMeXDjIRHqf1BgAnOod0AW6OmoVy150Vc+TOTUEqmGX8OkHFrO80aLm
MUuN0j/4elyOriydLNK/z8s21M3XJCLh5bjkol+GcVveqb7uZDYPFgqZ91TuUt/CnPrFbFTosyD3
oVYxmtur002DaBVtcnXzcd02erdqzLou3svCiMOYkYA+LaCZYCmYLHObj6i0VFxX6FnjMTKU1uYp
cC7HGZ/WJo8VHoOSK8MNFsI274ojKb58moenrNP2B7b/4qk6m/q4ehFQtaoi7cgH85JiUqKzu690
rqOZeEFdl7HdVDL5DGeYMwH0CEqqjkH+odzq5gI6vovZ30PqEl+vQfSl7nHwJiNQKUSziCjH7LJ/
8eOu9HCj9vZDvPciBjSbbz5UI9twFJHW5VXgepS+Rfi2zccEDgkNQKmgbQigJCiHivMYOV+P530n
ZVY31ksdgPIinAAyyyXwfAXA9vbTOLGgEBYP6FPDbMKxYVljwIDBGRC46zkhrb/X30vcZmx0Pjfo
LvgLcsyRetH3liAsEgVI9SS32RsBTWMBz2e8a/se856rTmLrgVqNcSx71UyaoS9HMBC9SivupXsp
kt/vhWhk/mOkwYmRF3G+NBV4Hfj5fnsLpCIzO/3FuMkURsyINj8pTXbYiSIovPLTMKcINaPXU5tD
xG8eVdmJchEJIXeX27n4bL4Z5anC8g/8rKoyOM7n4yj2LimuAU3dfXKpGV3teBzNui8nbC77GAl2
2z+Jnrre7bJm310Y6VF4+jk8qhrk2tmqAngi/P+0V6+Nk+oJgdHWgufPwdAFAxHV4BNo6g1kmi+c
f7T7u56WkifNXrB1zk8GtYUkaCQtZTgIVb0GWMRXCISrUzCTRsIS3fxBpEl9DGHdGbAav8VdNau3
Pl0VwPhL6fhSNR5/UEF+mZKuAxupR9yHsaAzZrTPEWie2Lq/RKSxTTlYaMCVlnoCXOf9K7miIBz3
R87wPHNmO70R7bChZgsIhpvFFdBMPoCFKSVrl3pLCsYubZrcGP4Kkgbr6FP4EAQHJlsZC+HLSPBu
EpTrdmXjrPMaNCxvZy9cNTORmGVO3T9nr1S5HqcSD8O7yqkDG8CosEloIa5rVBiMC2kIwFT3rTmL
64aX+hfEEgd7TFlcIlN+/3A8J0F6DYmC6tMEQnxg6aKgK7s0xCPCBiG2wpFJT3fmW6r3mtJ94gXj
Q4RCWgL+Ce4G0fney0pneKbn1TsHflK61t4O/ce0p+L1PdNKzajxgE0neb+stYvcEN2gRqRsjt8l
LsikHzc6+vTJZo0p0W5E1PS9GlbvaztnCq7KXa8DWDXLWdVDcbA8zwLI6dIkqUd18yJG29HW+6Xq
Q2wT4m4quvvH60iaPwig2CqDHP5bQPktV4Y6nw1n6j8ZK/S6f/NYkQRRPyWRtOb4bJ8YK8Q4WRXJ
vz+fK96iPIy4BT8Hc/+4TCbHtKq6rLy367lcrPITnhwNcKTTS3hIxPpvGTxNGlegMZVGGOQv3D0J
fPFeM5IWWNET5kDBY92sBxdWNtNBY2AF5b1/ySPR3/2Iqza4GH0FYZCdMw30VfvNNFfrxpFSeA0Q
rPfFBmruHAlIqUycE5gl1qY3aNmRBQs4OiH4NB/g0epcwgEW5LbsnKu9OUI37DUA0gVdZyI/V+H7
p64yESWIcrOodn1IuWE208MPwdThSSyOwsZOi5u+TbXPjG3A6StTx+7Nml5gsK5pnC4kwqbaRbTM
66YXQro6cA3oW4AL+q9MRfH54IYmTExfYNt/+MMGEC74AS/pWQOG7pqFFVIgjsnKysxPA5G78SAn
bGkfytNAPTqjAY03s8r4SEx9yRuWk5uzumHAQ4m4/iXfKqdYHiMufpHlKNsDRfOBjRn56k1oofBB
rUOez3lsb+fiWe5N9LWPTgzPT5ubcLJASJSc6MF9O3SgNSXUCxuaOr7n2hExnW3IFSc8pAVBRsQw
1V8vcSTD3e7vhUXa0nUJlBPpKFod7jMcA3pgrLgyUscNIg/vomp0tSE/ufqjFmeNzcyB7sCfkkGH
yH4YdVHPQArj+Zmg1/ks8ikysjht7P64+JsE967TLduosMlx2eu4kv+/7vTtOfRQU6ipBXO+FElh
Uy5sM7S7gPabfFNhKM8r+rEwl3AbvGUDXN/1gt9kZ9EgyrfwVzcCprZ1Y7OHqszZYKo/WeInpauX
LI0Rep58lRIHUDrlw7KH6O/Vn/hFn1y03Ctj/1W2njfgjUAsSvQXZHXgWHQ598rKPWR5hVRTL6pu
GRujkYAJGDhOiKU+nmZKmQfs4A8cDnWngbC1POFeVubyAeS9yLDYUiavXVK59P8kZopqKJNPxtqh
mR2ypF1KRFsuyPODK8m737+cBw+gSP1joyjVRvAzgS5GhpELmPPIuI+pASQqMs2E4uZEw/r+fxa/
H4tt7iCOiuYuizwcwz6n8fIEWznTINn88KxGYYsNQrtNJvm7o/Y5Fmu9lX56ZvJgTXDYgCzHJrJf
jTvosPtL+z9KowRE+accDSjA2pd9zmwOoxJYHL1fZJQgEZ71Dd9D6FhLz7p6GOG+MDENfeCh2gCT
DQXuFQk3cReRM8qxm83swNyoWDwWJDwslIFX4qYyXCnIZ7mlRCUVMTAEhQOqCc9OOXB/pY0HpThF
a+8ZVMi1+1ZzxBD7oSOKeUfbveAxzMo4JR9DDcgonJb3FYPTroE30rOhC1UoHcMIqO/rAjhOXhmV
PkCo0p/ssia+xlfAEPY0eRvp7dVTChm4Zx5dXJv9M8EhjYiItujC4eu4IjntMWKv+bMAhLukIq/T
CtFed1WGxPZwBpQjVR/1L2UNnkiTCYNh7FYFZ9Ou10zgCRee1iQNNlbca+VEvzvVr5dgWQojYZ37
z+ICNi8wAci3JrOeNMyHDhJGVEQFH1bE3F7ydcPDngp2TCsulhLykWfpvIh1TbIZFlQYj+jRveis
7vjoFKwT+dNc/Ov4VtUzyHCKz+j/a7jHNbh86KBZ4O7Q4+5Nq+mR/jCyC4wijLsSHs/JXWB8Fnb/
Aqmq7kBs8KJsO2NnT6Kxd1vUovwx6Df9v9KpmFWTwBdD1Kwx4EGDKBG5R20Ip2I0RcEnQcrU5Klo
9sCjntYw7vg/nLeDJgYtIR5WZf1pcZ8gKcRcW+UfA8O45qr3RUcD0uSH96zovp+zhJ4TPSGSHGIM
MqNTSco7Dj90tXrMfQ5EkGDmDSSs7cteq0nukPVcZNWPM6yQZ4Q3J/2Squ0+7/zX3FY9kMuG63QB
0gAyd5hfFUkIKgOFH8nQD+W67v1/359iCynIRVq48kQCPWW5Yk32owc50Ws8P7KQgSGEgrAo+3eM
qz3bPS9lo1CLxbACSOsTtEqArguD+owatUTUNj9WhNqp7vQ3gCCMh/KeysCXiy0Ob2V1wQKIyMG4
mMagyY3TEWAv0vtSL4B/0aJ/zvbSglxw8v2Ii/nu0H/+YoSxAWFVUu4ytgE5yWjoUJHo0fuSbvjo
04OsyxW8HPfgJw2F4jcN0MRZk/MiWs0TF+hY6keqY/NwZ6LUsjOloj2OlFpKGi6kF6KYMFftXn2j
DNZMNO8Z33oE2D0H06P4JuyJjPe5kwcqFAvvbpPXA9BrKuK30xySvHMXDQf55/nPuGxX8VTuYKk5
rLsBI0aH3C6FIyWgkmofzu9+Jr2c7K7mk3sdXGGQRa6XeUiO2y3NTZazCGAXlDJ0J3kPhRBoSVnS
5L0a5wWmnQG+dmWvjn9CXQbIwXopHgeAnps8Lvn0pzoi9C5ziBID1qNdEb683cpdlYgqcjHKdDpr
daYvgSOK72nm8X6iSOi9GmvxqsynutAVTy0j7Aa82oYQ2M2j+M+3ux5GDvsMx3s0DycUgIqT2/EN
F+7hV5Zj7bxbbla2cHoRqcZgeU6nAr7s54LCVgHxyruOWc8exwmP2NqA7M2Ps2K7IUWO4Q0ADHTQ
ZbBDSfS4RW6mm8e2CMj/SgjKy/QKqEooXC9ygFVoqrcgHTx7eIV8ZzjG5zoteqUt2xOYGRYgfPpA
V8vyKNP32uQY407X3ehY5099e/xH7ccGfm8yVCFphB2RgN7pI6aLsQFlWMZP2zQ3r5+ineFqPAwS
y3nnUGQKXDRmNGIZRLGfclRX+AWS+eooshmSVr5668G7lfyLSkZb1YpZLuFALUOFsQw8RXPffNPQ
62rWAItqIk21+D881gvyDuEZU2rM0jK82jNutoK1e/Cw45xc5QbCt6g/8qRAxwyqMSEDDAEqSvu5
/sT4POa8FXA5z21x6+V4oU3DkqVlX+yYAf/uklZyHojZyKBb1OnMp5FpB5ALPS774CNB/bexJj/p
xTLgzAC9+FCGe9Yk4zSw4bnwW+WhaHhDeHGlDu+c9IQqpfHzb0+WKzfU0ALjzf8MGlMkiIt4Z1fW
VguMcT/1kczRDNI3+bnkEqad9uNt8i/jYJPC+GITMSQXcsVRdFP+vOCRXhfyPdFeTZq7PT4Y1tU6
TvlQsNkou0McnLslyJSJmN5NKmSEro29RO/I8XNqUGJkG3q9nMdB4MzsFZS3z532ygXGaKjxx4mn
I6K+FIieb1d/jAXfsjmQiXnBR2ZCMdKZJHhEQktjJheSmVMTYvSY4kbQvj4X6uDAm1QOOlSa+Nar
gy+8aVaosY0bB6+IkQzusfw11jaXEHrjOmYnm/itpfooDIxSvjO+Z/lgNqP4tHCKqKitKPM1/nXl
flTfoJMWVxWsBeMFcgyTkB7F+XevWdkdqFEU7UaGtd4ldRx6YDgpl8S3NK/RKWPEGKBeHrsobbKs
TpunBaUKqqwH6JNwCcfD2fNkSSCP9IHrlcfVZw0zAy5Y/aM89HjjW/wIPMrbRARwYQSPFl9hCH1K
LslQluhW8k2grgIEJzWWL60jMkWOHqA3Ml/qMppNXT0iLaqYJJaa1TaNxTuJyUUSBtm102U+msDQ
zWCwRk7PXbARsvwtLUWOeALoS/eJc9LQiF5acGEL0DNUOlAMZGyS4PahfvpS27BcAW7umu+QmH2l
CZ6ZH8QCmcLgsXxcFYDssU/XTQvqGmdRwDPv0pNwMf71/5SD1rccgMHYhZDxd6mAtTVr9rRu0nRo
mQrkPrqmiXuXlX9aZtaCuywlORjhBXtj1VCAU5a/WR4MykSBsRm6xAfMeRNLWev2cRI5TxBVUBLa
sjussxiiqRZ8x/O2yhTkyAWIHus9Ib3QtS0gDAKlLT3GFw7a5CoRdEey+l58aCy1JDqUBi6L5uPZ
O5QojNOIRfttdjSDdUqJKVA89h3vEg68JtqnLakYYul4zE6mj5eS+dCjqRItt3ev23n3gqCXZEeE
ywzGb9eqZOLOdgWyHPyYbRig8KZQBXFNWp9h7wVcjift0wBBdaZWq+El0U83ubzYTPwIMgcpLuPi
MMIeciq0e/wIs3B9yxywRsEkxJL80d4I27TMgLejCBr/kf0u1p0ykA0bLy4TdzHxQAxDHrmFOkgq
bXqGTHYvnq8qdAtsiIVRsMAkJoNLSIZM/cW6Q4MIrE1GWfMuwED+ZjtXinCMVTVrABi+HI8laFvH
BCMfgTH555iHOQWd0ruC/OCvvrq5nemh66iI9t3YyimG6RyEq1//eW9vE18jZuegB+M4j4vXXYu6
b8MIm+IJzZYmt/iNcenVMm2v3nZAgpGfQWj8p3oA8Pw4qUzV64+2L+HcnOMU/5kIuxvxijRZIfau
azLyjAziMawnvTNA7qGznqpkuwOjJIvWYZlrSRkfl8QIaDxztSSQ6ehrPXKTbOIwBRO8CF+8eMeQ
BSFNXlzHNRpOPsuBEE+t3+j+Q6zT01z9Q5vQe/8XO/MWgolQ9ILnmDN1ucDG3bzytWl888k1J43U
UHNzz+AoAQRbXwHUMMQ8ipuAmP9CXR7Jrklw3KrrqMowhHCv/4NhRcmnco34IEYqRpogMb3tGBcG
/+RfB9y6Td1tTZuGOy6RLojmZH6LftwscvzGwOpk4yZEjF06JLXja021yIlzRO+9+Rnt7UJ+GHG7
yWQHz8g0YInJCLLmjciahfMFck7jHQgdIBPy48mGYcqXD788XcOvWKg7DBzPS0bQv89v8O98PQHF
btdj71KvGQJ5FXWRtI1LiD3edSVzdmcBQxp8ymXP0omEGRAzYS4HCY00bdowFLkB8nN5b3X5KYfo
BrZn7axOvr8LHZwcjEIxcgkg3R6fgwMaZbTv7iSiChJvk5y7U40qoplbq+nH9t9lC1GGgGWeX64Z
s4ljb3gkPovjzVigckTn3vlo1vqJKo6NIPq3mRll/G3+T4NKLw7027nz+IXB5jRD/Mw4hxr5oUBY
X5YS7HBAUk4QovG+cKsNqHz8iDKc4mk2hYzPbxNkp0nrtqKXwt29yFQrQOOsi2AelJZQ1jufgrtg
a+DHmKmRQsAFDjIGIt/Mh97WMxn6A5dM3ZKE14oXHygtsenePUMqO7wT9jykxz6hwnlKW8N9MkYG
RdphReQMBFzIF8/YCfkgfBry7AkEK44L6dwzYi2qDyEgULazTN9J95l6/1i6PDvhqU2pyuW1AtbA
bsvlTqh+6ykxVDpOOmcz0i5+/Ci43zaW90eTcR/m6xqKlKeWfv50aqoJ1JnLr1cipBlxKcE/h4z8
taLueJR3eBGE6FkUMDzj4JbfDA+EHDIHrXMiqKFqsfRK/r9K3cMpGDQTiKFkxX3FqtFIJK8zKFjx
zo/nbU49xJLrceNcduR/iciJL8PkxpZzXp6P5E6wmKjN+FS5rNrhCblVY1bkGtTY++nV9oV28wWp
0GhlnRxoPE2O/AH4ty7XgtsCc/bnDGOpsQFKJeFzKPV8eI6eFfmx70T2Z8qCUirYjXAwE9rbjVTQ
8JCPCEKaQooiVn2+FxDbCkjYZyzAZvxaU2zIsLOiQBolPHmp1zWYfNwtWnANpw6/z9plTXlgM+hK
bzsjCsQbnkMmQfG6ea/Ao4FmbgvKyXQlKhN+AtnBcSfR9B/61M7Xgt9EOmQbx/TdwaQrQ6Eh9pyQ
t1LTACtVZhEDz3xfvO9onVUzanVEdvdjky2zr+4sn1a2hHclPHOtS9m7zkbDpkyATw5yUASPSZaU
RpixhOBmqLsRAtFsil5JOsWRl6j0JzoqlTlTcFpitvuiuy62sNvG2n1UCB+uTjdngq0eDNjY2V8H
2MdWLpU6IMk1cxtEz8EnHgf7cELWedB8hNdTsRa67jn1Ancz0sLgGJkZmwJ2vzlZMQwsLgM5aPnL
KjaNR9a8zhYRrQtedQaqekOseGo5MpJfrA6Gv2QLzjojfn5gofzUjjC4zGghz/Nz83spXXTmzb4w
hf3YH1NKqzOg6Q+S8Un+uZGkeVX278uohXagVVp16DrvcN2QgyPJAC2qxYHb1O3ztSVoI2A+B24B
tNUCSSfK373MDy3an1cIEAPWyHvnVIVX5eXt99K4WVq7kOBXfLu1XINil/EBlkrfcOJr4yeSWv9b
5S+AghXwwC6OnpJkPHM+lu+zOUelu3zGvBPEGwVSo0Xi7kVSYlb6i67EgRzLYnbOsQAuee2DYL1u
J6zEajY/XvojFQPrSSoBYW4J3bVTEecACF8dYngMsmCzHMlCjqulwYggB7aybH8ahBPJ08iC/htD
dTqIWv/SlJUgNEVQxwR5GStzDD6cH1iMvLmlOwjV+KAxFT9zYYV85is1qI9uwSa3Z6KGspo60R39
cPi/w9btUatugxMLkfqumYE8ko6TUGYxhBVp91DgEDZa6c69A2beiv/RxsBrkAyHdAafIjuKJyCd
3/MvT4QyR5Ow/G2szq1SPYbPENJ+bIc7VetvUmR1s0lx0yZMuISM4ykGsZDQSod7SVD2I3upl72j
XSLxCrsWUCfB2LxvqHEwnLkRMFYT4lKA01ZZJKAz9WSvsUhc1gxTsfotSjIuEmNhFotbsQmDK1lQ
RpFB34s5oml/Lq1Hp1B9OMuv5wb6HZ3SWFfb0ZCNNgpcN1AxNdehrPKJ5G3pwe07dM8etQADRjCi
xbLvowG+2gBAfeNzicZvKeBMWatzjXtlmDrc9cXxfzhzi41KbvMfNO+VdhwBvgT/U3ibOx/tNQe7
xpsUH9c+Mp0KQvPUQ6l+RYxXzEvnFV6CDnqozRqPh/FN7vCq5s7vKYNo+rSVTHyZN8k3n42zpsbJ
O39dYJdGi1MYuFq8u4weGzkYBOfzFET+2v4/AnWJH4e3ze1G7QWPxYD2WwdpKPghahI0MOqDcIj2
l3umiPWxzd1hlESd2dQTUvu5HA45fws1Oo0G/YLkdbEYfAxqmQCWyyvBp4TM8376zHVB5hoTDWMU
pw366qQUqI6XezTpGFhhQkNjhy+D0yi6cfJVGl3y7nQX3CQZk+laX5LtQ5+5To8+Cy2XK4zlTtid
1OAxDIAnMdESlPGU4SIwmAgQGbkzGBPfO2DE88s51FlwSo5A78pQvCpd8ZJhc+JOzqHZHzdXEos9
pypQ92DZkHBDABsOc90LV68rnLYZaiJ6XuZdVIcxEn6hYFnESYMzpa+jq5PPW1hJQWwlfTvN08Zf
ykWMnl1E5MFTxTqdclilNZxE5IibwTS9JDnGS9zNiuWQn7VNl27NTPsuKgdE7bnKTqxDoHTeBlW5
ahDCZhageKw9tzSohFfW1VcemPSfu8/haTyzOf4nCZEVwcKzdcSvRSfhOoK+uy//gFEwOVaALyxA
R9zzgDc/eUBBOdCtZQyTg8VupPhB9kskJqacja+1xhoKMhAqaqoE0fm75YxbntxWUiuf9ZyWle7S
pd9DeWxaNZq9gFK+OImmXgIUhVKqow0f8tFa40gOUXTzEIJ3Q1es2PU2gBw5o+m3ZjQB9lta8Ijq
L2i/nDnLihKvzeXErmqtPssjG72kZT6ZwX0QvZhhlMG/aLqazASnvieRq4gnLdusVg0Q0aLU4460
m/ErKWqp2DqxjQtDjDXzw9PH+VGLlYPvgVZ7GoD21LkH3eD66LJ88H4e72xptFaOYk0VHYRC99yX
pILbrCC7wqYvvayo+Rx7jQIrB2Qbj6/ztH2PEfgrM3hD31i/qhvafqfbz7bcDmn74k73qakGsx2D
vnOH24sT9dCgaS9eipqxbEHWDh0pyDwORtTHTc38RavwbcGi03Lp6gD3aWs3Ij/NUHn/TBdRgaPi
r1cB1L25gSWb87SXe52jG7hgBvnl9WqzMCc7dH4u6Cj+bXOte4o61hBRHWlORN2dRQILx1A6MEbu
wQ5uEDwkleDmxXDz4OFT+PJSeVP+SaE3TE7YASLvHparznFHfaqLPv0wbv4M047rFt9lstJ5KW3N
lJS7Pvrh0Mrdd4+dtQCZ9cLD07EKOyFhVu79yZHxGpHpBBvFqGpfpUfjO+bbd3HeGdxNBY8wsyEs
9lvoT5vjVqHm94FMRpC21Zc6k7fM71EbPE775U4UiWpHWzXfY5wH0B3OPE5IJVtth3bODy3yRgfM
He3GiIgfanhppTtszuemQWKRuR4pI/3bWbqU1eQ5tV8Jv00lM0pjha2AVvOytTYs8X8DkijvYy5D
KlRUSdjwGgyDsfkVxbzoXx6Qq2IREKLrZ/xPnEecOoyXiCpQpXweThKzoETMaSlix5JGxXDM1sO7
spoIH2MpWLFzSZ3hoL4eTd9ENUyLscNhb5n8Q57wFxBp5gHuqUnSTSMn1BGp4SAwKmWaKXCCdjDN
dvq7WZ5QuTq57KtRs9Cr1VUbGbwucS4V9TJi1tpugb/E13gmG91ZEywnt0aRIgNyv+HapUCsZDYO
nBucsE1osIhuRX5dcYFRnRrmaH8SQJf397e66t9JKOD48gq8Y5ZTmGx6+3B6zfszOdwFM712PSeu
KWXfNm3ig8p++M9Pbt39aAoj070cjp8mo1uAoCUcIclG1TXTTwXin1h6twPHL1zaD+OcnRSk5xuj
8yqdG5satuR6mWlE19Dcr38HdSHMc/znxf7EPw1jh+V0dSKxSKZkEyZ//bfFvR9N0um6Dl6c8Rtv
NA8xPne0W9WwRHC6b5HsTzSHaHbdLQsTCZuyHd9JIu1KLG+tFFwBkiOM1pSbkh5LKar576KF6cg6
hRq+OgGrGu+uu9vJJ6rjDa5fK8jGKts07kyq6psYLsFlGTSHS+nr9hIfdwmk8TrVuCnoc2XB8s4q
hU8vur1+ba+75x4WxSgiyHpclaK6plHwD135JfQt/dDjHw2IA6Ui/pZiWpatADFDB3h9YJuWH/FI
TVMynG4JdcnWKpTY8QW34g2nZtcTid13AAPptznkjmXMJJRXYNY3jKvtkZK/gT2EV9Z3qAoyW/3F
9wGypnQG7DS5z13obbTZtU7QTT3EIJxEMOZEihdbn2rapqnVCLrIqkBTdncPGfHa8y6wf8IAOSkm
PisMIzm6u0bTgOUPhr4yryD0IIypZrLAI9X4xhSEZ27wy+vzd91lMYRJu59XNNnERxhLUKO4xGzo
O6um2LI+rFH82ZQyRSjbF5QIkaWYCiIU3Wv28ZBB1RBK5ous3aCjS7q+Vn1ZtqMXwVhshNQwSUjS
HJUDayUHipjHq46Llm5Or2byA0WjhvIWKvWyAHXJqaXYg9RHBATwvo9kbfH0JUbiBrr5seBcfh39
pmHJVGDZ5YbZK5UxTE0SNVg3FBPVpPvRI1JLFtOZrvaBjoDBo4xSykUTcOIOdKz/LYisWTUCR2Nl
gfRWQC65TrnCvxvRJ1DyxoHUAgG1qmkgFb4qUHO/wzo++wXxJRyJ8ce2Nf2jKE3nPA82g3Wx6ApV
nIvYbuirV3tC/wTYDYpjwtEoga0k7vLpNUKvvKe7le+wmBaglD67hNn+5gNvAsHauhU1Lg8WYBUy
vvOY0Xx1lOkrFEpMyPGIJb8ik6cT0SV0wTtggYUhIlDxELLREDj9nJYaDYjHZ1gDu8FMZGXmhuZf
js437myR7t1Tu1CeSr7BLIx7UxajIp5eJV8AP4NdgKAOhdLT8sgIqhLRvyXfim2Wgaxc62nyyRnm
emOKjI9JTSuN1RceSC0FxvZQVevQEEnMTVXBHhU4D+mKg0NzNtF/JUwuugGShKnD/+QsqesmoF3u
nXCDZKO6T+vSA01CaM3f6DXPxTk/CZQruCtJ6HKjpA52OoXU/nTQkVqlfET9uQYHMRX5Fae4ekWc
rKXOS7EdyH2QmBsg7n0IECvsNxRQQbEp/rkU79lXCHSDOolFn5VEXrFz/ecXWirVC/k5BFSZCOaG
U9D5bLuUCGeeaIRQBgx5UffEa6UtE8A6H19XDui0nMnnNxcbtR07gYLvlMpnh6auCg37R2aLEzFX
ExNiTH9aLTOlPIWs3R0vWDAlbUHIU0NUyzIe94BKXQRFUSlTqjcpeanhWkWWRoprdmKq9tykeDCm
lXpKgV2BpJz2ptiyiSHv2/FvvM4ZRkrTcMW7rojhjZTPZOn+UEAtQJfkjgSizBdNgM+c6nIYmdfD
EFcAFQty2JvB9XaXLNO1cHPqQUZT8YjQXMZtNcU3TNzR/l25yyrXlhHh27/Rn7dzHDF6c3vizGjq
9RsnXnxPy6kqs0iaqJGHkJwYkw8cvJiXU5FjtPapi23YmjfBul8uh5S2sm0CUHtJJ9SDSanM443h
gxdWFAnPdYhxmPSL7UMKKdeZAzVL29kxYlfQYxE1WaemM89ISPeKYIsCH0Xe/9xbuJPm1UQ5fvku
jbC2a/8LxVKzwKjsH1zh+yIb/zSWgeD81+cQOUQU984u0JJVZKocas9xah6N1NYcZVnsWIXzLk9T
TzI+gIlA5wYbHehUdSpKp+YFwZXxIs5GQPzgupAZfuLrgmFTwhZaJeVv3B9kvmvpFWl9/lEa73Zd
AnU4bamOn4CZErS+du5LrFmA6Yo2g/jDyPZ6w/CCsgyfdWA/LUFpowCycybSuTeVln32zzvmo/FE
i4evG9/QAY9h9D+g1PfpDJpKsg04gvYMeYz3uluwDdTqRMXAKU0H8tigMdlazUsG7CNzwnZbwyEF
d2wOOglowSjMQORf4UKN1pQfi9r5vx++wDahfeM+rymONNjMuRr0uyY+vqHJi1EfEfMSrWJzio5+
7/ycEg6wpC02tn/S6hC0PCblzeApNe2zwEr9Cxwuvq/KtOuTQnrnwdab9/qPaaII2YUIIj/rBNPc
lVEZPmWJRDdFkMd4jcCK5ph8+U3itEMc3N1OBFEyw4PkYG7gQ8hk06JIO6nDSd3vuZmYkIWGB0h9
XG+c5/pwjtLNzSaZjFQs0WKcVUpzpewSGlBlyVkdUYhMjxEMWvCuOG9nAGUdlp/4bdLiFxGYI2Up
5VzRQUWOmIzQIy/+Q6IVNUtxMgqKkCsF1yNsanI4reai+5qsevGOG6RL60YVqqVWktSar90GVZV5
jgufizTj202Wc5guXNDuG8Amb8eGZRlLrRWJcvGmE+s8T6U7ePBOVGhEOVj71vlt/U1lUAgOOG+6
ih2YwDUiWBA7TsZRfcV75ST2YGVFTLuPvWomnpwzkIw1WRnE63yoCz1Ptn9QQKAAojcjAj+t6dWP
EM9qRuc+QnE9wRJtUw/JHu67s2TOV9hWGxhV445K7SkZHIAyznawWqu+XzS8unFoqjpGeR8ynY6M
AyFQZZ7F1PZeeVsgIgK7OmRvw2Nl1ywbt+BSKs1hnSG2c8e6c3sBG2c4WOSBtxSYB+rnseAygitR
glauAQVEuiFqKphGLvKGCXzvPWwC0cg0cDXAIR+nxbsouZMMN9/EmInjY1AM+GK7lyNOhfb3tsMB
KhYdZFqVz0l+CWUApcFzzMTLcCU2MDBYNB3v3w8U2ySiRBlM0hyJA9b41r42NUstcLqEeb+HrCMY
LL89o8IjXlPPvBegKauffX70UTk4gVQABfrUinwkZY0p1vrg4pob4ONcTiodIhkQqWEHMVxHCVrA
dccUkRODV+IrTnoQ1FxGcfkrmHIH+AX407l+MOcz/kmedF2nKW0GYpEgayg+AAyD8u0x1lkjZ3Zu
0rp565mAg/SGU9FInPd/lKQ1RKcBWFmgAJQq1Ijy88dvlWZXQrm7xly9jwKAgLWP3tXeWUBxH6cc
IqfAHLuCGHuBoLTDCQOcWVyx2SmSvqrWFaR1OmrtB6N1STgQSCJ5PcjB6BvCgPAbGm0Vwnh7OJLE
Nn0h4EO6m2JhcfNuXIg5pzjNXE3M7hj7pULtyyLrxwK4LS2jRFyidcRUILG5FZAIKevUp69izYT5
vGV7BShBJkEPUz2ezfXk87xz4wHWcHQ0suozbFZKkPHFgs1btvDAedRfbcz0/6rqzEi+DvsS9F7M
vcXgkbn0bVgNJf0k7Jl0yH33gU39rCO5TuaoxyL0G8+3QwxPJHIX3qCQHov1q9i8B+zB+3gQLdOE
CTpsTQo/c5F6Rd0G0xw2m9dvTkD6GeExV8anEgpxFPT5aEp00ZReSIo+YMjEeOgvV49aDHQ1fvvy
Zs0BSynDybF+j0c2dFlpd/PHd0Ij1iyE4RPRdhTt4mquaKP/u26Wi++kae1G/Rgh/nQck7LUKMcS
cwh+8I05C7H49J5ZrnoFe0KFRDEgq0b52f8Cj0Ipg0qHyWBU8peJnM7+f98xgsVvFK++2sHzeKa7
N22d9m3j7G0as7gUWMcbJV0v1Tqq+nIUu1yjAxpdm7Gobi+WTRB2i02i6tjkjmcnX5rB4o2Td8EO
QSqGs4Bxu6fqtvZuU/or9B6cipNpF+k5tA3ArQXhH0ql1/2AyoG8XSUpa4BokRhM5ujbtpHlrbng
lrkonoR8TIsy4193peiA4GkeNJn0z9JFVihajZxb6hkTu4w3Cz1SMbBJflNc1VgqeQGhZnMXW/MH
gpH3HxNWr/2IoyScGa72Jga31GTmLClMNIpbXnbZhEf1u2vJaQWB9HBjhcP31Fd2lKvicf2O+TpM
n+B0vuTlZqP3AFCfIReWXYVETGjOsbW9rNqoSU7sdx2aJoc/8AAoJKqG6hPDax3KuXm1QBuX9/Rv
sVW8vvxljjRZCV6bR624bLqxNILRaEIWPJAxBC8Ki7jx9L/YWcaIDbSZEBJuIc+NvuyzTHX8DGOv
VAdJ40KLCr7d8IATxUNnWgvEll4oFsvvJVoCD7ldWKhOrkYLQJwznoUmoQnSbNfjSJQPM8nleKs9
LdasrpDu5Qf66kWYZgpa8tUCgwBDyhrJfD5YjoeRBxdRSR637kMMzIU1ecet8Su38eKKvrrBilfB
Wp574MnQqnhNE7v3y6Gifsy4kq3hzeXRtYx+MSyCgw4Z90Xv7IoRYPoDxT9KylwM6YBCWfDdTHpZ
+BB49K+8l8jHlYo1jmb3M4qvdb94iyeoeIGEZBheCw51A2SW2jH7bSJCCzRUdXpUuaaUlGgPiRgv
IqudffwB/BqUbfgGyPcY2n6ScPXl8KC+0psb5Gqrw2FsuFJ/bvQjFWyN/ZYlsNGXOUyE7MJsup7D
Fm33kHVGkeQDabdbx1e5/j8uZVr2+dL+X+rqkm0OMxMrDfdHqUfo8LQYLpzCdSekAN/EOyIeIiTf
hEMEdVzarPtae3OKeocvNhNY2QY/FWNX6NSsA7gRnDNa+YoYEb/wSB8Tm5uPJgGMp7AymK67wLfj
6dvKMC96m9jtri8uRe2Xa+AMMIBfsyvI2vP+Iq9gXoU4SPYpuW2jOqOdbLLk+bFVVT/dCFOve33x
Bvy+bGR12zGaIII+c0Q7eUvvbNnZfaZBE8m1I54/xm1ZP2aRQR1Whv0B8yzFfaErEjotbHPytJ/2
5rVpp+WHGVrUPNUUWaLdrIc5TftALppi0m5ljFhd1CT6SGQb7i6P8F0sYlNB6O95sYd7LLbTWR+l
4NohsuW+pJNJq/AUbLg8rbw/QMGzQB3r7mXH3j8F7czGiTw/O0WlGmPL1DJmi/uVsb0Oza64X4U5
LESftbp2C4yK8bi8Ou6+tXS67Zyii2alDf5ZKAAijZtVUUQxE5dHBJSQAf0XxKD1qSY2MYyr+318
r22WGYKhKqUeTQQm8Qv8/Tw0Ia0ZNk0eXUQHWanADMsWODSE6dJruyhPjtSNSV9qiIxK1Iw5F08M
LHpWX2TNexKTN98sWDmr4y+rQT3nIdy2+4oQxiuSKr99SZmePy0s79SJn6TVwahHMfhj4YXEWCgA
Sh2ZXB/og3h0L12xuXDepwfJYQB/YYcX8cZxkpVDCOSe6O4wys/p5tK8hWI5xx+f/mXjO6BcNq3e
RA+bXmeiXMxC+SoczG9gvfSmkvuaw62p018W76TUAggfuvXzFOaoj+mLsKt1xTyIA92kbNXeKtdd
n06SLPCo3ohQZtDhul+DqhecUvmvM7Sp2n/M9iseIIZnrhLVO+a4MRcIeOxC5+NxIcXbef0JJoNg
tEpwY/IHvdQ8fbiyP77IAUwxV4SYhq9Fx4CJVSNRQUIwdlWXdP4WMrkvdSNEleBB78q5/RTva18M
8vtvth9G3KXch98ctiHbCE5j7mdjTyp7I3ktL3ba0BgjQsNxDfTXq9BSWB4M2GgNaZP857Sty/Ix
7P/Rs/25GTl9YtqowNTmZCYqf+ertDgWvNCVgdkNELUFmJMx/T0BGjsoZQQKfuuCJoGrEhE+cdSr
+JJnwapLrPR5SP+R7H6DFMwbAeDNlDNFymdtgKdosYlK8jRCvRqYyTDZGjyset0iIpOxi+BeVzwk
HGR5UxUXMKcRVLtisjbwtq9G94qwKSNdR222LTSeFpazuCD1hXHTi0y5MlFIG28dQE/z4X6nFqhb
1S2tDvcRoe2DW1Aca4hZyN70/1CGdmoB9dQvC/pyfD3cMpSA6KjvAOst6Qf+LFg1RtDF4oDfiR1U
4KDo9oCFqCKe0y8fVAskjSKPPa50vnpjiKfw7Zd5hB3V2+OMtqpkTj5mwx7DNm1F8K5hKrvm59V8
/eaS+JGKKuhEpF562BQGjy40naphayKhuYm/1gR6WTrE/hIvcJcFNq2RO2p5K8EYTXoZxFnM5Gkx
CKT7ZMOpZ7FI8a3/FIMjdT9lxnzbfjAtE+qRHnSL3bJx8//VTQHvMDuZ3EQQJkh8pEqGoQj0exOt
Ecgz66pKIIjnJqKg/HAuw8KZIvcWxgMeIJKb9oiUY1YuHOvbhaVGfyEIljqH9AH+i7SLxPRIzJOu
pxJgHOX7v23eKv8kphtYPb/OrIOKOa+BZEyArkhUIyO6JUWvHPDEgNBNJ1e+4ZcYEBjBRSvW3jqO
BV7lGeo1xcaFNsZvds52HUDCtvDqNaCD2SXXWrwLfDgh9bWW38/qvqNR/ndDS/VT5N9lL6RhM4we
EOPcIMh8z/fzxsXuI07jSsNMmYeZI5AIlhm9W8wODWqb0S4PqJ2m6zv+/RyYJ38NGNcku4QxcYqI
W+MeEGsXNFouz4t6Ln2GLZJnntA+ZAKQTtFHLlUMPZQnsGwcG5LLYv1fuiBoy7Tzd7135LKDlnmI
I9VXJaMEgyA7sf2SnFMMmmf2xFkRYAlnqCrjnsLgvyMISObEsNAmda8QHaZabsWURR4GBXh/5e2m
lq5sbrOfcHr+2RhJDXQTbkR1XBmajhSTsfKGq6gVxfeykYc8iV83U10AvuFyh580amEcIM4cQeIP
58+O00DZryI6BpQ+r2pjpf2kQ6El7kY+RpJbg5TYpoM9fTlb0ZOazSXwK3FAksTw2GKC9MsRkQhw
J/+Yi+NveKGBs3z/rIIzpDyudJLz20PkO/yB03dMBXsaS9OI5N2FW4dDzcsS1wl6aKXFhn7wLE6U
pNI9WlYkg3HAR0X6lS/l9dc4e5IlWHx1voSKlINvBdhSXOXRxCU/sOY8w7jdtTNtQWS3pZRNbbgv
Ov2XCl0x9uerb6YNyftKMPduQVg3n7copx4eR0mqODeGgbadMXNIbNdsLcMZUpn/nOg/ay0WnwBQ
dkuWw9lKG2EB++thqYnE/zLqicHiGBa4h6PYmzy7owfI/AixFT2M17iZ1/P/ShseDlzRl3nWxSHv
R7t+PDpkGBN4y2fPEIlYwcZeGfDZY17AHA5t4YnVUmbnheM298sYi0hRvJZnb4nqrqy4H+uNBhaT
rwu8FfQ0wJpn8ec92CVCA91NubocHg0zP9aK84cMXiCEicsobmUusG71Zbv+kkgUvLT2fpvgLnlJ
KHr5NrXLtdnzk7x6boOk2y9QqMmrm2n9JzGJg9RuP61jY7s33uNUk0BUR1MByA+JbnvAYSL52KsT
JClfT5qanx2qeg/2UpC4r4uXfpoDheBWBeZ6QRrZJ7si7koDO3ZKgPd0PwCSKZum9kgxc/bygRvr
UQTQKOCY/RHcdJK8RTrbpdBBQrneAkolgQHrmtd0GFHgSvU+RmNQ5eiLbSOrVXAsgzsv7s6WX9Qh
qrBxQeRDiLphNM2LfW9ZQtDmqqkzSiVNAeE5FBr/Tt8vlmh6rK690X2RfGIzlBpgRmME04B/QhPr
1nqn37njK1JDc0mD/TnepfZGS1DMrFD7Rv6hoUJAS2AVgDYpkHpRNrNYgK+EHFhF8KSFqURciaeO
qy+IF9G3IuDFNOhYIdIZ9eAG+/JfZwL0Jokfk6IcJ6z2ypzs2TYoU9FQAePm2GnL97tSHQzD/qUe
/G6TwshcfSO+1aYmOmwg1x4uVeveT+Fk+gNBe1KYMc9ch7dp1QhbXU9iEwmFZn4xi9Ayi4u5ogcB
yCVNyXh7Sn3Gt1fHcEE1F9yx0nVtthUVRIwd82vxGzDGS43aKMtygwruKhEWtNFS9APTVB5SFMjM
gDyYP2XY7/pbO+WXmqkNgZiXTkmHWL697mci5l5Ct1Ao3908i24B8Eqld8yIzzVs/9qNzfGHaWwh
KB06ju7yDb0fQ3pRSgHsxd9e46irsh6++9Ayf0XSj46ob/3JkqjC17RhM7D3Z+0v/iEGAdUt6weY
ZLlvzCxsmO4eg0PXQ5w02aJNoTf4x/AEl+R+l9yTTqm3eC78Yp5HBcJlgl1ktcLTjA8ew04tjvnV
oqZm4mmDZNZwZr6kZTr8H85TYfhJ9bOSM17TTk9H4yoW6ZmEGDOhFRmNIldoX22l4MAuhpoxYpLM
g3psOi38K9TRHTEeLjxbQA77HX6zN9yWSAzy54hVJqaVRmqNlcygxzod8tbz+3bUcUf4aIjmhuRj
agNHihrUHMEAw6XoXD6uIe4FIqTuCVNLIBll+ZwNp+XxeYc/1Md8GaK2lExcSeBHC+GcGaUss8cj
hF9R252GflDWR37S4f+KpR1vQ7zK6RnZPAJ7OYt5FGkiRcgXVHSa7wFT8JBPign2iPpqs9Vwicho
lY6OC7h9jayKlfOxcW2YOc+jl6FT+3eFjQDHMZbVIiZekCIlmNYv0p3CDLbSmAN1MfCr8kfHxgzb
R/crOAsYcaFrpYcSDmgxn7zvgN088wbztIi6R8G5R9J8VQDEK6plkY5PoDMoYGZJ6S8v8y2dqOQt
RN2XKoxgGpM0wEZ9gjaIJIHvKkLrCYguidW72KGdc03N5jcYMHabG93VrhAwiMWsYGImBZJFxkez
z17urXikaXZO69gSHERATtJU5M8R/YdKhfo/nrMnfXfqS06ZogVSXxMplp70GxVYNRDVUwWpPHhj
rl72bWCnSNW5jmCtbi5KYSIsvrAgZVFj+NNOElrkTbVMMLF7nwwSpbEs+lXbtnmt3uVqBRYzPUsS
Xdi4aVAHTBN4/6DDzsz448/aARQiSE6YbhlRiuxYwxbaS3e02/afz59CnbdKkfC/uCNmFgWHwPST
vBj4qUpesrXsEmLNpZVxxm5xGmCytIrsOMsWSpJWnnsr7dq8KeYVHPQwc+4YZCnEUnt0poucWAer
/7zsCreu8bfQMgx9vDe2kHt3YZpztgECmiXxVgijcvC+mq114t+MQyOXlaURGBPrGVLupeudT6Et
9srIum/8j0tbRRxbIE4BXG1DFGun4sJt3camgtfMS2yVLZ9Mt0dhQGJgZNfsQfZrLl4Y1ij+OmPM
4gm4ju6u6XLszzL65SA/Gq9ct/LDq6ceDBQKkX/5g/dCncXB8wTP+3Lb+VK5u4NQVpUSMa6a76w3
xvQ6aDX3O3mz6+MJZ1mrA8iT4f9/UybwRwaZwT+YFloeJwU0eK4UVbnTvZTZGfRZgTyuk84C1DaH
K4VlH5+54t/qovrzmS/9mLJEdeml8U7Xqn+bDiF0XINX3k/JaB3jWVoh+fOS5mWMj1n+Hry+UVga
kE+5aOvYKfQouFyCyvbJ/DtsxBKe97+LOuwtMThDB3GjWrKA8IuFyxv/Tm3J8Alln+1eZN6nJooY
mpW5cbSsb08ZFUZR8BJd+ak9zeDSxktC9QAPK2CYJARcteROIqVKLk6eVBPNKmqSx1xau2m0Oyem
z2MlzwJiuJOxs/bMulJKBIE8LyHQpjTtpcy3b8XqWSf/YIZgX9ZejT38Iq6FWGYdYrOeu9+hSqh4
qRQOwJaW1YqAqKd23B9ajliH/y+kOqKC8NWjA8q3p37+lxqe3m/EeP+mOFXwTW2p9p5zskdI9VjL
JgAetZuvq/dwvSSSa78gPNWP/EYxj/UOIS6DeV8q5ZkUJo3kY8oGaoGEfTrPv0vK4Q8MvsrZneU3
vShJfjuZZW0whjYnM1Jvi6yI/EgV6erQgf6xTHPEpGRzoiZoo5aO2BWoWeOnyoWM7kdk+448OhKS
F8Yp10EYgLBItj0Jm8GekUxSP0uVhrnglypeCWCYlBGcrNiSZxo86iE4zUjMYtQdbg1IcjM8OEDJ
Yhmid5Uhj4YH8YgnWF30DP07yslkN604D4BXq2g1QuBcCBuj2TY6/5ijVZBloPk1iSAJDRfeoSFn
FuBWW+1+f0u4P+ZNwKe9mDbQAEq0gFD7NVr3bYvP8UfhGonFlUXINCV2rF3meJdnpxdLwRVLPcl7
srsGkn15hMfGE5hJIne3Z58/TjtcXzTtNCk/4N9sfQE+wlyQmqFygXB3Xw16MPbEU5wCIhaV/YmN
ZFmzh+0H3FCUXweHvlsaAev1fIl9MH6MSqHHyyXGL6/FFSrqG13laazlaizLhDKLkdhRziVXGGaK
sVZVVGOxHi+pXwq/r65rEw5XK7r44ase0/Zx6e0IYFoG0j+TlNNbjJcuGTLZh45l0ng/5AhRv8Zu
ZVi4lknHtEmw231Q/RUJr7PkRM9ysb8h3ePIZ3mWE0rncqeRZz+JvyuusXdLVkSmrbK/sv4x/3+6
D6Zut3sVwDVYgs77Vci6CD75Olduh4iEu26NtnirnZLl+RwXUxWYHXXHs4nPjo8iZV8daelSWkRP
qF48b2U4ctL1yltjjgJViurhD3KdvpfBisw7igGDYNb6YlbNdL7XphxQcy5mYUwWQ+IToKo8loOe
k3ExASUgcBhVEy+QAFb1jwwIhZZ1NtUTDzOpRS60y1tcUX1zW5a5WwMmXhEcImlRehSO45sZfCNg
7YfzlcpF7zGVn/yihuf5STiJaRq+M73q2tmxoXeFn7hBvU4l2X4G+M9r0E520tRnhlVapriTXQJz
6igDVVXtTNsXjQQvcXRo5owzLR6s8NeZRUJ3IMiEXGIuozyBPkE8Rp/XgIS3WdOq1Ea3oDBzj/oo
p+23gbNztuUgxuZzMCKgfUOUi0tDE5RYGOoii3Sh3dDW9hL75o20h1w5NR+nwapB1F2/oO8u4x/X
KaWR0XODaz4+48gurP0W59rf10oJdbK+gv2h3mCsTIhr07Kse8gesKzIkflCzNRIxIFmNvCrQB3m
uyJb8H9A+vCqamCMdlM8u5qTRSSRIdtgAH1k0ovOp64kb8peHjTmzdTk9I3f0OLKB6UMoXIMzvUl
tMzCJCjbfFQCy8nHSKStHwib80LtwF1BDQsKov7E+lAd4yOe3JSd5uSEhGklD2tHdd6BvAVauYM2
t2ZWQfrIzdBeLAP0gk+S22Ce4YmWDlVHDYMcxSB+AJ/p+0QytMDUPAvq+MkUcfMqil0csAjY6XXs
a+mPStvhedqFQjU3qgtMIhoxry4W8vfPbATjo74ffaUHP7FsvBk7VoMIcyNL8RB4BXP9Mzx1XGsY
/UdCOoXCqwhD3aVwAvDc2fvGmNWJ/g60eYAmBTRMYT/+UqcoZdQ29LeJCRUwN5vXym7DTolMIxH/
GaxvOd1iXFzJ3tA6NWiUdGtd5a6gFZfPzp63CVmpr0pEouPynntAX/v4280DToTZOhauzkQPbEI1
ftUv87yVpzuC0KnJ8DVMLehEw5WDHH+g7Ve2Z4YAyHqAQAYVnQRWtKF5Anf0jZwugtbQuAln/k7h
vz7nj5+nkyTuBXWbfolCTFJEySXieKooPZRSBjxYdpoVMzmhnEi//pqAYC/iiN+GsJfqHOmhD36z
iULRQeNSiarJqei6Ru9wChDyk2Tj5ow/ZtdEhxle2ENicNrWpO1GR02Y/lyUBSF0JKP9rFNYoGyl
6nAfSup9WN2+KV0gIfF6mECXE9Y1kl0CnZ80Kfte5t5uJ1hI9gKgemFNbLf/+Y59+BmPS8RGSWzk
wkTiRHEmcit2hGFiLzuG/mhiD0Xgv05zkLCnSuc/PvPqAoBkLzRseADu1MDlzJQKjR29b1INaRlS
aS7JmI3ZXonQeWwt2Norfhv7GZtNzMPJEZjGWvDdcVqP+kwhZEOdkY0JHkv/KMwNoX293d4/3AXN
OrIILimB5E568gryPvlYT1/E+xUKOCPtWRkvnDrScl0IFM6ENxs99VyIt7Z1qKbwTY2U411X8CJv
LZSGtuJZ9pplJ757i2bwERLHjmU9J8Tc4SSjKNPM8QwwvICMz/+RE2MVeTZ1Nr2tWyFB2RAjNeMr
crmTqNgduwYnJV7qNwtwqBtXGNbNUVxxJBLFnh0KuaWJmZ9gmAO6XUYx3c5zitA2dPZyhbIGqjpp
H0hCvNIaE0q1lO3K18C+hzpQvGLd5LCl4GCqgY2AIIVtusZzSUNUQbFDlRvI7H+TEGjGxzglihvx
HwwN/wXv4iPY1Gjn4KZIIrfOO5khcRsOAxQNbce8yZ7oQrG72+ZH7nGBlk8XMJwngdbg/Es+kqEj
3QB8Ip4XvoaeX+f0kBXg2CJ4S7TCicX18dr1DIu64wYyeWNfzrEEU2QpV/+0RKtRxJbGyyg9lgmc
P1dtbgQ2fiGRtmHaLRYC7+w750Dr57sdRAKBeqdrca0PPoFUful/STrJfjhwzZrweK5VrRmiP6Hf
AZ26VDt1SKHk3dD30yXlXb7QQA4q2kgKRHJMNwbW3F6Dbr/oz/R0y/d5ecqL3KjAzvQ3XHtlSp89
Vz7j64itfcPjo1zKq4sDP3Bxdm2lVbPm5HEsVrL43wlVA+P1BOUW/zDM+J2yvCTj9TVYJ/n5ANYd
zahNgNgAJBICsb0rOIZs1fiesTfnTN/5avY2zQVMutBNbfpjDwcF7jB/Wc42YXA7j2Ysr7nlI5ia
1HixVvS+I8tuzuKtRGRyRFSzfWNvNeXBLXsa3K7nmN/HeauzWudI8f8CAag0Nowo1jnHDcwNgtmI
/XOxrjseU4TimYr1UF4mL8jZOTqTFVHeatFM92Uhn43TcAK7Sg6/dwWGUHLQOfRI3HbCyChxOCtB
o1QoZfvkcNtDcAKR5i3XY9BLfMiv/MXG4HBJuMdMIRrm+txlZsVYo9e7BqEoTpOFxCkp4E0ku8ps
LlOqIhw1Cgeq3HDONXQG0/8tgIzOibnY+1nktTipA4de9Dyo0zlldYsrtq1k+aWWFGz3cw7sWl0A
zRTFk07DNaVM0NhVM3PqA/Vrwo85scd/Sp1dNIHh6fEMIrNLvT1jercwlvHi8dcW0IK3tgZRkHyb
BGGFi/mwz8+7G+vSv6o1ntEthlrzYV3EW9KiY6iwAa8Wz/U038rKkfTigBgZXsaNjtTYuBmgDBFW
zXUzBT+W+rKhTiDHKpWC6sMMr0EcUw3UYwH4Q/dsDKsbkzpdIYUYlfA0giqm0KuUVBNMzYN70Cta
Dtlvzhp8rRIQiiwXVvpSZnmGIHZM5A0IXiCf0F8eeDeJKk+BLthSUeJXmZrLEwRCV9ATFyHUTY8p
Gf2cttRdO9uDQKiG7zZ6fX+m/Q9R65pIRD2EYM9tU55ZdDURil57SEdKCNzW1TDVvhZhp4eByc/z
a8/9+fa9plJJ591m/orR++xD+BZGzgY9bj/NxK2fbOaVDz5FdSuFIreLfAITsPd/57YUOK5auUWM
VJcFlRakn7IchpbnHmd8xXn7CRLBq+1wYEe6RzEO/p5/4gpI1PyH2I6VwTpAVzIGiK65mcSFFw98
NDw9dv0pPaNzv1H92C5e7MOyYCHiTXp4zHf7rKWVnqCj9+TjuTV3Y4Qcu8Tg/BabLctazYbxiPV5
0ImLETFIpak7NKSri7LbDlSwGbRjwDvUQOvd8zIQr//yiYAypiMVv44/E0yuYgpxFtBy+DPy9xO/
uTDnejNaNVFRzLE9tX1ji4xD7Bvx+6fYOXR0wyzXgHx7Qw2/+JCryLJneFeqSpVdja0z1VaFhOYP
OjmkvXRgBD59H+Y7DFwaLPUr81xffgC9A0cDCoDqYmIkbQ7kDPXUgQE4xkY4IP9KnxJUEXMa0Dna
Ql+owWOsTAMGnqlNUGUyBNltmrwDYU7uaDO6tbKWgdEn3PNyQjI38U8vr7Lo2b9FGPMbwdUeLUpB
wHxKk3i1S6RE9zzUTRmGoyenlr8/7XgVZxU0O700HPa1ZIoYtsAzoeJdQEuviHitPUv8gMzGwDUs
HuaHLYeJ87dvIX/V0rAh23lI92RVCC67giwfxEaPX9z6TcPrKUT4gPEs86HgW8okRbz26i9afQni
UdOD5QLYFeJZ+8BLcNxKvXMtuTHic0UFv8NFEJAhjN+TqqxrsNZbbeF+s4MzokN7HnhncpmlMwIZ
AfoUK02XR88VfT8EDK+6fTz7joALwt8ooA91mpZrkzrLKLzB8dAwF6KedJK4yOvSlAv20JCaivN6
C/RZA5RiKtV0qmI/3Gau/OQRbNZffzw5qEakSMvPZoqQu2Mzh4/PUOJuFJgvl0wW3jl+b8vbQqOj
4MmOw4UMbQB8PYElprSwgcHBJK81n+wzsiXS/nhDOLxqrtYYxR8FA+dkvXMBpbdQy0gil4qabX2T
ERcUO2xQqdkYFe2lhDQsCQAaUcVPaExNf9IbqNg/bEObvYraBeF2BgbvagKM4Onptw9yUo2BUrVr
MLyESM2YQ6UU9+e7ml4jG47tXO6lBtjurOVkHzpnAXEZevMnAyROlMjo2nxGW3e0DbsXsAk92e3J
fVpBE0jnh4ND/Crmpw62tiOKhLvZ421FSWt0/O0MTsEN9G8OAAZbdeuTEcytnKiMzyt8275Q0KrN
O5E9QHuNnQfbroqTYrYI9C8UYydeW2MekhYBR2/JlOAJ0w90+nzl5Hk2b8+eZ8M4xbI19EaGpBmV
OdCGObt/77DJxEwI1i1rFwhAIFGfXLffZMKfT7vXiJmrwRW7QfUeicZ1QXAFOX5co285Zy2Ka50J
yoH/wofmdchxtbBB+s95TmWavuS3q/CBxxqgBPpvyR9H0qsam7kripeA1PcQvy3TvxRFBojHUpad
G7JSgkPv7I9n+Iz3KXCUuDqonntfyyP5V96VxNH+48MeUw59RKKVMLwXoXk4598bXpZ/1pVqf1jE
1NyOoSInGtPCWTr9h5NN/sSj4wyKGX1ohjgOAU7QFwuYNQUauN7UvAcTsjssl9d+cZF8taJgkEdA
QKN+IxamY3PcPt6l5PtWAQZqyewc+BSTjM79VELY5bBuWT/d7+kp0nH1hgUHoupUCZ+m2Z0xwY0n
xNsZVHvyrxnU3knqyxKpZs/F9yW+IzWOZTvK+tbHpP9ZyHXiyxv+5vOrqDzv84KXGnPe/MuEMplL
9A8lXK5IPXSafWmWXoN2GsU6f2rQf2aRILQh90WmlEW7xkxOvFnZgt6vTdCIK5nopzX/CquYRd10
NnfHjMXIgcpwmB+wSSSBALZkZOXlzyKM/sQorGZe3wrL7uDh8s+O1LgTMeZBS5FP9svSOrQhO11u
paY6h34JfFmRvY9RnSoUTRuSzDi1rQ5sqTXy5HnUJDQoneNYfmSXm5MYd0beAfVgoZk2jeJnSGJo
T7XrqV7nv7V9snNRbuEcyH/fGgojnUmlB3r2Daa3zJIhzoQeH3LFVY8YrO8Zgm7Ygma67/BlXffK
4f0/nCMh8VW0LO7MOf49Ns3bcJ5exNXJJKZsDPIPJhcttxcn3ZYUeosll6zP+8XTPni0mzrTl3cW
ImxMY6PTiN19t1pRFGEAeUD2nda/GSFNXRxnztQD/94rR1q7pIW5W55qFOQyysRDUJlRL0UNTGA3
7Dif1ySYQJ85CSZV+CJD5UH/NR0V/4iUSA2f09uGkGfSvik3MMFlR4G5DEULyNfph85Sex8NdldA
8ZD6DZ+Ly4aM8nBdZjl1oJ4lQuGW/Yp7iDUsmebd0TKW4v+mblD5BTh0627hxFfJOjFvYQnZ/tV4
9kJin9KjZhE0B3WcyrfY5rhbrQ2bz3raicR1nLKh/b0/jsK0Q9fK0ABxGjYsgQUbXqhPfdnLLGGT
s3gRX6E6skfRLUpy3lNJyC6H5wy4sjRxMy+3WkhPOE0sqw3cG1jbQHwV/dEZpLWyH3MR3Q9ey5K3
j8ZbJUnrq+x8geiK3XV4NTlIn9BHdZY8z0jcojL9tvMlaXrmOL/7cdF26qwzTVpb+NxQVliabaJT
md1dwvWztOtlZQ4Neo/CTVBbTF9igx0f2P9lEu9XSuN8gZAflBCIFVa5KcIQ24y6QYB1BMPwzdnI
J2eWmDg+c8jAsaJfFj0lJWapQ2KnoEUD8Y/a/X2jHXN27MmORmmgJoVAkvNSh02R5yFUzv6gmJo6
2wlREEh5TQB3y+it/CKZq4A/Pv6AkQNKb4lbHCbau9pYCGMAJExX+pGEIQsQQe6+Am5iD1PJOZC3
glsrjwSGMEueT0dAFl3UnvXWJjDKy+M2muJhCw8+1mQ9PRYHpBbSxz2c0n5mpnmmQXFy8r7Ex/sN
z2mi16FYlMhhQyk6M6XB/uINnKqj6uXyHQmdCxESriO0CFZFWmMtWYq9rtHP7qtho+N381bTQU/N
vT0eghx8t+nF5JJootEKDgE724j2BI431O7mZqth5xUdBmf75z9qF4H+k6PFuNZ8bCtCQ0ECletO
fI0Qrb34Jt8uwfKsCYpDeCvcvadNMC31Re728L32/USnJtDwBwk5s46adzOr2mCLADbz7xoIRDbY
Wp/MIYlITm6JgumBKoaXH086S1JEyiv4FGPuQEDpZgcu4RbxXvLEAOWhmORsUPlunlNhC1ItBCxh
zPZksZhFzwrVxOwm/MWI3cfqEKy/UduanTDjU77nrLYYaGsUak4dGI/bKsaHN6cLR3QwIZiKOr9l
U9g3R3jSPCJLJOrPKjfRsEh3zQcs+arIkmG/7crQ2wm7+wNHFJRHsVrtVO8342mR+DMD65z6rIxi
8A7EJSGA7W7YKmbh3GKbNli0HF5ZakqR9YgEN7Ceq/a4tFkaXmhO8abj2FpDd00b7qqg5A2Z3dN9
H6EFlhWj/NnxdpIC8UqoI3Dla8Sng4r3TA7rRW7GPFx8nYRAglq2BvxBNN4sMOBZYa5FTPcNpGXu
9iNl+5caR/7Osm/jwlMUyBbRnBlRX8SsDPoUrLxH5J2IuI/a1SzaUDl/Ax6OMHJu2Js6xBwIvVJj
9Gt6FzchnpF7VzMd5Hk+gxYOi4tlM2o1cvfVTkIbd3S+0whX3VODd08+MIhXSekLDt8p/iz6hK29
Q3Qub2nW0HWl2WofKR1jeVg+i7sDKpYZGC4dJ2patEGbCBH3/zjqIORQzP3HuLnfa7IWPW5y3jHz
rZGSJumBI94wR9vJaA/rdSM0oz/vSYweP1XByqzVa2S7OqI04K1X7GsbqG1EU1FpRq/1xacONZHN
LeUALLx17QDazN2UiWOnda59VCdeyiJftyrfWE1Q0OISE71oDKUEd5BZeEVrC8QIf58Ybxw6Z7EN
k1SKGdxteuzqd0vWni9zTVB5i3Bmp3wuE4aq/UBI9ujnGavv9rsGTDgs5BwjvuFDyZRt3DW7mEeu
QA9Ig78GNl+voo3Se/fVkHH8juR/tbHKIfbJkcziWAAZFWJJq8GFB4tbbea3DnDu59/wQBc6l8Ex
kJz35JLDkNl1cfmfFvK6IHm4XYOh57I+rm5KZP5WUyOMOd1vGNk9OeuqSRXomgiwjYSnO3lqiv/G
1Iy9XGxMHdlvReXpes2Y9GFzKXOlrkxgUB0hJHlFUK32OGZ99goyzlpU6oT1QxHXP3bcnEqDUc+Q
Aqzyj0m98+l24eWvEh9VZNEgdBjNpGmTwvPvDW+DxOUYPaQcMcmOXDJW008yHAqU4RKf0NIfe4Ph
2gzY/BawuFlWVxxDFQyyOlXvQSHCIUGQItGhHaM1kZknYomp32E32v9HdsKaZLAYTKz4cSuwDcXL
m1EeNxUMJEwwD4H/KCwDLC1U/FAsJeIaCr3l5yLvhF9TY4IVMDNtSLoOEI1S0on2Oa3dlu7kmW0n
fIhY/7KUjNl/oBxQt2TFw7pefKSjycktg+HTJKa8d0XlYnDNcEcUdiEO7H3oDkB8MwC1U1WNNs4o
f7kcQDT6vTVa2p9wBpUaBdFUTZ3/3N14tnIJq3vrRVTTW0Z0d33xPxG4Yk2aC8EteKCNTefG+UJz
nf0qXHPVNkMPcMrplMWU0yR1FOMly0WRlAZJJx6/9pLZNFLO/q9mEZYyYuNR4Nyz4fiUAj2d0ETb
Z9cod4DNIDlEN2HOeePBE573vdn9h5GCoq46s9pXiFsuYvW1um0wylvBar9vuFbDRrl7eGXzyQfr
nvAz8M3uQqSsVxDBJOqAUeCdm+k14icSJDDK8lNSvN2FEVsE/8JkeKsGmxakHDrYclh2oypDdKIJ
mCBM7eu5hKKAK9NXNG2LcCNvPmOQ1aDO7redJC9fRhlGiLLNqBaduzfkba9RH5qM10XFQXEqSVpJ
7yT18LR1feZLf2JlsbOb7uGvT70m4Oo3WFmHuwWoEX5Dv3m7LF31rn1AIig2U0uesPe/+ngLYURV
X8eQuU7UWxRyJ3QEsIaN5dh+Rq0UbF/Na93H05OzDMdm2oHSliTaDW2krdyPN/AvQ4t3lJ14Zl51
dqXqiuxb3i5AwR9FQEfrNKgnQSEPd1Ac0L3Wpww/Y1RG4h8+KuVSURWnQsgZ8TlJ7YhUp90U/7L+
tL1XQUZfEnz62rJFupqrAASZv/UcHcdoVIELLb3Ipil17+okd+FFd6SW97dULlFh9ycjoGj9ED3X
aS/ktP/93KL6M2VGanBDO7QZeQvuo2b5PXmz+qy+XDXXyEjjaZCHI3NdRNnAZG2teaeC0rAIM8Fm
RkLgRxlbRaOJwMWOGSMG1Fz8TQQpyQflreC24hRM1BWgcj3ZK0ScJLxEZ/+1auFeqtBd7KevDHq4
/tppnvxzvjFKUWk3VqyUzdUPOdmGE/iRM26ydS8DQumMBfrhCuI9A7ZyIe3g0AsoVztgZSYM1EVQ
o2AAoGIfns6LtvEhOBBLH0csyRiBKkwas574iRFnl0o0zRnW4RjmKuS6o27JlUA7bNSSUInoxTXG
57HpMaazuIDoGL1PX3nDp4M8OdV/kQhdCeoqfM9N6lBshkDN76dPG9fgXC0Sijuw2jBMNm1I5Fi9
6krsJ8D5UbtZsd7Mwjmdk2y+9zsshRfLjd4aOhgjiXFy0K1bP+3DQmcBD818IG7hCg447daBKK7R
yfk3G/SGrTp0DQ7Nfy285NE48jbXEPIxhUEowxAx+yXlsaEHLb+FIth+t4xWs7UQp27LJTaT8fmn
T4gzOqwtf84zm7vjy8/1ottCGKrcO4Y3lNZ9uJAYFqvL+RzddRZjoYYM0KhFf7Xi0Ne2yo3IA+hm
nmP+Y02gyxqikgd3gnXVFdPWJsq5+LngXqrrVTcSP1lFnT/LzSR6INEvPYUs4cHOKM5lhbzbDUO0
YLnWrWWEbm7PXjb+s8ShshROdXFf4TJsJ+/bZjyfJWi0fNQCeyyP5pP9z25ZF3h5LhHEex+lXXwU
evU4F5Md9psfpY/yv/yNd93rcmx6bP/kOqnX8OrgDClKlmFhwMJwvYlzxoMGMDw9XZ/iCA2yMolB
FuYFZOrdzR3hRZTSUtxkgX1zEYo9bCVe5DPvLrfsJun7TnTojXrddXMTQYrfI094KZcm5zOcJD9w
AzeN/Iy/zL0f22+oYwpMF9aouVbHdICnGhN4O9cMqWVMYwMe8g7ur0a8BXd9CWV/TRc8Z2dJI2Dy
5ERjhTyuWwYsA/RFze0c4saUAM2WMl0wN0YSBMNOOXZN9EP1MrybHoYbre/MMEyCHLR+x8caH3Cr
j1ZUwWPnDMjNFTaA/spNZ0tzGUuuhWv5u4v1Z6+4CmCkjTuee2o7P3tS7J90dSXOLJtIxx7nrefO
IOg6uG1dnhzIZ3AQKXYzZOW6iZu9EqHI/P4QUIUlICAMME9Rr1XgOv37mtPJkGbepYlO1SzsuaQb
ail4qho2nwGQsc//QgVN044RwGMqIQdlzCqOOrpnT2ilraZZTePIhIpwe4L7M7p4OHzrJDeqH0QA
C95kiwz0Ht8/PgijcHEn7KgVVD1glpETtC89gkDHACKg5bdfBytwMiZUMJYtxoabO6PMLI1B8mfV
3/WC7NZZQ5HK1HQcjVHzzZVNJ/1Gf/aHfB/3CBLzeQgcrjjGKYY+XzkkqgjCkBks0rhc4jdpF8vx
AjwY9vjAogdY2xitgfvGza1fcMjwxb6i05V0soSq3mfD1Ue2daOJ1mDX2vBLLwB5dYKidtVpVZ5C
GMRa7OeEunz+KSZuG0WfMp3BTvyhrdq587iX5CCAu7sxVErgGGtiNVCkPlkcCpViA11IzTWKCDXg
YOVnWUQj6C/HGo8TwMu+CZ72jwIoPx4TnChS69JVvZ5XfrjN6ESOaUldCwiNnYIIqGGRPnK/u1+t
Mak0JdmvUUmUknZul1poYMX21VODjCs7SqB8jlhqvywaJls3v+0Cg0UcxLGN99hX1F8KITvDs1bx
ARJ4F3o+swCqHdEjMLw8QFYlTAlr5ovxhSLfMucY6fmxV8iP4aPHsn4/yknspl3Db5BgekRHdH9R
R5BeZDEMv+F+5jh5bSLasimaDOaOZzGnR8KTDfG5PZooskunorFwau62hbdFIoXt1wcwUngpNN+1
AmSgh8A0jobU3MfDpxl6K7MqlxnRs4H0X4Z25Nt6W9dKqTT6bAqKzDoKrMrpTnWeJ2ePk7ovttOC
NcytaL1yBxVyiHPHbD7atQ3IKUmEolkc/PRSpPPxwdgYSEuYwCC+7QaunJE73t94IcVSCrgWtfXW
lkhGH/CTX97XXzQftjovrlUnNGtxdUeAcKaPL+tqu7nuoX12XsNjKHbaU3OJXsqxUlAS4VKZC73J
lRNlxkU7y00UL03DK73UCixOftjaP38LK3whF9v4ctJ5YSx4WZ9nGMWhZaAOTCgJ65yVxoqGnqg/
i7quhWr2RKW+Fx5ZG6PE6HHNCDCdN8WKMtSkX4Euq4XxggyB/YMH5/e0rLVVbnzsP9LxjiRbQSf4
eeDVJp5lUGBf2UI7Rgxzv7s8c1zQ52tvbWsh9e9Y+Rvt7IC52ArWVvI6G/YZzxZWGR7KMU4PnmI9
NH5viZtm7HkTdmT3M1H62CqyI/6m/4PTqCl7UU3QhxYL+Ln3GqzhsQc8CmXG8RAR+/w9sq8jz00+
O1x0doRx7SC/v3T4qxbaVCaDwQcJvcH9z7Wi+XwEZbYwA04C5TNBzt3DbAihNw9JUSMzNtk23b4c
D5sQq5rC2SnRNxEtjoHEJ5zxODSsumy4EnMAOylx+eUU35B21XJ0BkfDQlXVnh3hrxyoVjdGBSKL
kH3T223VHXZFYCE8mTvBzuf3HRbV1qH4a/Ez97a02ZFo8zINMlhgfRnTeLvAjifcFkWOBSWoZdnR
A6RCgVbBN/Ea8ZZr2Ooww/DBDrb6B93HVA/nG1eSpVsgeChYU1VZPYdpnUzAa7dRmDfS9h3IPDke
G6M4de7h80UU/QIUzex4tmDiLHZECd6T/zuLAqRk2xipwoQqc6zlpB8lNjPM/rAXZ3H2oF8ur8ys
35pvHTNn23JVJVKvPe/+MvWxZskqtNqxfd/FJzw3and8FFaCyKFI5WzsvX/OESm79XFh5+vvNgVL
yCGItjljwT+blbnBADhdH/mqyRUUCfq+6Zw487k5Rb6clhWAb7XFV9MZ2ghPhNY6TdKIMejuYpS2
HTcIogoThb1WtOJfq7UlymnxbZc1tikwNgsfwQljLc+gRix6Hs469rO/ykYrvvTu0h3ZKirS2Rm7
J1+CNrHjBHSAGd4+I8YeXTiLgOYNwF9ahwb26JqR5oDNDfM99SDMUfmiwl6JmOANgXVMWMyaeQIo
mMFUFk1VJ1TyXhzSyAkIF5T4uq12WPR6XtRhFfcgZaS5/mLdCQXH9H73UQ43I+jl6Sl9chikKDN3
gWvzsGpdQOrjU0jI6lqLNbSZ564xWE5bOyl6rpGImqclOrDiKga09oZofi9ptLkeZ5DXX9w75ZxJ
PccuxHQS75Q61ceFjqDFRpomL9iQfakD0+98Y4msmsv6OcFtJK2J/sjpI4GmnvQsCcws2vadHy0b
PZiGJPvxaTa198GmKQDobnwFVJY9tJpkonJuGUysL2SIY/0KKxHBZEG0GV4UjX6VOuHVWOGPVmaW
NhPOfRuxqLOgN/F5h0aTQKReiO745NTRKmobWRVI32h+pF7ObFBygDi8lOj6GYyIf/k/CYE2ZrgM
3Yw6OpZl+KG1s5a0BjnqqbQq8O/WBXy8NextZ99MOGLCH92mPpLlIXLzTrQ95ApPqEMBu7VKuOcs
NBj9ZwiDFSOHVKmZoRoGe0lV9S+fDpfLj/BLR9zyDfpLILlzZy/RzTu9MLV9dAOOJ60ueaqnvH6f
1CbquK6/4wWZZSoDvZ7HKMdadBbcNOrAdlzxzhnbrKhTf3UrACOcNK9pxq7m8uCfhY8/VEEVbWbl
SfmdWL2k25lnLfl00xQNxp+HCbpWhYZiRqkJLomuV1FQQt+UCSLDbV2N/7CsRkc437GuGg1nMGiX
M6yBXEUG7XnreEZerLvQGbs1Sd5D/Y08Dy15J86KrzDKor5u6PxKJBm/nXX5SyaPUiCJK69dJm41
1ClgGubNiNwsvopuMg8RTjuzJ5xpGWINzgI98U9OV3PsITozxSfwC4TfDI3L5aiSwtek7nrTtj5i
zJV8HBkANrN4Iuosb9rLPUj2X8eWobRWKrfZCy6IxFmIX7otJinMZd7cxQw8tHgQUl3l7vcIs4NZ
TjCaJxKy8c4ZX12zAXdgEHTmxWM/VPbfS8p2BzwAwtCFc5WzEgZYyjqzf3DIDSDzfKq9/3mUR9PE
B5hpdUgDWJ9D8GtSFf8LmxO8WbrpmTr8PJgY53/Jao5/syoUE+RQtxmpY0KbdAcIilVlBcH5OytO
7X5h8SMe0QhiLm/p8wWSsRklhoTgfGVk8HX3y3Kkuuye4gxdTB8ECE8kfIh4MS2PCuDm6vryMCRI
UJdhlu+u5aDti2w6zctm951rmmjpLFnhrZMzgwo271cdF6Ny49L2byshiuG1hKXzwJIpliM/GePw
BbKeI/zb4kBnVDDwHuzclIUVVQwNtT0GTlWc/dHMyE9Ka8JZOqmLIczd/6iA6Tv7GUp+Mvayjja6
8MgUmqfLyqog1g42FeDz6zPIYVNmnuWP8jfV6zF+4ySke2lidbNjpyvBqROkwrtAcQZtne7Atlkw
uGWPEPlX8eiqEPYU975uDrCLZ38oJS6d7S1ah+NA3+FJf/TQm//+Cbtzc4HbzUYT5ytQzXkvEvps
GUvI82QB8H1N0cTwb0RNiM2CDvzmIeBIp5/khtraDr7MsBzNz2oKI6iHTtXeGtvpWs6L/EUk91VU
i1mQwSRzYeVKa75YYPpPF0br867mNSvAHKGEX8hT/GBv5089ycn19YudIdji2MaOWlGSPHmbB4fK
3OCtUw9WVq1zeQcPnsNiNTuuEAYXZsxxl1HITSSCxTT98hfiOrGN1hsOq/j8nGHhV7fJTI74zNYr
dTN3k/0iWKVqeorP4w8AbqLsquJKNizILPp/gpgqInbSKCDsLpdlcwymx6RlhYCsLuad/ALw6W9J
idcV9YtjfAUEzIJKyan09EbRS89m5yVM7chWC80u+ZfiGoaAq3WqCVA+IM0k+4IHW9TjyKMXhoPe
GR5ZlQnh6sCeW6naEfGhBY028W0Z6FRbUBS8WSLbKS24PQOO57Npfv3RlA1cU4fYNHNrvb90Y6VL
iEIqCLfd914rQKfz+hFhuO7CDEOSfBsoUWwL/CDNLIuIe72i8jwdHXXdr6Xwj0bC0miQSGoc+HZg
UftmUrMupRgmVck7Z5+lMLpvxYvV6uytcemxJmgncLWBgCvQpwx4mgGDryvjKVGyrvRpQCKHB+x5
sNQtrn5uSGBDeH9sO1PM8eba+TCHUV7LCvgK+ycJMtxdZfdphE1FfUg3sPIdZaU6/CAtWEsgaBIv
hLPnAeQj6pJ17O69fpb6dTuxN4fH3St+LQpgwtSTOoQXAHCXC3c2S9AxexDGtSn8TH2YG956BHX7
nk8tGkfHJwEeITPIBnqtlRCjW1r0WTh+En8V2GjuCb5lnnh2gOszIH176Jq+6znzjef97TWMo8jP
Kc3+q7B3TROXLw0zS/Ihb4PLkWzMRo9a4MZBG36Pe+i+iWOEAWLjxja4c1NIzgAJgd4Epr/g1Lx5
wdIVlZMDZlItZUt4Agr9RTj1dDjD1pvsqAyWHzTZJxaanwkUoaYCZPu3x60ZNqMbtqFRTOmGYAo6
uDmwcwiQYhrR2jmvP2T2Jf/g0mTyTMZWvuHul3oxiKCoJJUHzJ58R4s1Vc8xLBVaThxKj9Ijw9C3
zpG2KJbmxWLwNKfLPH9aJK6yAO6+SK3CIFS/jI0Nd+7A5ImqNoEg7rssN5DDOE4rUMRghzFwcwkP
gtETXONtYBDbQfjia9TxwLNLn5/w5JE78TcmsehssWE5DvVuvf8RhxutbSL3TSUPXGodEfHzEvmi
3HYMVGQr0izw+Ba3d/57bCSh9HBjZMLeQO2ZZCGQcdrZ79cPNp27JD3ehhXy0DRLU+aPYqA5gNLq
RQ8uKxCiPqASnlpXOHZ36fDKP/7O9028u1/qTjfi3gN55myhwieQFoadmHggKg7dcrVFI+1Od0uS
FM/i7EZnA/PypsC1MQkRhwcG0tWJI3epRsW1tA5ByoP+5DVew/fvNkViZqrceJYtQQ1ht2OAH7q/
DN1mfAWanimOwgEOBtRBzJE+3UZBrlVP0/OIqwXHfg9kzPcDkMbDQvaFPv+Hgu0UcE7AebmDcXu1
MCycGRA6cKtZqMiiqp/MnzGQgO+xWnA6Lj5Dk08P26BR3eB0mtVZ52uxu1l0D3rgybpYGnCS8o6A
8coFDK88b0RS3QsfQ/07RsLvTCj1RQ4Dl6Cfyz4/rBvDeWYCSo9KSHx0go19o26J4ZE7qrhx8lhl
2riNpAEkQuYd11nsGY4fth3M3bsqE4UVEWmdac1dmXok6asIrZr1x0Ir/DnZ4rcpnq3KITH1Xw9T
OGm5Tab6TORQjInDCUrYxqJuqZ8pFCjZ0O3wgnhqWHum2XVUisZU83DIFmYU0UR/x+jet0bf7Rf1
Ixfzuk6hUEHauBQB2oZ5cMspq0ugjphPNepM9TDFHpDOcUeKxXwt6ibsWK+EU8lSS6k+SiqPALZF
JEcjW+6GzHag/DNefy7OJHWHOFAcveXmy4I5AA/dyz/VANh+bgXKteoWROYbhzOw658xbGYHzzA1
RjYblxXSzs+lExSGuROax9rTES8S4KYM/0DCNINkKScflPc/eJztbSYjZen7q5wuiHHfwncrk0fR
N4shhMoB/wMeN2vwFiNwaFGSCaUt8wtRM0br1M74huSiLCD01n02QI5CNz1ToDZ1wS8lE4zvx7tQ
3ezwK43f1kqRaWbO1cy+cAfj2EELbUuC77WFJ2oIjeDaPmwWGxmX6aUkUWzVosGxcVcAPHHM9QRb
0DByQ03e4Ywxw716jzJV5tWc5OA9G1laNQAC3Hi6dtukl0ks6RTXVBo0OSzRLFQUHtnZGoRdHZB0
HSVQg0Mf7qxouq3R0c7RnC1IiFqRoYizUMEJzpnft5h+HPlbqYCnlI7xc9brp0rkT0ZWWf1Tgv1Y
T5SGjrEDNA5MV+ikGUNRIylu054h7+LS36TFo7/pD/MHawv5BF8tfW24r+E9gY/cQIjKdFa+/uRA
QVJDwtL9ChyNqqQWa8tX79oCW1JAmT4qVVZ5ZPUqdwVhtr/sSISFLNx+bd1yxOlLrLVp6CN4q7WG
isOvmBtAuNITfryNh2fbrLk7Msa6SJ/jGKADBJTk+z/VTUqax9U6HRTc505Z06xhU+5WvBAulP0/
IHlFzQbkBFts+E4vEP6UsDYr8RloxwJFelOwmDZkgVtXxB/Q/2JGsMqewpeV1StsnWeVn82Upr7a
B61GbuXTAdPLwPaONTeWFL5Y7uk1xl6x539zu+Ra0A5L8gWQpOoTLbnWE7gqfAzOuQpIq/IzvNaf
xPyUvGJk+J2Ja2bfeBI49MAS91ExL9evT/k7evo83urUolbt4aHrmPm9cv6IQ4Nk+tk8mEboVQk5
vZKnoC9TUYrM8/uytm9Dlu1az9xiwynCWZlDj+ZSlqSAOWDja174QpizOvcVOs+VDG8M6Qx/vxvU
9Icsa3iMBgERVXTFONoTRK/FWOO31+3/VPXw0iYHjVUezpB+c2ZIhhcsutwm2AUTjhXhVSmVdKcQ
pR1H47H12Z5jdSMdQv59nmvOP2MmNgYQTpgczLBvrv8qUovbFyB8pPVVHPWuWlsow9TvcHRwWbb8
EE/hd/A3YR8l+hS5zafzWd6moOMWlZ6TpcCV5Mj5jsxIDdUN/YYNNR7itdcu8FmCJoA1Hm43M+xU
pxMzRkplxAAobRBHZL4WT+5Gg1ADTVfXeh1fkKttRuF/wVXGeN9pZwOGaf4mNyH+QnHJ/hqA0y49
itJCbtW1tGBXXw24BsT90WgQAO85xCBofwRVLYePzPO5XXrY24BYJyEniXX1ACYcFN7wBO45niA7
Z/OGdAp/dnpFIx+xZ1RUVFvUGExJ6MKTY2IdlRBnI8nDyBfTzDaTx2NWToZov5JLTZ1DGUogpGKr
xAOaI0dQ7hZ04kIvDkL6SjpZTq3GlZ/UXHZUvBnFIcGocEI3BR4nETw5noaNvdE1Uqb4u/Y0t11M
5SddTkrj1I8uFtbNlyOKxdG4mY8RWPDpngzrtswxWZr0olvQWauffqlVriRjpBpUPhMuffRha7+e
0vyy3KLiIjsrRFmcM39ZpjTWAWPMx7YJ2Vd4oU+PmP90BTGMmpWjexdWkemIjRukhj+8o3UIxg38
Hs6dYPvR2qScKKih6WFsjFzGYHnOcqxv4tU5IfxFp0O8p7fdwIBE1HX9B0aGA3O5pgZbcX5u0LOu
HhTJsV82nBvV0tU8HEi9/GIKS2Ypqwj+ORUBAIKBtMhMvhV1JZxp+o6/1I9BCz0CbppjmuAMkm9D
uP6NW5pMIY2Z+ZFUG5RhSabWw05dQmz+Rcxte485pZF+PLW/B68ZoGkbq0hkIRtNulr8unjfH2ui
Y9cW8fmGbId/Da4Xe7WlmquNNDv1RZwlGaBX10Qf/ispUUShPozYzibhi4Jni+SQelwix+SKeJiQ
GumVJCMC0FU3DCnSAOcWQP1LAOaJRv59wbGjq2c1nwvSey72MphEpqx4OOvOcYnbWq34IrPwBju/
i9zKHMmEBO7Yr+WOrGt1vP4C6Fe1Pr3lcUCCbp5/xmGJMN0E/9pkx8WeizDdA0Jn2C7Vm3hW4IU3
0yWz8MwKa55NpJ2uRb1aOnm73xcPbqj407SjepFyJcOW6ln6FL0Vi/KzvrSW0P5VdVKrjoYdIOff
wAgKITI7gYeRzjqDhfExfDsjeYJxsLhAQuf7qcp3VsPaq4iZTe/IyhrWJqUAKAWBqd+Bn8qiG393
9RR0JBvbYj5ytGlRkRw1TpLbZAA5i/68DObwHgp8aAOfq5y0vin34URHL/qWq06TZTPOFbaGTcSq
ie1Wmf5hu4X25i6M70svOpgDKoRfhSjOibX/mJAhcM7OV+i05et2wah5fmWkFKiq7RCOM8ai4s2c
yZrKDaUOa0sizoe7a0GSWKlACM/+Vjb31QeNl+VKob/fguqFdxgcrUD2WYMrx9lNWfHOjvwX1eYy
mA6dfkqV4xcZaevjxfzdL2RCmJWU5IRnrdo5bAXuwTal+R3WT7mxXwwndbN3Csw0+hWQRyn1nn46
vZYPqQc+3QtBwiwBeAoQcClFM5BevpPB56neGw3PO9DCDZPyAYOjT3ErMd+oXkexJIZLrBHItNDc
qWN3zNugmKj71mMnZ8i3BehCNlBStykgTX9xwXoZ+hz24n0lhO0QgejeZvVjH3CQi/ZXCHP70K15
awqUu1FwZLhRDNc8zIVr4LXPVXrBN7FwooRLJLhIwmOYYBFIa6+Uid4uAjvrDk57A1TX+NykZmth
djv6VD9QP+WNTJoQ120C79me0Ghp7ewqO0dBI0Ys7YWK1sTPCrHLUaS09s5Sa3xDwCjB/+OLIiAb
3L1on+G/t02CXhpbULA66bCHosdGNbeW+uSJ5jyicjFT1it2FEl4mutTUCFw/i7NOiPGZKQgIZKx
QbPidKJhZ25J0gtdODUYWmWjz3EREQ8moIMDrFqJ9Z8RNS8TtiZtbDfJM+snsCvGSmU7mccBOKqa
17dMkIw+cgSiRcD1bIRDGTaiWTuSlaCCxC5GI/TxwR72ps5AkkVvLj6RhMFjNNg90egiHuYnoJov
CB3TIk9XNCqCxcT99VNmSu2GP7VNU1cqOTKETAcPxVC12LDfNCbtSqQfAQeYdnfxTi9OeSsuHCXh
5MFQ54ggKj/HkX/4oYsWy3o32DtR1S3NWYpmtkaapK6UfQwO/D0hT56jkchIGw86wg2QICAWRW13
0Boi+MRBoCMPTr8xydy5cH5b70ZHNwAEpmvtiiMXJ22bTv11JOASZX1VbVCNiqu0K6thlndlf9my
cwSZBuNAgDWFFaA0ZL1CSPo97vCUymVd2oo+JFSq1Qr7UoPjyK3oD99prL2VOUri0RehG5nZaYcm
TpOGh8MINav4afXa/BkGXCh8tdekspQ04VcqVeC5qdek9KjjvzuAEP+pN55El70Sby1pdXxpHZ2R
zvcW7hkAlybTWPsf5AVeZK5D1dGp7pqq9Hph9X8fGJYjzIXuhhe5AST67SfohExE9by3FFQjovlx
hraLz95Fp8wbmE3WhehLmYksTqvPa5dgGy4TghvgLoeo9E84t8GK7yMzyqMtsjx3v2VTkLY16RtD
W9/rNmj2Qr3W/RGiq+74iaZUWf1G3L/75fRILiahNcSB0Ai5f76Hci9SDCufhduQffkJoEQzMVFs
zsdZdN+HCYNsADd0PQkSZlAFoTKvZmV/PqXqwuRXkYCoARMWjIi5dVXGHsXifhrKv4VdyovZMlUl
1EDQ/bmOCcRfYpTEkhlNclwM5s3VDexHHkIg5nCil7B2Xr99ZROq5crTx09kdlhqiJMTEKO2WSDn
nSJj1p7Z4Z/uBpYxJ0LozoyCuOb/dbh5AoHB+hhSyQgEMPXOBnWot0/XGImSIixIlWPpu8d6Uwyc
hDO+vtP7c/lyy279uGZ8o//5DKsYGXM5bGpB2tDM88cSWZOglSkGnDiyrS34N3NhCHBTqE6eNa8W
I2ZIGew9iZWBNdwBnQbNiTf/LhRYV1QxfErcbsMJVnLNSMbg3+As2/xhwkqh7VBJI8O/o0l7Gs31
lS6lhUOSPB1RXIIMX+tYVZAWrY4Gph0GfImePWPpR867USgCWSjX46os4IXu4SDJcgqEhOht83mJ
QQsy+GpQerggzlE6FHAH8c7Xcj37mXfsca9JGuc5jUprFRqVW0usi3BmK4E/2Nm5jr60kYJTb9rm
6pVPpU3hIu78pZMZ7t/hPn8unoknZxe+P5xCrspTqqDEME7AavMAZ11uKjiADe88UdcG3JqA8YuX
MiFC1g+Kc10lTTwNSp+h2GynQx3bJA09H3WPXwR/RF4GasJxdx3b7qbMkyX52PbAsG1Z/raWubGX
QUYkGrMSMp+gVdum+1PWlRUP2/S3tO7+8XNpiiR7qeTxWd5LaR+LafkXvRw8cm6reV9+iQ0pyM1P
fUwktLHOtUEw4Nimej9SLhqtKnfDHJihkHiwomR7ps9YHR5Zz8zSdt0Za47PBVObSVEKzKU9IYFZ
q1zdW9eCn+Hs6KAB0t2Y/11Ddu9YCIHYQJ42PEzuClbRzgxQV4/sW8OhFVECi/6YCu2BjGgT+j4m
P9jhfRDC28ghg9c4WZ/AEJM8W5xoYlcsjJNX6XzRjGJSf/+5qs22MYGkcjd0xZ/8hFqsXMHiExb1
X1eqz5PILhRmJGqmzcF2SBdE2Yk524G4CvUTuBEAUfangAjps5g+8VO11HCmmnvDr+e4CT0z23TZ
kAdwJ5PKZ9Q42RnhWYcCO7h2xvzkBPa+eqd1rImBMv4fDWsGR205rNNTr0ObwvCUjdrvxNzgPzqM
d9c1L7wFQJ9VOCP/iZysmbY5EetirI/XLOsTDXNZj91nnqDXTlZRKcAZ+I5njGUS7Oxe1eD2fivH
Xd4dJN3va0fR5txU2R74YF6uTJmcxOoZawB6Za0+lHZMVPSNiudN3tPmiBma254xUUrbH1yj8738
K6wARiZ/TpIOOkzdmrUSN7FymcwQyhypMxaNVQ/Tk3qFC7e59AAXODA5QaTIICq97jYeBA757rZ8
gjjd7fwyuB9j7vnOI8CDO2BGdi03ZmO6APCT2xjiZOaCNtwRvuQqNJ7Ve9vERJEYurjE7c8q8d9t
1X7Tmr0jZerWiX6IYlpahevKlMB9Pd8CT7FTD1z14sq1csGEil0AiZIWXeeKgWDps8bHO9CR/w5/
MvDkLeS4NfmhMg6G4Giy4hruR/e9fun86b1LHwo181WhnMO0MkcS5zJcI4jINVo/cosl9cvsS+89
pnSPEuuBhu+u5GBFda4e66+vjp3C3U/oBIkTU9PUyZB1oDu1q2J9zABnmoNswoZnxf7QlF0pZgRZ
jF8atLod6k0tOL7xCwUMJ8tXlY/fgDJFS05ILiHBawPS5wQMmAmt8JduHh73Q1PyP4xvL5NCuuww
g85ld8wC2fyaDt7+BsQOCLClpc0ZAU+b+FZnpYgQN8DVNWvVcMBOyatId5yvGef4NUlkb/z04hK9
WSNpjOzkE+x+XxqdeKjtynC4PrnudAYSDPw3aTSV9R9xZSqPQIsv65MKHcgCJ5Hb8rBO8XPSE4dd
HZPBTJMpqTY/GZUoFHdxYJtYquB7VlOtVkELUGosL7+EAW95yPrumO5btamWNuwPT2nonOPYPBla
YcsOnKPU1upCKlYt/Axj1UReiBuOZ1XY8inVLf/gNIKS/0ajXI2l2IVll7vabKO28wQO2L0eepsQ
hPWdZEGG7lncoF4A06YvF8dyYB4sl2wsx8NcKB9KU2RScVxfAgP4eAujPHi49hIzNuXoGP8RjJcU
xFzhCPx1je/AFDciuN7j0vhnGrrWgY/EyQhc+W4FnDZ2rL970ut6cCoJdCAIwOHsjrupnYgtHnN1
zsGv99yuwADUoQ/RqbRkJcj8uO3LEYDpx4bjuOco1IReCdqQorGja2OlYDci2LD7JC6Ix7ei5hxX
CeNDFCmEnzyyzpYEPrfi9rRbMRMqqO/pIyBNYsgxrMsLT1fIqgx19eXdc4PqUopJZPpp6hugjPSr
385XeMPzQYqhGsFO7YH4rhDGA1lYwgv1pk8Op7v3VSEBz8LjnlzbW7eEccKKFWsnulusR4l7jEKN
SNuUEcwt4O1NtdM7RFgGOkJehizCbDtahzEzE72MgSeCYbXj/fsfQ6CKeseg2dFFPVonuXieGDrE
pQ1mzGsyjdNPE+/edZfe6+tlti1AYFBuVGIZURrLPp31RWPpeHWXXJxUVoLsK+HZJhFjepHWiP3t
iPpgcQ1Dqg9TtvsmfuFpZE4fji+4q9Ld3u6r36JUWsnfhc60cEzZ75APPv2LLKhe+wMQGZmY1L69
KuwmFBjgwbwN08veTrMDA1c1wsi8rRZNl88s+h9sR0XqxNFO9cPiylo1uVGxBJg0Zz2+jNb3ecU2
wPhzMF1pfch+vgmB5oWRl2ZJKFa6cmSsOUS5QW28nn9MeI6ORyWPiOjr6IaPjjJpq8DPlG50S0H4
P9KJNHPr9/1KuQ+J4lwdfYSYt4eTnDfJTfsvefB+6URInIaoMjN27OcH6RfHKpUs71TMw0KJp5kd
YI54giNTfVghhZI6ANZ8ONufYCXGSa6y6Kab9V2CfJYFgNx3GtDUzpm8GU6/pntD9aOSGA2pcr7+
/yZjidO54nCrAbFopzGdWpbkq8O78EHIouV/XHXkGq4opOgyyzfrR1MeFbeydC5iab7i0aZ7pPCD
1ifs+UMPzpIbXHtxpaiBvIDJiyNRi+eys+pSukj58dRZRMghGDWD475UftqQRNPSA8HitC5aB7Rw
2i2bG4pPDwRTY9FhnuQXwGLXAjR6KBCYF17n6ucWwBmKsDrs7nrjGVpOSlxTIy4kUOXIg4SwwE9e
9kkKQJVy+Q26ONfYkiNPCIqRffdHznTQFLawlBShgwB3UXTLG3jQ4UpNveP9zTFGOhNv1Gxhp60Q
0/N/G+4KG7kOzdHZltiKaY8U/S9Rzkc5tpjNWlgHLrBpGtd1cG0y4HMZj83tZqG/pr5Zw8b7ofNh
+qa4Dr/Pc2oV16cSE8/4E3qYT/bmW7pYNW6SD4YmlgRerTNEKv2lykY+6CEsGLMWOPWfkqAEYjqD
ks3QU8YuAisbQ0Yp7C0RWZOOgeRkZks6CJNAHWU31cO+copt9T1B/v8fNXhF/OD7Fcdwddr8asaH
0UdRzR7KeuAq/91f2v81TMgTQGEEc04U7PPhvC3IFBKQhe9mj1ZnR9MaOLfsPGIjuBXUXnh+XLD2
ebrzD2PPLwT8Y89UtkEFwaLoCzw1rMryTg9eO52W2axwAxRx9M+Aq2aYHaYNCuqiJdOyhZd/Ep7J
U6RRcghu5jwp/9HDrnqLe2GucEYW3PVQTElDbT74DYI912AoehEFCVV/icGsVknjS2ncMybiEJpG
Mb/5bGOQaU8+YxVLdwNxvJfQDcgOe2D91yYwqHD8vO9usCSjR5dFTOjj8owgohBfzig8UA7EQ3wZ
OZqnxM0LyZnZyjp+7WB3GHoDAGLR7+PAd7JLsUQF7cxTUXMvLJ8dB+GQ0ACkWR152205GcXCaTQb
U6K9y3GP/4IGJ7fIjrgwQ+2wJfsAFcaX9tayI31gZajvcdRNodN9uf6anWF073coIKbBJpQg3K/V
P2DikkJ987YM1gImBclaUCj8WEpGyxksal6j5Wx4oJkcPG0zZZIdh8nk95RdfvPyT8ePs69VQRIp
/Ol+k9Ll8e0oT5w9x3pBVE/4qAxlXFOvR9IwQWFn9hhZqkHmnOSP1sdUUjtoTZT45UYYPI3WLPSI
NgHWI/UdAM45PIvwAoAlm+yb8J2CtF/8BDp46AtgyuVhlup++7I9zxNcgML2eyM3c2hWEu0GVxMe
PMuoq80vU++yr02wI11d5ElEK/Y/L9T/vOtfdUHp5Vsowkw4ZZimyBHPnNsxIYBzpvuUjpkUrYsR
e9CtX0oDKO9ApJD7kFdvbX8SDtPePAX7nqfZ2mcyuN79OwoebYn4QsuLCDF8mbDvbO9/ghCzYUus
uby+KdSzCkJiunOQ+L10SIU6wWZjpI6ycUXPrUhYEfX7aGasWYOeXvbHoMzfW+tKYF2InoBRltHV
Eiba0mgNL938hPYxK22YPEvQXdTttd01u9Mn3jAotpDx0WMepX42qnm0KQoYz4L1UX6Wpj9svppN
gzed+JgC2Q3zNO9y+7Ho6wxbzQv/tEbbDK2HW2bNfKQVgUUn7oM8J9Ow0Xc1IUj8HHMALHk1Y1aC
6rfDvh9fRsoaYklCdYXeDuHOBTF0faDQI5URLHlJbdc4o+secpBwQpSNM4GP4U48RSdbOzz7j/TE
hwdpDXCkckx3qgJOvJx/PVcCZsv/eGa3F+ip35G4it+ryMwy576W9NRr+aDHNuXH5cffDGteNHkZ
4EyrtWsSu0DjUiyQePpsEHtiTuQtZBf0s+zxEOJLpCVWg9CfRtqeHY5aMXqT35KS+RhngEgPD2gz
eV+2Y2B9BkQptUMsaxmOdECdw+sGCLmXl952D/UtYjR9n/6r/TpceAHAl7kcW+6Tjg9+h6qQqAeo
jujdEB2eMOeQy+2i5Hvuq3lYx+F+tubzQp/2/voQKMuXHY4DQlpf5lFvdmec8EUrU4zLdcG/FDEF
xuFz7rWJXG94DybopE+yUdaiGUbwC+GD2yzwtV5bN+UmRrQwdnBGZeT6h4v3rpma+HwUAUlhcQ4p
k8snTnoa6CG3Wc0O2EfYywIqHqUwQjQH8CRL8YDns2o3sgOcoLNpPDge4TH5mnW/3AytuPlK3Z+Y
EKJ8ep3GfQ3KGA7b+jmPH044EdQ8/eqRT0oo48bTYPhbLcj6jUJGA17R1QMvdvoG/6mPZMFYwfJC
aFEqpLpClAS5kV5PYWpIWY4czBRCQ/gOl8uaIi6h1iCc3Pk3cuPFw6Kg/jkS6UJ5uZAh6X5bILb3
ODtCzE5UljzLFNW/xb/8eL1ibJtHjezbeslVxsvGZyCpYaxl3nMDo2zmE3sRZBCvG+aJSG+6uiKe
2biChuG9sNmkJVcIgTNPZwu7xVJ+9tMn3CQJEZK5r2iiRwGYDsDXMuxdzB1qTPgnt1IMOY1o6po7
5He6wJrP8waPoiKz/TXSUHuYh/IoS9TuyFjiEqK0ues52XB+sOtmViElwdj2nQiHPi3QIfa635AE
LRjDONHX6mYKZAvuZqeC/0UOALz0pVtgK+31SW2VmK/mok3xQYJAo7gfT2IHe4wzK1H4w9WUAlPT
d4HUxEJssUsbacFgTsrVIVftSshzYw9RO8R0R89lZD/BNYiTakAlJs9rUtHn3G6LKh9bz++2vqPM
5+OMyWr0uFOxU49XqFDw5QztWNyPGzIaK3tExdq+9QGppdJsoH63B0cAVRrKGdiYhEEReW23Vqrj
o1CqbkcOUlhAyejG542YhSNykijI+Gorkq5fULcO/D5iNf8o+qa9XvJhzy/MGK7C+fSOzHO5e1KS
3VDlYSa98w5m0wcnBgLXN6JSYS4jf683yaz34U8buHIuO8M7g7L7wGw0Lr66Eoh6J1jFisD5tun6
2kSlLufyv8dQqdNN8BuKykYq1sGyo1forSeQelHNaagV2c97gteyau7Zo8s35RoXFUCs/vJqcigw
PUmqe7jzCH5/1/cdmoZcpiT5UGadB36go+oStBcTT7ZvSDrjEYr0kvAzbqZ/HJC5mwdu80peU75G
aqtIooQIJzUuwaXhH6y9gDp/RG4rRB/R8Eu6grb0b+vMY9Bu0goUZaRLB/Fk8XKZN5XTjr0ufha4
MK0lT+f4leUzRGku1kWx5APYIDyu0614Tkvxo/m4sTsTVYXjkjyWi5Z+r/ydf8+u83YgmPBJ3TNW
20gsQAxNqvbVQYdBPhi5lMYTrBG9l0jX93WZ61/WkN8uz0shvOum4+iv0RuFyzJVp6u/GHnvLtya
42D62Vjy95Gsgxc/srfiMRxF1ZXX5vOSEhoujLS+vFGqgNLP4GU3DrsYLhaodqN0/tbMeso3tx3P
1A7XtZ5OuYGf5BJM095QJwJ52iht8qMPTrmcGpL9sDd7vvb3jLLCl3mTYIvhRB/2Y7rh9yUvAIkW
CuKyNXbZCndAURhLtvbn9sQxo2u8T3k5nxjSW7vGoOE3yp1HICveZFaOhZoYU59kICzjaP9V+lPR
p5iwpcUiteRpOM6+4jifzUrezZDf2sCGFwm7nxifUJsteYRtwwILWEeb4valcQWkce7rvXZMRZoK
orlTLvEZV06aNiUZ7DKkVk50+zGGdMPoz1m2SOmiwYsGVB1AgwcSjHic6+W2kq2yfub/AQc2+Du9
a/R62Ung1ireu5vuy3JNKnvby3CnLF3D74sIpg1+oc/EkAC5rAxI322lg4SGR1gRvGOhtFksZ76E
IvK9pu9U3y75ueS1Bi1N3uA5QtbyaJZDm5hpgFySZDBr42Uh2PCW0+phtLSyea8kk8akqOygIt5g
mfHW7nF3xcYutX8CwjxGdu+KND+Yg+TKPO9nDAjZZ6EO1EbPirHMv/ee36K0hJ3WCfqBajJH1QRS
V9ShAj2vFObtdcJT/ISVAod5e9ElphaH2/vgh8VVQhDoObZszFHO2J/4t0yCelhSV0kVLkhIVcRd
lT04uHdAWtx3p3qRCUj4qdvnZhb77pxeGb6nt9b2ixZHzFF8e8y3qshlKviFiMY4tBkKhdPA5IH7
RHUtsf7eeeNlJsd7hAlt+w489MA+AsWvF8i1cnQrWjz37lXNoXkjE7YV1wCTOejVIAAkNwDJfSOO
+6XV4wb180dbkQpDNW5ojLzS6fgiGlzMV4j4BiO76gkxOS4mWW7Qz07i3YJX6Ct7LH9a66LMn33q
BQZFdKEQzt7JTe1An5scvopmHTueu2/QJMmSrZ7Z+AnH7gVk6eFBNjCQSl6spSEtzZBShMqpCTnD
I7/TbukO73R55UcqQhNbH8q5xkqZduRkz2dCjtf/zzVebE7iCVX3ueIxLlq3Qkg07i5dS87CkWDO
45tCACnwVcEumHyyoSQXfZAXWsaIiEZbF5ggc1xsh4pmX6iVLQ2XUvXqmnxy6LUCnKc2XR1XP4lD
bcOd6twg/IgNMboG9zZY4jZWri0jqGUgwVMB+0bASKvaMSkN1bUa3Hh/dW+Yt0ARz7TvZO3w7PS5
Rz/oxNjl0E02qe+Tuf4c1Q4WSQiGCBKD9SLEkgUYA7D7uORw3g+Ms7lP86MpUgpIwEqZJ0pb1LXX
GPtW2WLNfqZ2aJM4xnJD5HmcLYneBWCqFgRfG2hGlCmi//+nyXTDMftpoM5zsTrdLf+zmPcMV2h4
WUxFF1eQ9ZheibdLPvwpPww3vlJUIWrZtwSxfYvg9DM+HONEsuCQ8O36rpz9UEt/QEz+XAXWmu+r
iY/oXhzOTQd6XA/8dBx8mIWyUmceEP+Xg0UGyDBfrqGXhMGjeVAEzRntCeCklL32YAEi/fzXox8U
m8F8Ppav9itQd+sfB6ncSVDas3Yuyr4DajEP/lvdE95nUeCOkX9haDPpknONFMdeKf3gNmv8uhsZ
wHn7QRS1uV1Id4yUt5DsXdbZr8eyBKos9Vk+6oMcKm3etSXBJ93HJiZBqPoKwaxhvpsveUR1f8Ai
ZKqwEjMNTHRvA075B5S8/5BRgGO0izLkMHXe9N1C0qEwd+m74oWsZydBHndZfnguvHhCNB4pSlT9
X2XgtYEFUEXUOnzgi0e6C9t0TfnNBSpwwMl8uokcLqb0pvw/X5l3nyJHx27yxiIV4Ma+I9WzUHGS
wCQUMhLk/h+3l2JDW3biXk0YMhRZjsJEjYgk3fHm0CRvL9URNHI2wyZOsQUqeiTwGh9PU69hG7sX
/pNVefyhz6d3wfr0LbTJtJpHWD3TOwozxDKFa/704ST36TqckIOjDEqCpHubvdD2ggGVciqjSwQi
1rts1Ft56EjocQ41p079rTQeTCIz84hZ0u/3L+uES2i/IbJ7+wbyEpJCAARt8YtpST4ftldKL+X0
9ruViO8683sDNOc9+AAmyh4ffMlrYNxNAY0AZSgwnAEkTlW2V6lkHfmGDofWJERgHl5A+DojwFtx
VKfFIoI4Bx/BAoj1QSHtcOPNr6LTxdqjT/vZF5T/slkvq2xw7WH02/Iiisdpc27omh9ZlYB0nB4Q
m6V33+h2BEU+MNi/KuTaMfEmO+TFajxj+jzte9kaKGUHc2RD9pZIig0tyA5geNLnPFntb81Eph9K
/R7QsotaikpJWNf50TZXsdI4wmHw3DWrx/9QY1H4R/dmoeK6Uiy7gm1cZrPV60lGwPxe1j9QNfKq
jBEz01KZjELSH0vQGXoHce8M5eXZfl1cYZ7LV96oPDFGC6E4pCMPYC7MZhDi9NmTST6PLXU5OoBO
TSPvlXMUFHbKp8GTldgixXRSGeKnEGEerhFRFbQRu58qnNVvp6rTQB4Z8yu0TxSFVLXHvE5LLAjy
HIQGjtvM0sttYr4U/zUEpc+kZNeDz0OdioNqAi4CjS2QIpSTG8HvxF97jKql944+8TIp7Zme94Ox
pSBJved77G1+SnnLeKbacXVrXNBap47JJFnWAZqgY6aJnsgt2RsPlXsUYCU1JAk+ezYIgPh8KNzF
Pypa/WdNEltyWMF9vgH4yKvnQv/DZEDh6A8DeOkhU7PWArTB2H092bHa3q9/nWT50zPusPLCXX0q
0TuT2ph1NMq5aPJVfm7hGT0EDvt2kPURge4WcU4vg4aV3WFvIofvtaOKt32iQLj7nxLa+A3Qg0EC
/KOXfCoFZwjW1irZYl7slS72ZHRX+zHRJVTkBHFAmcs9kDSXHDR4eSsj638RnooyA3af17WpwxaS
lplfXr9OKYhD9v4M2Qdq7o+HmfB+QjQZ2OXW4KqU76/bYv5JlC9jHHbYXVPS7uqxqQBTWJ6abnqc
fU0MAI+gxqNENclD/QrpGwLxrNy2V+IqecyN440rsQIr6ejK9wPdO9Uhcl0z+vhLmvnshQ+DOL01
Fu24XjifE4xAG6yyGFUvIIMvWs8r0ulng/CrCiyk1zcwPHA16J93GSAgA+8Z1XWBETzx4WdPzjmN
lrGiLhfLj6MBl0C6mIlXkXDSsJZO0eZ1XMLxxtVzCopCprXx7ibFmEn3iCwdYxL+n0tgR/IXkVuz
fu3lF3PPoyeKbypewrN+Bk0O6mbnYTCCVeF99KDuL6Mkevb1oPo/iVUNQpLndd78ir7MCjsqf/KY
yZN2/Rp0i2bRrxcP3VmVY+ljutmpVc8nGYJSLrq69z6veBBTyCHZynYKRg7NGVu1w4ZoaRAjaZ08
2ybWpEv6ZcdUC+1dgqRTbU9QJs4d8KeVQe7Xzi95SFIFRthJaKlD9xUr6gDpg6oXVO69fWp8YKx8
UlwDzWnP/CyyQ1aB46ZdQlQUp5AmqwIUe4g2Wr9bjOaYZQJ8SeAOmMJwZz32FiHVgDUMnHx5riuU
W/HA8Hm+GPujsrutYDm91cwKlTPX5uk0BeOnV8ovZZttOGrmA6W0zcwdV2ixPKkMSrodT9UlCNCr
nUAVLe2GO/nDm1kBcdvKNY1596yL4d1j0i3fCnigqjJ75KCvxpEhv+CBntULHSQSRYF3JTfcE1T0
jUi4PJafRtmvgSRYadBSTyWtpksSRRTTLbNbnmr2x5tE6uDgTO/kiXOTttoQmJzdMA6c5wzXXIXQ
C1CDr00wJQmSO3FWSvO7mEOMpIsg3MWVCdexO0++BeBPfeTtrbPEDTafTbSRplCc6DQLilRCanHR
Alj427gIrd2mphPhnieKniTyoeI/w2OaW5iqh5uOynD/2OMIRks/t4xqtfTTFB9r1Eh1JAZiZo3S
ml2U1n4bzzuJgAM+KbBc9sITt1lrgkhTp4kC4XTdiuf3ksDjBGvevxALCe70cPpNEHT5SaBfUpEM
G14LTmEm7/HZqFCxZyVIK/6uVS5iVwEg28pdSRrNhiqMmPoEwukdIdrAoO+HfIO4ZgwQqxhJWrfu
0NYllRIerML5G2mZqRSVYvGrfNdrvbckf34EMeXa1H4sfoSXBZUM0d5Jk1CdoztTAIIPOzhve6z/
J5expLO/R6hZVaqAPmpW3RODPzRkqMoQixiRp5DJ4/xtvL9ZIn2Ozz2+AfvzSD/b8WEuGdaiJ2/F
tVc74YS9Zs4yKYxN3ZmUvx32QdSbNhOEVqAuIAUaZ3WF9/YGfP3Mqiea54CYn0Wg7lXZH1POxWyb
0SL0TnZQf/j/z0IdZX4QPyllm8gUUyerJE6TqpTs/T/F3a5TPpMeBU3rGX0nNOP/gJHLdYHGWAXc
XeWkgvsw2fkuKMhaq4Odcu0gASQP7ckcrXFygLbkjSNWlR4CleoDLy0JHMvZJHEtcJGxhYRYE0R/
/1gL6td1ZGuqcPT1uTsDHQK05yxU1WxdLHr5iZRzm9sHbIY+JpQ7d4Dv+gf4dLvcn368EWrw0L9o
tUaDfQ9e+MsMkcjpXifmh2Hu8+bs97Vuup1kY2i9Z2Fh+ONDF8Z/+Z/e7yM13j++X2/kdjeJufnS
jthWmDPijKhEow7QXgT0qM0cDjng+6IshWi3W3ZfnKaWSbPtVhBcyNxdMauDZxNVppyEnxrhuhhx
3t/bvmCLDfWZDMJSwIfB6XyMuX4cR3MpuDVc3KuiAcY1uexosVn2uYLedsbG3h9CL+b7NTOqzaFV
Qgr/AaqnSg9W7PBFlAB/6TxB5R8erpIeCWGLP/fvxh5pICIQmtBNJ41hpmcv1x/w4pOxxpzQftPJ
TrJNxkb64rz07vm4nxqKVe6FtakqVaOFVzTToYQcwV5ikxrWCEHliVKbZyT6qOLlV6SbupBkLp7V
rNN1Wk7jiBO02C3REwIiv9EsYdAuHOCHcvA/xHI6WkBwFhE9n1J4OlMQ3xp7yoPs5WL0pw6giTpi
Nlj2NWJKMQjhAm7DinjkxeY+tYFn3CvqtcGlaVrWbfiNMsTuW6c4/QXiLlc+mbDxSp3evjg9LkFk
z+qWV6xqET9yTItyFU0FXevE/ELX+a0zrvguiN0//ps1WXzOII7LNZS0h7SuaGhCVBya9b4kCkm5
UhTe1OYv6272DXnNSYggzZnadcbTmYRLSC8DfR6KwTbq+IfoDYNMCJQQ9I7sWl+6Kbjh8311Tj6S
K3sFGfaZhPFHFLB8H3vid2ETO1OkptZu6qAwGZ6/3lwAdy/fS1F5aXLYHT4FhElaDcMxyfH7fZjX
yOl50/Br2S2NOgwQdqh96gtMyQ66tNpThGmDwqnh+O19ADf1s72TWvxkRo6K7z480FZEHcHA3BiV
d/FDsnkrMbs7O+rgDvK0YwGEmuK3km2Jm0f4bP8kvEtN757KTQelYFtormnydIj/jnU4CmI99rkW
Frr/QcRc0qBnioL28oNOBRyhQGEzFf65yCkKOsuw84ammMSjxsZ/SykyBFM4jpYWYmevHyWJqU0v
SXs/7eJJS2MJXvkYpn8/LMs3mvfp+GAQSqTI8Z2L+jIxFSVEyn7s4HuVu3sjMT46Qgxi3J/00Dkt
3s4Y02q6XnSdcYVcJVCDnf8ZREUIYU/7llRd/Pk4+jjzW5sW61WRTbL3p/wmrPeOgI8cnYQmvEXz
vrJuFNSo7ecOWSGyG2w35+YxLC+QDTcmzQsWii5EfO20OMy678dIhzC3/dE1jAAek9AmbxkbHEmw
apVe869/MfDdcpcmKdhNgPZQykYwI/cz775DL/p3K+2aN7elZe2255u66E4xA2wtywb3LqM5pmuy
g6KhUOrHTxXKYxnevxiig/f9FzhLSbnk1AFe2fZO3AJ8hu1bTb3cvHpN89IETqHwwtTBKTvGSaFT
XImNo48M5c5zdXkwEZzSE4vNBhDh3I9O6wjg0tnkkLaBsnHRtZ4DY81x+mwtba58H3AEtUBSdcPd
QiklJIxPh5uF9eUJVH9TTeVhewQSasb6tsPXCnx25NWFmkEUzTy3VRYrE11JTIZhsRh6RI2q8R7/
ArCBMgx8bnxMu0KeYX+PRAwnY1Z5jVzx46+B7suRWnp6vNmGgWXiMQwHc+P4Yru3foiu7t7YBbYu
K46cTbhITyAg9/tjEtAX0eiTgQiryjG0amFjbHgpK/mku4pZzc/67OE4eBU4wf+I8EzyqeEKHW+F
xxOQZqGSK1xVZfsca7i4XHxO+SExC58z+GIRP7ZmniYNe3G4/6GzSrSMzg87i7YHOwDjhWYexsQT
f2ZmgTxahze+vD3ecLJLwqPttkD0TqmtWQSS8//GzOQjMdCAjAbaHgbaKnH3iBYhhLuHon3y7Zic
dOyQIescgz6BKL9OfrAb67a6dOxcIBQwUn61RNsTTXJ7QsXsw1zlXEg9g5BSlp3854i9CPnq6o8V
7P/XWCE6468FKBIK0pTAQvBBLehSubQsFjkqjuPLnabEPI5EvvBsFo6TICxrz77myVaHjfFQnIla
gmwBGEGQkZFY1mgrQFRdHpRFxyyk7dDuT0Ba/TLJfYPKiI1rqpUDckD/1q+A4x4GTmxRQkP9Fun9
1RUeWcEdQsuASlTOqLjN3o5kSjs4Se84aWGlK82aveeqseXDt8n8vVQMHerH4RaO3v4XAKA0j/2K
5OvcCbKe+3neK+lbERiIsJ15Lrxkj3KONFRte6SfpSDAbM+IeYcKQK+7N3FwdzLmTQpgW8jxZH4p
hkZNs5uwNws3EIVCUpid9OLncPDLmTxo5Ikr7EG5ZA1MmVNt8FvKl4+dgqcm2rLDdqeNs3qv/wGl
HxjZLkEW7wOiG1V/k0W5UmI1YJd7NTt1kNrglFnGm5NXgLy7qmSCIXVCoUzIS++6BIQHgGnS9T7z
N+jsW8aT0izOPqJkVwdbcn5L7t6AVjkpnMcFYd5SlVVS2EpRYfaeVLWp0oGQC+lMFEyGK5VgFILg
snLIoGJ5Sjr/B2GwV4cykioJmxWGc4Uo7A9x4NdIEZtOk1YegVzjeH7g1MOuPpbQStUmLeVboT0R
9O5uBiyhGaM67VF8UUKFdca0ZsukNGJheoi+krLqhWZKlKXH8zKEdC7okUN0sFYLgvPeTM+JhR9a
+lL8DAc4tbJeBH7/CYs9Qn+SDKEkbDWzm7aNX7AmnTCCA5h9JQKqnMkPP/vc6WuVjdx2V/F22rxh
HOU7rTIsmzyTRgdxBzl44KEZIEzQJ/dco+ky3C4KAdDLtd9nHrm7LEubxB5i9rWhGoJfXLQzpQz5
dRrxrNxFN4rEt0LPQon8PBviu5a4L9Btnz9t8pC4vTDpVwMvb9tEpZRyt/84rd56+GnFeqnwsdAj
EdfPp95jiYgTnDpGymf68zWGo1ebmhFsZknWMRb4bAcjhcOPeejmGaU7TXhVZh0zcDAq+IPZmz8U
ZdrgI7etPyQL3vnOkoB0rHa27k1DdggTAaggrdKj1t4qzBGFRrTji4PTIHUD0pDzemDQDDoLTOlw
Y9k2cE40FkYdduaYpY90zj4F9mwBWIwEdExz8FNNkl86yzSNdLBzwSikaB010yY1QDD7tJ/y/rkz
Cu5ZBoMT0I6Tmxawx7RsTS3lIKXLHXmjKmItFfVMSDCCeaLeAjaoGLfQgq110dmpJ7+CvBsSpEcn
x4r9TKmoknCysGGE7BGd5iCXDI2zSoNoJ3qgta5RSdpmm4tF47HfVlXFQWmyQTKbSvA6Ct36YuwX
3eMeq6e7jg+kDwytLukYzDjR0oAfbVLkJOno3pclbBGBBT1taZUhTTpioaDNOm6URcEI+uPU5Wix
eDHt9cej50eruMWA2Z6t3n5IVL6Nz/OkHYOZ7RorkPXJ8Xw9/Q19muwIgoeP07Lcqgz0DvAD24Ps
oJoFiXKw2Afy/T6IeQsYmKmCKlVQAqARpeNoPFxGvGKUT8hOXnpzKdunojwkmdZR5KcKZJbJHX58
AMTVxYW9+djyLxKKk0eFlwSZ6OKLgdTVAMFiEnf4P/B3MD/jwP5i8RN014gVgV6vxrISTSxIuhjN
fQfNDgUBgUvAyhuLHFij++CyEbujunPEVVfSnCojvkmhq0bbpZbZDSe5KyAaIaFJJRxdfpcPYQoc
g8GsSNvDuYzQApdh4cDNbRBf26YYMzQFekPLSV0xQ3t6cjg71/Wut9TtchJbe2u5OnuN0zHdRlt3
5xDZ9U7lmIDGdXbPV119So+3gueYj3Wei0nvrtT+8DbwSD4EGBXDQijifkLNgKkk9WAj74FiFgoG
3I8bi3rTtRzqNUoBrmEBEhVPWxj/1Cp7iMTXwnPsejmY8wVYJVpH2Glpk7yV0TH21wod8ZAB6e0x
zYeoO++6HfiPwU17vWwRD6jijwV9nWnUU6kI60+/mKE7F4zjwg9rsL/w1SBtrWAiKnH7qQBC6F2U
hUXGOwAr2ksb4lByF7tS+mRglNIjJrAVoxm6DO1TJOwqjwinCyEqSwQvP9UQwLegLl5BgJ2Ah5E6
Eb02UMj9kcM8RKO/Qup9ugeeUIen95NSZSORFuirOslgQ5Sul2Q2EpBdUMuksbs8PCY186Rhh1R2
/eeMmmN6NBHro5379JD9c8ViGBuq6DFVdGsymWA0r6quTF9iW8TDAt3rWDqKsm4BQPu8sRWK/zZm
v7VyZ+DfMtdvpeFmJaKx4kBqO/P6r2N7cb7iegkAbAYoUhiPpO+GXs/Q/ogohByAhC/WBkz2wRMd
I+jSZGiDZyX0hS702ZpgLm9tWmgXxUM7+rKyfecrjXO0eIJCA7ZfhN3K5SNQFXtqpbt9YADfGjq7
aPG4uM6HQrEbfR5Op8dpRJgTheE9zTgZl286vIvJ68mz/Wv+vG1FUWnbTq4go63eSjSpS0j9+s2l
G5RRx/T9x6wqKvfs+h1yizMw9++8uw61JqcFMio4f5a+6iPSgKZYtrXOw7AOLSFiT9OPl1QUl8IZ
IP5tJvjvkzKJYyvEWThqDMUqIXUYpBdTqkb3PJdKPasB9DNfqu10ACNaVxY4q7nYhsl4WpFk556J
wpr7ANscmDHLwqJpq5JkzgMV4BymOIrZsyLrYIyegJWJLKiQoq/K4BXQj6+tPZpqumzf7vptdaBi
hMiFRlUxO14/wIPqNWU3/bt+ap1GGsnj5bLz73kn/6/9EZo0q3AeP5XDdM+HYqrfAxpiAEd1lxqP
0rO+Oge8lv+qZLk4sNuQ2QYnnwGm37rlg7fIb9QC6QmLLlmACPpOumpBdQCD4WCgBCyB47YQiZu2
rcSXPMbbTCUEwMB7wzcJmXeE0TN+hQkGYtHALhJIM9yRbJvSBLNY1+ZCARI0h0r5dPc6C8vBayvt
aHKpaQlzUaVbZZ65qUMBx7P+sd3lYCPnxdx0FkyA1hB50pi31l3Yrd70qcspI6lDu8hE3I5O310F
CvWY3VDsmUkL76DzgEXNVPgkFJ9mwoFX+QXJrFmzhF1wzFQUpKwcEXBGooeX9Gw93dMKVmDP6Nww
oKwKRRpcOWD4MXYKtMfCfmqrzvPbvRZVvbf03OBy21NPMnIQWJvxi86dxfk8guZ8TX0FnIdOv5Aa
W9kP/TtpzEYPVFEb5vz7qXG43bDYCznXFNNmljlOHi4qPKdP+HCBuXBmegI2uuvAhBNEfYErgVUE
Xzglb24cO/BdtSHoeokRkxUeuBXShUCFXrP53yGYRdTI8iwsJhzE7Tm0rz6iV/dT1QeAVr6W7OM7
Wk7NJ2korbvhCcrjT+wsKOKnRw0OZNmG7eUGgmqaOCRaR7TNBWozx2VJjo3OmsXNw6e9Jt2k213b
RIBGhhZIGQ8ESHLF6om49LhYhHpP+xoma0Vy4ksMUpgGtWUWYWuJ36AC3GG0yJw1GFHE2eTazCqJ
lmFE0Jvkcfya9dw2BsMc4Yhomq+GzonG3dEdOJ781yNT4UPvrwH+w9i4VhOXHmir0od3fg84NQTk
/brd+j76BRZBaPX4lRbeoO0NSSs/idDmsJ8faAh6tNy/BEmq7vmySn5Yw9FGWUBe2uTjb+LeiUaW
LvVttIl++jIb11pQVKVZ92hASkdWiSLBKH7z/Gq8j1SnWkKSRi3pE2cSL27V42n3+eyh3l2H0LFU
hViwlYcPTcz2JFR7Zc8BioDYrIQnP9IXp9okvAbgjERPCFkqaXaoiBGWIOqoPc6W/YdBdT4Pdq4B
dL7Me22jxeo6o5EBDb2S5i0tq/fRpAbcztKRN+WNqc56f8RSu4idhUAHkvQ1elmoTmA/HMeutIup
t5HLIiOcAcVlHpveInqoZpMUXdyQObzaU/oR/8wSXK8DJIqL3Sd/z20jFvYlifH8csBy4dTdefb6
IgZuDiSqTWW4qbEgvidJ6oBngRiiM20hPObYwcyDd2IZaFfZMqiL2Hvc8iUFmmZp05SKpOmv1+i+
PZ6P21yCbrpo7M5kmmReHQULIsSivMNFD4f/p36ECgxBaVjSCHevNb354QCTbInU6h+vTzvhGd6J
O4+an9FrLt6tDjX6Rxooh5eDKF+aGHoNJvoOfIlVRMpR8Bv5beFp9g4RB+gc3Kf2jTUCy1DV13iE
dV6+aTp6VGWi+D+63VNlcnFWVTOEdaqlSceokAna4l2JqTmqnPhT1zAxtjwGbrQNOFGeR9B6mlTs
D+VrNBs71oiboLSAxUV4DMR2B2xZxV+l/a4JEQeR8C3G1dV2oCq2OywMJg15sWBtJGOCC5eGxGmn
xcUjn+8bBAM53QJ9gTQzXsMgbm3vHB4KCggvWtN2tddjqXJvUsinsfzrs+daH3UMv04E87eds/zG
KNwAabR7Hz6bQ+Qva29IOmYKDGaH9ris3fecu/1pFRgA6hDAdvSK7ypMmCKD78hXHbCQTFffHCMI
T6SoAxXOmjOIdG3TPHdGui8OQ0taZ828I3Wq6kZs92KFwVVBVuGGCuRj4aBz4aFIcuoqQLn70ebg
sWDoah6gqp0JJ1Yd1G0o9uKz2HeVXmj8Z8ZwrpHnfkWAlB6QOhnCJ6xNt8+Y32mw7yHFDTV6e/ht
KDs9b8R+XH8Dr+M3o3LXJXKlJBDfIPhJIHAT9kzbTcqpxIU3cJSxEo6HwfrUs4AUaT5htEgptOqk
0qI/1RgFYMditbD/m7Z8bkgJZ1v4gZc3HRxlPcOlWcN4HCQ4wOVBm4NfjmmeXPtwWqhVtKDLOq2W
EyveWSEGbDcZcHklHzxvMCxGUlULfv8q/5jJHMLrWuTj/ynYVX2PpbQpP8f3tFD5ZCL8Lsx/2YOF
CjqJgn7YpGEt33UHLaIiIDKQOhOTu3nQyO7KufnfZuAEzs7pqjQEIQ9zz9si3fy2NhwG/tJkppcB
ThBNZZ9rTPH536q1R9/KaJdxPOQCNbmz5t68fHHPiMEQpXt0JUkFkzxTaHtHJf4KcC4Dx505ejR/
H/kSY2pEeekliYOSScQFGHxEhnzSwmKf+Dj3qseb8+0LoXrrAAnZZlORt7w2J4Shod0cS3JwEDwt
jhOk9oPxXoE8KbTZ1vfevSnkbX5whAiyABMCaTD530mQ7VEK/SCin4yS6B0mzttQu+AsZyfqxOhe
iLwUKlZZJMGYIrpSKh/5IFHvLAzEVmLzPUPVS1NUO4sxXPrWprmeqxjQdLGXMe6TfPTYDolQ/Hma
z6FGMjsjYmeQsyUjgKpzbEFd6CutfTk6BLDcKCZIUL1GgX/ceSUsxJvjmTmpLT9vJ5Q5/niL5/mi
J97U9L+sB6kYxo2WsI3QvhNY+RdFzTs02kYhdu+gAhedgX0vNw/ug5MLV39OBdysjHw7/p4rcfWB
ADRTcMNIUPQ0ou011cHjwfzqaAp4UNG+8L30DkiUgOmKjzeTBbvLYNKnVSyx0200KwtmfkBIRCPH
FuckKGgmn+8mbyBmf6yuvIYgPjwJPtMICRC+ODEtVPq6Ue06T6XiyeqhO6wqPOD3ZjZXh244p0sc
cHpO/dX/UFtFViAGzl74mZZ0v9/AasdhvlIfDT4FeiM77baaIpEDtDF/Umz0pZppPY/i5uWoXN3+
ILRFYM9FQ1SNdkHpB9A1KiZtiSNw1/lrP30NnemHGQAxrlxHu0shW1ksgPH8tEUPBCvqbgbRcY4y
xDAAlmywItI6MhoJlpoUH/zqBt2wbMIrAIx1kT7YUjFRHo/gWWbkZoNGHAIYb/cftu/mObOGuopt
aHYl+yPV3LNmQ34jMwkKleGd5TrViGD2dGowNmvhkaYrqbsmyAi0rKo2HPbnlIitsfnAbiD2iSFs
EJluMOwtFmSSEYA7b45S38MAN6vCewPzZ60zph/7Qd4KS8cWupBQsmZgENjmSzavwBGMe9lfeOyJ
zchpHLRtzqboSc7O91P8s1F99igtoHHYD1N1gNdf4BwBXoO5b0dmTGFjUQiCb8NHdEEqVSLTu8I/
NQH1i23aaebRQVfmsrRmbOfLXLXaSXND7Z8ROSxD6drlvqNBrYDMh+4gXCVZQQ/fNqs1G7P+ORkE
URMXwFjNYPfEjlBjl0elw5iJZy7oDtLtykkKHoCU+zgHxI14K/IKbfXa9h+6hdiD9r3wamhN2iQG
ZfM7z5wDmOw5Own1Fx469IzlMcIxXnEfzYTnCDtIAnY8i2C3MYcOl0wydUwAJ12qBtXboxQkhYos
+CZsbSA6tREpSflppDGE4B0D2tOOcAeaj/0pka2kHmLKEhNwy8ReXz7lr7JgTlWkK8JTCP14xy7t
vQlF7A3d5cEHNM6bUZXX9UNDJvHJgkfMksMynBA5SEYzS7MTUJkos70ffN3wivM+4Jca3uXsEgXx
35cDlLb+sARlYHuN9C3OwNJDE1zThWmUb+fA+QvEhF1qWLeVp6LE3h6gsXVmijKCLYZgZSh/HSnP
1U1+95R/RSjsEodQXaLB0uLEYi1q2s6N5AJ7sjIaQdUWBsrUW2pArxWn/H6XmJHcQ+Z1LAaIauFx
ByI36TUAJDES5WqwfQGaDZXjRUve3HDcAKDPWnN3ScvnE5zFn7Uf2sSJJgzjlnw1H1FkualFhMaI
lwVTQH3FvovtzWSFoBV2RVinxd0+6yloQ4g/ubrnJLa7c9c5gGAzhoPu82sRb9m0OPLLSREs9gMC
u7GRHTxyqWZ/+tag/PnfRTlaLral6IBvE6GM07tSgsnTS2mkeMmaCUcSb8/EjweWJ5iPF4b6oZKc
W/v9CDri5gsa64yhkTY8+7DeM0aiM5z5ShlpZ+l4x0aBhlOuw7YuzYcRmmhPK6pKYfJEnZ1nX/ey
5bRAcqIUHUEIr3+AuMyO6zwhsApaXJyPxYY1bLK+ZpjNpTzNFLSE66s3xJ2yYQk5lETu8rOH/bhW
QeMqq7YIByTiIz14HHpKkWokFLHoqM3coF+EkZ24TRFXVJ+/3/uWXzSo+IHMDtMb9lha352PQtdH
Pj3olI0aPUCBbaPZ0m7JWubhJ9WWujiIhfncyl5UJqZ8NVCm4b8IZiaDHVky7qPyJ/pCLEApcOwN
/iHAdcWxLnPxt1P2canhOhaDCrngWCsTJuFKwT8QS0K4Ts8ByV49m21+Nn/aBb9fNMBgQZ1k/zM9
DVtTPc/LKB5Niy1DSPLctBDsO7J2KerBpqo5Nm8InB0RSLIdlAiF6moAwakOi20hKGqIJI5BTofH
D+S5EANgR0QeHpXKeyhJK7+Ajw5mZgaj8p4RcSeIIm2sYhQbUHRV8WmjhtkN+DBk3P0r2MF7d+eU
iT4kOya2yefgfiBjjown7XWusJrLOCDhNWribnWoSUD0zmyhE1vO6K3b6EPGZ+Pz9fxEMBKgmxmM
PSSug8/d6ReRI9JFO/PI2u5jeXAhWCloDeEOqrNnQKGn5X3y1rgF3KxNhPw3gAwFBRQLkKFaSV+E
WtJqnpYgbdk4DpYb8a12XrRP1YhyhL8Z3A2hIEQ46/48zlbaVYbr8ueQ+k2MlnIvJ6V8fg3/cf9w
pc1VwuiN605nkaU0GwvwJOXtH3jIToWnQ+0dhd+LI8LXDSPsFUaMolUaKd6B5cKPxuQmFVPyY5Sf
oZ4zeCgkDG4ZYxidSJONUmhQ1JBMuMc6Id0gh28fUNagfa4SWk8apDtBtzLnPYFZS+O4x2CHnLcX
H+YDJzL4EXSJRZE3MX+T8qfpa1P1tVXqH4b5Ht/Gp4lSK3cRTRX0y9Sgzs/DREtGBmfgw8n80Rs4
/27eHZMqVQEtHCFv91JTv5yPH1+P5x4KKrgGhmAmOJRprHeY7nRsuYOnIs9vXnQcH8M4aQXWPot4
jRIz/QK1oEe9QMze55l5rvJh8RYRiOercekTopstwtqLDGoSG054btj+/P1NSoXm8r6LVz6aXIXs
soITxZMZNuE2kQT1sgc1TzmvSPZJonARVU+VR4sSwrH9kjSvSekaOylZcnd3jwF3z1AhyTGowsEP
DXf695ewwNh4YF0qckjx3yf1jefiOuC5+FXZP2YwQ5ID9GXt3y3juiVxw0qE0jKonLunu02PI5hl
CRuL0S/+PSwJJnRvlQ6pu825K0hn/CQiA7Vn7OiaLa+kUBKzHcMNyyxMrQdyvztBTBnzl2ORRZH6
sNwTmiQBCkD3URoc3dbfTs9HaKMJkiYhojF3Pcta8yLHUi9vzjyPQuWkBR+3488K/UnTyfq4Objh
Wzvcs7OUVROgNo/leIVwpzY4G+tITLLKlK/YFE72ZyI6eVxVTvY90bDxjVv0mYpWGo3wYUD8Ikoe
gyXT0AT2ruXN92xc/qDnUQBXNrFwUrsXbxa+z1YcPLNugqN3S18KqTWTDCmrbKuX13l5OB+y20yD
DezHX5vE12qjn68AX5aKcBw4keiV/Cc6SupSgYzBgDPISRZXYN3D1YlOys6uxnc4H5chN0ZbINbg
KxZOAAKHZR9tQTUIjjfHDOJz5T0ZVL/EqMWtwc4OrTx2QviKUx6PxV2yUEW+b/Km4BEy5g+fBpec
xeZVD81muhVp4HXltrtYoD++m/y9ROHWfkco4nMKcEDAmaqog46CjnaatUuKnmH0lpLlNYdFPINv
oVh5ahYtikrMqZqN8sJtvwIUTkFsF666aszIFAcGwaaV4680uDgPbxwghCPm4hVyDutUfRa7MTdI
83ZLLDzjmSMrs4efjoq1hR588nlDfzUtILOvmoBreExg/8W87xWaqVzZ72SzFb3xE2dPQ/g6ZRnz
dSMSimMoxgdi0q6bmMbnpvg1lNTChPtNfBaX2cQn2stGzWGxaChmTSd422MttG5e+H4vEl/XOWtY
Jw0zMRFE7eIrxwr3h7IwJNQLL95I8SHYRUDW67c7REqIXqYnaElCeyLJCrh72OAOGKlOTiuO1cBi
n5jyEWGWkqWwsGWCklmRvT1Zv6RYCD/ERYWvuxuL1V7w7Mz2L9Mj9ZX//q+t4bv4/CQ5+NevZSNV
fpztHTW2lbeC7czAbMg+s8I9BpdfTVYOF5SBfRHfhcQKI0j8QcYXWDJAfKTPZNn3xYSEJzRavJBI
F3FZ1+vuaGqHHUN9J5a16tDGFSICVX+OBtczR8YG5aDet5tMf0C6I+HWQHUpQP7uoFKqzMPVajLd
nLAiFVLCxFsZBU2Pkcv/4fZ/UydtjzXzO4hPum8BFfNPfeA5JOgDvAkT7MvNZn7pWYB14gMCRd8V
nKQi+D4ZflvICdySNCcCwjgELnhud/iDUSfiio4YCUNsrW6G3uphHy6cxMfyX/+xTMVc8Le8tLoF
IxvmU3GG0YsDOt8L5DBm7jBSJMB+uqaSSmDhjiEBGq6oC8m3JDlfM9zSJHzyEhnkIqaJoLUBtX7I
5jgVluw7wCesi/ahm7eemuQuqRjcSKlCk7zBhF/lf0k+Zl27FLXa6hTwlu/GoUrnBr1e1QLBRjZg
Fex0XPsddvvm9NiurD4YIIDwn97JQmwpRs58zOeGIi0quWI1NoeBxnLpoFCtl0A0+6/bw4zPCwMP
hiOeYjqt/FsyESiJ6XRDe7yREBYKyle0ijXkpmKx2p3pMh/F5XYFO+1tcmZogt11xtqbIxn/GAFs
7p+BDlGlWuJLuaPD26iU1UMdy200O2T8ecii9ihxDH2+uVTr7etnSKjoJdiM5AMLzUxTEpp2VPc8
nzo7nKe020xantoFqVH8eXw6b88pfH4jsnr/ZfY54KlqgkvKfXmcahdUiBAphLfRBwhFzEqLVVZ5
9yPT/l6FfpdHEl9sWspXsfRTnuUctoWFRRROF7DTDXv87Okejgo/dh27c7mtkqrSyrud0rUddYDY
DRWuctgHhkreyk5hJCP4xgR4Ji5aGg8fsASES6NJdPaZyyc7Vn2ZTLLpASLwzDRxrG6wVpkM1SVl
CSGAS+FRNGrArEukkh00l1iOvpsKadWS4ikzJD1omQYYrxGjE0R9i7p1BKJ0K2ZhLhdQiAVegX7k
O015cjJVesNzypLDdGdI+8pqy5IRiWHL8lUGh/FFw3EAyCU7oSEKICydtxZy6AGUqNeRCKGPwayq
VXzmwg2CDIwlSdhp/+IF6FaEjLRgTqki6GtYXTIPlcopek7ebKmK4v6ioCgxbtxvusW1Ctoe6Cen
UC9t1Uwe2s7oGMdBjChyZNL8/0OrWD9aVAzoI6SxQ5xrpX+AMCNMNYhQuuDk0VBW6fxlci/rD2Kw
T+K+i0z+dmIqwDt+KZBAJ439QSfWEKeM5qnyt6ARup1bxDtkPW6x440SdDAh3guPQDERvGHg+3bc
Ig6K8tu0XcDtOyeqk6gZlVr7OgRChepgWysoVItmvE5+zGIZ1FF4JIPnhEyUlOciJI21XTyXR/ON
CNbxM1f+4m9iD1z21F7x7BwhXDHfKSztai0AsRdS1ZJgoBZfuEE57231ol1eJYLEdMkB8mP2bo4w
RA6AHlnDNw2v4VYnMN5SbAg/xc6wxgqOwvwEm09MUMCw2OQLK1kRXLQM9ZrCmgsAnkOCoj9LBF2e
JcgpAo7FXgDJdvlT+eE6AP5vp+cga0cfCFKLkv6YtP7xRRAZpQjdvcmNv6FthD9z0aSGGFeifha+
UmO/Q+c04i6tR4lYRBXXJtTcCem2gMsv4SM8DIp73vevYuMAOMmgO27ORDcX9BOUyeuQO83MO3RO
eMnwFkqX1yhUd1i1/y0XZ193Jj5Tz68sfPOJ6pDzbMxofcS8fNk0HPrk8zSl3ZX1VzUXfgQn6hb5
ebb8usClrJ6C0xMtTbVtK6zdUePrxZViuaixI92twRk4lXzUsH97D726GtHTqHc0ZQBKtqt4pRHg
GhjcWi4nU89Cy4rO2B/FOqTbhDThlCJt+UT3N4aqoCrdOBJPtwN8BDryU+yYWzfb3KtI88yinT0J
kzkeWW9zoQrYKhkf3yPTej5Ln0y20+rinUH83YuoY/knI18iVWuynrr0P8bIrsLUjvIdkW+0p2gG
NErTtdST/087+v4fbzayffbwT+B2GrtLxhe1fX78AvXsFg+jv8lZaFlrtefHf1nLpHXP1eOXj2Ls
/h7XY3vYG+4toVdLyReerhNdyGZGa0Yq6pj9UYZUW4jQNfIAkYjDLDr20rB/QTr/WxMtQT6r0u43
idc2FfLapUPNZIPPo2ibddoZv1AYVS6uUdXAToXwcHuPEHdRPUcxjQcPDn3Y9cHG5c8C0gv5dFwJ
OpjhI9lzmbZY5g0QFnzrRY/9Ci4MB2IG9urf/VME/4VHlQslz25jlTVs1cP1syqSrSnokH8J+2h8
/rA4g25fbpcAHRiIWFlJedVKpWIjUBOiSl9kaAjjYHlO9eBKfvKB7lA3JKxZpC7/qgq/vrBGK3GS
XbKY9RqIq4Z7mJL5DXHo//llgJohWvInGrt+Y2yzAIC2xqqrjRJziOVlifozT7Q0VvJhR5BAr4Xg
ueVo1DMQ861MrBx+5+jRFDcG2qJ5TjRv7HVoWqtPf/3mNmMHHfCKXsliGf3ArkTtubZ7cSDc+xq7
QMBqPBrVSdx2l3qxBnLLdVIyqsP8unPbhzLWeE3jurbv1PR14ncxQscOuoXUfL6yKeRpeMyga172
vk5IKW/PB7Eqz683/zNyQpIsQ7hFIV2yau4oJJyeJB/Wyysq4TYGpW3HQyhAvykvvIopQeMQEDfc
rwlX4kykB8hzSB/iV0TiL8217zhjT5a78/nZ0mro3Xt7xa1MYcS5cLi8nglr3mdTAuL7xUjq2Ekr
stOQmF03sJIralu626ID1Nh0Mx18g61Kv7PU7mMkVF992mfG7NIqfeLh7TLtniCVAYLWpM6jQWJt
3ucURttP7//ZRl2mPKqRX4WoxZAGZxffwTMfAlQ78s4MEP7BKB+kFwTU+EK5MsYI2eAt0FZIxTWI
BB7toaNKdEbFGih9zTiHcpAR6jUN2ZfhFQfjzYMvbg9UCr02FQHXYSX0/cg0tHi+E0QVEuRQJ/Vm
Ffv4fe3sWiMEK01Q7D3gTcUm3fs5OsFtshINQWR7jHREbB72ir0UUsxMcRCcb4AhKQjqh2/emxIW
+ZBASa3AZCrwczPsOUOoDn6RoKGKdPUnJzVWFktFR48sjbrkslznC7EJtQUkudM4mWgk/yvXQqkX
YrteEJXEIigEj4S1Mv23Pp2fCv2b46OSpl4xy3k5r5i4GAtOm4FkJYYxao6UaCp/X/HP/mgUBupz
HKVQgh76YxO9ueg+IFTFZ7FLodfotm9Xi7k4TEDf9VBUuTGZLJgd+5+Wlicpk4NdxpegSuRj4f8Y
1iH8UXe6JFn+X+nBGBthPwMhZsyWYzoJ6+lCtryH2uqHfmg6HcsZA/y+1Fm3yfFOrQrR4RSEtGY4
ppKFvk58zBGOjwBHb8bl0pIT4TB+aY/1Xl3dt0TaeMn/IyTJ1bG1IW3VZpKwMjcouemkXt37sDrE
fA9P0B4/LHrjoYj/r9EB1nyFhi0qYHcm+htDY+EwJ7Vmy3iU/veTk+8TwuoJkPMIiIpJFS65NwUr
YwymWgbrKImesJOGmpZOCvJ3qqxNMrlU0nB1J2cvlx39dAJvopF26u2tjNWfCAm3Di125k27H2Wr
WHUcNcELmwnu8FBGore4nvvURykfxdTZYjzODwHnxwa3ig8fDzd5tf/zeVxF2AtXDibTMsAh46bH
vCwFzmo/FrQu17vqORfGMNGlv5rmEXEwJCwzY97q/kbSp2f0SePZ2a/Ab5HjQpo78f+CZKj4L/Zl
9RDxlYDVO4FrkWhE7Txlwa4ZoRaiopAag61GwhlxByJs0Vb7GxdmCQW0aPWSEvoZCTT8o4IaS+h9
PX27UyWk8bMiZMjssRnrkjQ35/ZtPe0mDJCzrO8LgARGHVU9s171DBKR7w6F6HFodmVR7iGZOUyK
Nzql3DwpCQquUFOh5nEXcmpFt8/4mEdmnG144nj8fAcnJ7Tc1nWnU3fgWQ2fE1yDp8BCjlPSo5Xv
KybaLiliN6EhAR3U9qeDOhRMCGU9P1Bv44/2S0gIrg7g33i+EJVRXr9056thiEC1VUV20e/ulPhZ
6mWYRLR/tLGHcnfG5oPVtI9zuVHpsWcKXHYwRq5PKVRhsOVPoBtZb+Ufn9fcxXnsrbWmE61TQhy9
eDMGfg5qcoczr0d+IQ7AejLBDC6hMqm0qbEEBH7G7VlcfP40HVL/cDOBwvV19QxsCSZBDxw2Ixv+
MyGi2mJVAY0aU/6KiPioo75VPdbNZmzHLfNZMrOBHdRt2UCLXete1Pwcx71NUutGjsHrfC/SaRjv
BJK88oL9+Gv5Nf8r5pYvJjERQbQd8xWBMw1XQ2k0eJ0qt7+XEw/hr9XtCT+3Nz8EJ9Z1+wgFpHeW
+b7EqlVVokMd9RZsIcswZ237g+HwYAh1Hzel+Y0lNLNVa9ApXg2gnUI7F8FP850VbwgvACTFR4Ja
xuMyHGLnrvSBNKVa/dHfcoPWl414vaCODwi8X+IYQMKuMuGCPeJShvUS/Mr9tXVCWAHnc2W0Y4n5
j/aRr8P7Acg7xbvseGcw2h2rAUYGxYUAzcoUMJBX1jFK4asvDlUR2urO0XgUQlUv80pDlotjgW3Q
yg1e8zU3J4GZiL6PHAFbjr7Inruz5De4U0KU3JbSM5xJvQseyHmPYP0JfJR1d77IuQfYkECsqIDR
zfl+2fKBBzt1hXNmBcIlrUycFovZQQQXwf6Nw3LwQBVTmcYQl4eUdLQ80BSVzHbtyTNeOG4NlLlp
VijIyERJJwa7VCR5nP0E4mNkxF08oGEbp0gvX8nra9XDftye0GDCvskEQTh1fzyNeiklU/51+Ac5
TMqVMmDvt9DgvJ+CX0txp7iaol8zTmx3gsxcztlBgVBSaOIt2UFlWFFdRRVpwHacTt+wGmZYFZk+
kQiFSTciXEs5feWdilxWmmhfGFoPZbXwwDSNf7NZQkrRkzj1vVdNF3noJBpxaTB1/lUR6fD5LPKb
aARNonD6+GTBHLVJqxA7P5jqMX4o+sXG5LzdAatm3qGwg9uU1LyY9rczEERJjO7yeE50knlmmpoY
TB8Tnv68sp9b+CoCdfMZKIlPy6tYasMKrA3xLN09qROqEV9BmdAxP4KiHcjL9W7sUWqyll5Scsdx
YgAzvLzyN9X29SsXJ5x7IZfbjWjoLn7YJ7/ejPJ96PYPZpdArkUOeinXDxaBruCB+Ok7+zmhj/rY
JUfEwc/Qq2V9/gQdrVzKvZOqlT/skcZKAveAtB2/D0lW1Ii5R+zO1mn6vdBIX/hh+VClT3UA/UfZ
s+K/9xnGUhx+1Y50mUh3+4UVqobqRzlV/AfhoOS/56uzu3zlTpPhlsAL+WPddep4VmLCVV7LYIwR
BnyG+oJUV2bUzDG3qRLCVWRQyNcpfHxZHosZ16NxjhkxK8pe3/KVn4a75kmK8QeMMsLZMjw16kNY
BAQK1q/Ww/Lou/sJ1XY+cDEiQzjaILG15LGg1YyQKqMFrzO72/bDyuDugD/QZtc8bF8OFs0WQG4F
9mMw364jcL8RMFrmbbemz+VJI+OEqLiHLgF6A0bx6hdoaFRu5AgYxtOaGRmM/3Jf+4cuJQ2+7AUI
Cgpyg8wf32tOB7enfB9ZCs5zAamA4meAu6DM6oxyenS5Ug4No9uoJ4OdKH9VvWFbglNcuZlSNn3F
tpjXHfIfQGHNe+HInBq6pPnrMU3LP9d6AlrhBrhNlZhvdeidwa4dlP+65tY52YfIoWqcae7a/dS2
DWJNLj8EtrnShPiumi86ezmJCz+ef9pGXXBivoCWPNP3FspBnl7cAtbjvJfIyX41AlMdPeoWAJu0
UmShH2MWVnyPC1IQfXyfHanOHDImRbPit62KSoQwqbUFsm0BS9erhS36DAtc1xuJqsyHka6rlkVD
t7jyS8rxcDqVStOwL4BaseLW2W+ThfvXGoRDoVbjjvQVaY26Wt559vo4cqLOw66il3XI7TGTgdBC
xGHlMsl7Wy9wKjLMoTxmiKeeKbc3b/sDcB5+3u3Ha0biQzSvlbyYphgXg2+LUaOtvIJMQMhD+Pff
ixdmqUTywIUAmM2Bs2gm/mO4mps1r2kKGVEQwxhrx0h1KBMrWO8QHHWAbxAX+hhLwpggnYlnU6Qt
VLrQGHKYimBt5rGJqcPXILCf7MbJVoOtXtOt3WILro1cLWzG7TUEHpZral8xFC8xgXQ/GcitM2pz
nzqhumVEGVY1L0xQKQ4CjsZ8mv+PcT6Ujp9ev5/3HGDQabTr+HBSdXv2rR3nKHIxvgmhkECYp7qT
wtqvSosxjORXUWtpAtjbLOWN46RaMlxkT77AGykP53ozzWninrc+dcF/i/lTiaR9Uvbd9yvsvXyj
OmQ4xgthFJfLJYpzytTVyeRJi6kw+CQpRVqqNSOC7WeEknS147xpWK1pUnoWVUwzoJ/ai4t/AuzO
iJXs0LmVe7ZH9YaLrpWuFzjwEZyfAIQSRd1T6//p7HGDjh6R+OBebOWrQ4sOjk00fUVgqNESLjIq
xUxWG+DrlnHJ9Rpcqp5Iovrx3wnE+uKXa5Jh6AC0yJjMtdxaVNeetLaZVd9zV7qT+YauxL11wIWT
GNt/Xcnlb1uMSdBfE5WbrtDiaCYA3JMqyqVTNbAJ6ANpvEe5P8bkI/5kz4k7yFvs3d4DjmXhlsgw
AYZBW9+6GLDFLRc1lztG6o8+EM7c/dDawY8IF2bBjYx/8VOax8wbigloEdTh0ohGocYhu3GqHoDy
aq4K1WSoaeHfb2KhlbUGYaOZBziGgOUJadRBl9NmJBQI5m2jMVvW86M5qJegNUWDMaj9sP3apJdC
MUgvawxbDrqYIPxeRhomqm9REwnWxKqCHA4qTUKseqUnSdm0oRvjyusAiX1sp0GUv47Kwa3vHIXi
bcNWh6pJR55tNyvaGYR3TM4vCZbecxV8Jn9Ad/iT9Ot1bFEvxQS4HZxiJzdrD6CpAfnJwQL3nh9a
tOSfdMA0mH8TFsoyca2J52ZEm/i8uiNCPkTQCdbb3dSCvDHGZPImoqavmUqirfwpSTOJtwaJasMk
up0hNsqjvH+R0RiHm+YUKGVEAXuiLpo4rCToRzZmvcxjj+kl7Hbwr+SXUhDTnmjFU4P11PnUeRwp
sZo0+Z857avuXl0beAi5eXyLVw9P+aYs7H7rhudqok+FmwKpzX96BfVMDwC9yKVjW9Qh3mK1mJBz
yUHuKbkDbL+aw25Vo1MQenz2HSwZgket2cZ0m3Nn3UivWONbc1ld7SAoM76220IRAWxOCWxwYjNn
5Ap1t6n9SMp0yMqsiAXVnK07ipXDffjVrA5geavKf/s5LeSL6HF/dMMxgTtuSFcUSUu5PlLizfro
iRkYqGFoxtAbndrMNuitIRFfzvlh7yRoqB1CT9ALE+m9M+1h4gwVCodAw8RevpwDLON3jXgkX0FL
uMeQO4ijsrHiqX+imjJKOutBOe+zRhV53mcgQsbJinH5OwQZ97aAVbI2/UsENkM6z7t8veBq9diK
dR/8sGXWres7EfzTd5lIObySnb1BXGt0aG/0JwF9nifISxZp8gJ2VoLy2oU8WfsJlcYuxPG5a9CI
sPCORb53Up8Q8R83gvzGFW74xXq3WPYMCmX8/8yk+ijfZ3Nnhii/ckgzWyV6cYtFDdWWu1QC+41k
aew82kiaHRqxN4gw9RM3rxF+BRwFUX3vzqOdX49Y0oWbZnhlECRt+Hu6tZ5El6OmZto4nHxRFg/i
DhH1Ioiz6mZjx6Gh5Mghyift5IaT9tGA+p03V4XpWCZMG/G9lNvBYUpaifR0jkbg76Y9V3cZSjvp
op8AEeRSg5r2iG/MvMfXPA8Xp7mkeqfpooR6r6mFRM6r8VpyJH6FbreJHkxt0o7yVfJUQztL/JB8
YAe8E0Z3O4sEuSq31D6pQ8arhEapSeGKmsc+6A1eHacXy5C5HymUvtYAF3bWiTrrD2bNj4RE6LuA
XIGef6uFzfKZVzBQ6DBBJIRT1TsDLT8m3N8UhpSQzejcQ9wmazNACBSDKDEJgseXeq9Mtd6b8mlM
jievTopt4mxZrf3BiJGojIdsAK9v6H+6BZnwa6sTQVYpqy1NqP77ZV4aVFAkYXXnX7nQ6qx+b+gp
6Bu6+fd/+747p7AbdNn1wRSYMKJAlrJbNUJEbYJumhPebt2L+SprpakS+JvGKH/IsjorQ4ZXwgs8
9LCT8CxAwozYnKg4mmm/0r0/HuLhDslUJfWtZFsOJ2sRYmaf9Of9QfXclPZUa2lIp/yZ8T6Rgnvx
uCK5gvQSJDxLHm4oyUX0louh/r71aSXxGQKeV61LZpDOkbRs5PJ3QMpKjsWfV/9uaFGJw0w2wTUm
IhS/4xEbBKzaCHHGI9PGQ5yb3xXivalKw17VOZ1CRtOJxyFzlM3X2lKOQ6+olgEFhDoXdEEzxLrW
9qVm3G1vzdZpUBBZPpsaLSyAKvscsTd6RdAqsf5RiODRuxwZlhIdDiso/loCCGcna1XBHmX8sgph
3jkLvmVxQ8tp9s7MidplXKu0yFw1rfwKRR6w49GtEV0LAT7hEIUJInyJbYjweCDD7kaJl9B2nE1t
RylO5QMpQ4elFtlOnmHFVIlVcbjeWrj0IRy7spjFjN7+wcwWai+TPbA4yoj0NadMSGyVZLoZqtHO
qEPX0AeOa4yK/dmFSk/y/E+5jth2aWNtPaQzONPW0mFi88rqeph3N/VSbEpHKX0B1WPcuXMhLkKn
s2/wpmzSuMC247CO7HH30ifjAVTYY64ic4liTJUQHc7Li+h3GBzei5OlW5k07Vf8x6mGEDDfsIGj
lezen1Es26iLNcQdowo5Jc0zLlee8Qk8VwrokVZcZflS86wLa5TDDxMxP2qwz0GXK+Qzjc6kpzw+
y5ZFi83ow1qyGVwRRRlBwKE8VMFzjJjVDIPtNtCPdxGxo6X/5wgLj9QroRFpiXXyt0BQhfn0FX6+
o2r9F0uzvDRbI059OlXMQMouwLTbalAu4GhVrP1kBRp2AEl32gUrWDZDKMRjuIX2Aky9AS/ecKIj
osLkuw+/EexW0ghmXiyNqp2RzeJeNTwjlO00e75Jl0CMMgTCSKsHZIkBvreHk8B1Ype0EierwodL
VPkLBKT7K53JeKGx4ChOHhu4zlgFrboGTsn7GhXmoDkx2XNqEbIDqg89+cwDK9Qeq1MDiBjK/lss
Ef+CciQcVXoE7FaPo1wK0Pw7aHqgZlj4M2SDgtkpQHvH2vqtatFq+ZBhJLgHzlNVnoaPZOBCGo1I
twpXdc9ghpwpcl0yFwCwy3QrayRwOm4dFWLn4c90suvoGUzD9dAkTJyj74RyGj594fVgTPdqAlGK
nsZpdDuyv5j8M2VTrSAS1fYxxt49WScmL2cDoWNVG2KNYf5cYzkfWlFYYupwK3q+rWP/hISz893B
cslGzxSCI90OMxu53extygWqRAs2v1jHyKCcdGpNmcNZAsCrqTmMzcphyMY+4gfw7hK3YwNiXazS
LpxkpBG4AxuoKV2pkPzpypAqYFemTqlGsMjMKHLAb6br7JuR2WX3Bz7ZmwnyA/7/i34qoGzQIu8w
12Q2UnPZwihgYZWExR2iBRCkXOarI8opzp7dr2jBdNduJmoFnqHDAUj6W+wNt+RME18qNYQpkyRp
5rkNF4cRrDL0ivks+AzSowrT3x9MKPumfdQhexPbSq9byhila+LEEjoNwakAvU8T9vWmImRj+uqB
Qwd0WyhwdPseckvOREbYybxMlM0ha5uzNgt523H8y23Rqjx4HWcFdOvkWY/0stbl6qqoaQKjV5jx
nNw+Wv3LOweC7EHo3+MOfcCtLbcyRwDLPDgtSwW0fjagHt6f5wiIcdnPblQaqAbhzPuGKsTuM6m3
xuE2rXV08EvqllZkrbe/MWq4z50fjkZUGz5tjdlvoZ595ZEZuFfmSrp3KNF84KWruVLmyH8CG8GF
yobpLm9v7hOFBKC3/zFR3h4Dic/Bd642u714puzaHUFTIeCRvIeqHtuj0JALbU969UhQx8CmF8Qn
JfVAD48Z1TELxgb4P0u4aA6OfUF5ceWalgxLiVklqcqCbVy5zXG8lumFKIcz0vf/EVTFxYAeIEjd
SPof+1UAcinKZls22xbvH9tW+7YkEVkoJBPV4avorNzt8iytCAJs2GDk8ixtxdMyUPtLs9qIjD+3
WqpKztWLhtDJQ+hmFMgO88GDUjMDrx0FKqT8wuIRBAIqm2m36O+yNJZ6iwMN//21ltcCTc8ol98Z
cwWTNpT9R1X0u51H2J1YKXS8J9PVk82y97elnHrbR4i7LWiVMMiXTTQpRm+skR9a2CFVjyPbmZ3R
ajQ5C8WI/dD93UeTlTs3op2e0BNqeZ2OEqSLwBpDQu1WeOzYuJdUHJdpY+ByZBdWDgIWQ3Z9LfDY
jFK0Qy23uFnrF/kKz4WE1o85frYjktwKcUzMeU6dhNgve379bNw5c642yb4RjOb/sBdHKFKoPlVf
Psexsvmfh3TeInQORWjM4RI3JsGvIboKyO5QqsaGyijkDx6aVtoGQu8y1FnDpgfFUV7mh1TXhuA8
0btfcGq+lnJ3ODEnXZPGggN39rR/Obn15Q8c0Gh7vE7SXo7w0eushB/tAtZtbqsvDDMa1GhtF5QO
d3z/DVRXsJFJmaj5gd6r397vSL5vs95h94+LfyACzqZ5coQ4tTQbZk+3o21y9DEJNs3KjCTEmCcD
QYMrvZdvBZnumGYVPWAjwWe7QJW0FyEVurj0KZwqg+MDEL6WE6xal6+WK7AAQ0jECP5or6hk5nUD
v03PcIW/wo1BAyFF+p9XX0anJNcHoLEUnkfj7acz/YpG3MTYW/vy1c1h7lPgIo08cNaskjzKPAps
prIdteS1ijwwfiRUW6LqZd28vQyqFp6PKpvLDFzaHBM8THBb37uiXrVwJM+Hj0CfzgJWraub691j
5a0wUP71k23hj0IGCJ7eL7G9NtCQ1O4hgo+/zknHWa8USKWY6F4/fuHUe/d9/7ZVXC+5C2kQ14Ut
YXCBe3z6WeDyjzesoNcdHCkf3gspyn5MNUGI4LdwoEJUmqf043SDvgY3REUrkYo4CyBOQFp/D+5W
TzSfkQSfZ87ubESliQK2urtc66TjyoUo+8LpOWW8R8AFT2PqE1LB41IywgduowLAeUh8R6JATLek
FxXbYgf8Jos6HBVZg8XzjS4mPrvoRjr/NfelTUh7B6J0OpTZpVHo7v9rq5obqaDyJwGRprwusnAV
tY60k6jeCteMKltUi9AmfzVvJOKz0kNq+nb8xRVI5vBJvahBy3idRPbXvCZFRyXKQQYFxPWET9iB
mdFsYzPYWOr18Uf3tytX2lW8zbUz9GwNfLNgfluMqeov/n0TbAKNrOvRHjA4wfS5zhGq6xvsM6LE
BCr4W4fKDXbkn3u/NTNvvcKV0yrV0Vp9Edk8Hb3F+esm4E47g+U2Et9k8qO470bkf+WPNIq+kpJH
7O30PwclTHhn5VZp1RTiUHJOW6IA6zSWmxbn5AUzizmX1SUyXUEEUjJmsQZK7PucnyvGmYC78B5O
gqiggc4KaH034zdxLwYVbYgW4jr4+jbQQaoCgUWtzVxlRd2vKEkcGylIdn3iFBmHeVmQtWK7UdCq
dxpop0ASyDNRB/E3knkQRAnc+CFLljBYQZ/c2hDGXSkk3SIAiBrnX3LaKyYu6Z1ZC5neTJFgJaui
jFCtZEVNY0rq+m8wBuqJqfoJUjZNJnjbbfTYe10uXhtHqAZ9ZzR47xk0WNdW/Tb/2tvG/eOaJNg2
KFdQkiZU/Om0ye+7xAIzyB9H9sjNWC1d0ee4jLwBwX0Lx0VvC982y1a0Kz/bdHaEKWWBRgVvzI2+
YnOPNzvDFLUj4yFBEyA8tHn/sa33fy88lRmeaeUV9WL3t9PAcsHoYaz8yPsTmWe59RLbdr2JTP6n
pCzhDAwQvpKL0VK60HiefOFyNAS8yCq0ol0YijYPW65eS2yls3zgwe2sOroxmjD+KzNbsyE1S9vk
zgFkeoL7gYIkR3LS+axzXJBxVkn13vn8yEknHoJM/hhdZUFD7yo3U8f7O/ndT/EToVPHzFAaAnqj
CHlwygyPwlx74lC/vHHVNpqaE0bzmPZifHKV5yXePujkYVmQ8AiWdpJYOlLdBroO8p234EayHI+z
dvd/N6Y2qtNCITwoAMeEzmcBnmkA8WsXwJWlxI3bzihLR9h2kqyyeCOFJzCi4nlqjXv+S0hVF/mq
YZ2vnH/xEFI1zBz87HWzf+2UzVtNMxp/p7WBNfx3vOK1WsTEtwNDBOOIfYGN+an0ftJh8DpF2jgh
h0Zrxoy17SpRP/IbLqtfXQNGikApHHGvm0/huUGU1OKeIVQzQxAu9UJFAzwyyNzU55LrVi7kLqTW
1m8schDZ72a/Dh2QO9h3GyhpzQxR640Dg6t34K1ktc3iU0yVayKKrvs4QNAEFtfh8Uvi+dreN1J+
rimiPbrlsGWidX5JYTg12YLT8sdedU16G2o7LAo91UCcypHMFWIDehcJsWJY2dUnLOvodKBu6WPX
dD1ndOVaancDhb0JoXgXmVQ+NOs3QZ9zi3jJYZjScM72aCcX+W+2Esa66Ean+nmIAg4KRNFW0j/X
2n2sk3boW9rzWx9rLOT5Wl1P/fyz+dfigyQsWc0Us/mHbB3xMhzuqHZ/+lpHIr7ZC0OokU02ALIX
7iSqjFlQCQyarjVijex9iPiYm4IItFqs1YBfg7MU0YBzY8HBVujxTVmMRv/E+4ImFOR8DgOvXKO/
Sl/4xemIpw9nC0xKbShDAgrFq7wV/j3OI5C2997sszKQ9DdfzWIz7U8bgqoAlptd2dmLYo2jtAH/
+hG0G2WgKcx4c64qcws64uTIxgDz9ZEO2p9zFuucKTeSMN5yZEml3xw93HrqKmhdgFf4/7gdQZvD
+BOBvzVVWAlRxjO7uLJm5ezId0gUn1WD4iDvM32uBS1qXycma9bFyzS7ZesV/ACDJcR/l2UcMrmH
x3CT/O3vtBSojE+x9VV8vUxLjmI1prLQPalRgPcffs6Oxq8eSK1zARNiK0sF+SbbyqGs7UuD7D6l
6vcE7aLnNrdjtTcrrh9n6iD5ZSrdDnvRSDgz5o/ZdKcP2Ka1ELI2wMEaKP9SCdGfNSx3X1IZLHqV
rRx20H+NEaEJduz4dCL1Da5VlH+tViYsjTqEhtLssHBH8tNz0s+EBXy4oXALwq5m4uDKWaP2g9s1
d1fkTRIHWV/9jBk+F2u0rwDxzRMkZ68lgoHfTibJswPFp5spstmVBGoesyHeXhKYLgwiZEQSoxYY
txlH3Xzkfl0+eFDt/qw4Hq/zsdFGRsax8mTg9XlOOBO4CAUgVolS63RkoXRKno7ZI+p+kJowDbWh
z4F7PhtXMqVnJPHzHgikECPP/ZY4Itgi71jFbWYNDHsnJa9Jg2rbeJ1RX7sni50wCiKhHpzDqrry
nwHAspPCNNe1gqp7ITfc/ZE8kbhI0xjWo18wqBr0qAzpSV55aYrfzaTdfDVzR4wvuxVqoCSKQ6Rk
Ub69qZW+qfiPwyvtjNUYIwfKmIds2EYEa0XTZKXE6EYRKNcCHp+0adOsRTEHztO68M6ToRLZIwdh
vfgTcAR0w++xRQQBeTuG13loCl6VsFQilCnzhfQg+cCfqWFocX2lV4BI8fD8JjWoq/n1mVzhG7UV
NGoo6JOqL5tsHJvHzsVX1LSl8+cf0qn1oFmTkTr62zYNrMOPJjI2ltkZ9fEAgnVnFRdETxGg/Se3
YNfcYMQjjqF2WhnuDcZzjZS5WY6ORav5LLOG7tvdpeaA+5Z3jDcgPDDLK7nXKMT0voP7sosI49l0
uK0kF+rgCexIQlbYXs7MCsKTbtx+/f6+D3bXsbJciDLgdy1zWaGj++7lDruFfblt4v5VOtMDpxTI
MYhX4X1ekSZCietq1iZw7A7daTpKxYDEXGkDBW9ARwehMigtFE4f77k/slEsCONTXwYGlRujq7eh
lSSBuBYCTaOqFlsalr7sqihgQSOm9JD96VyNyOnYNiNb8zEo9Qm3msNakHq45uoY3J2gusNtGDzI
Cti0iNnsGFphzH3HEGnHnPNaHqKOWGb/v8EiP3M9LxgC1I3dWeA0xGOGR91851T4hOps9QZk97Rh
qoptCUfEOBaurIJ7tL5TU4g2w1qUJTNia8aDjZz0a5nSrkv1MPCmdMJGM4f0pcebgvY5kIL43elf
P2Ve3/5F3nsjqlTXAembndUgDuMEnSajuYFtkH0egEUsIvwTOxK3gKsu02SIWa3b3tX4CzDQB0FB
QB3S5niCAlAa/qSqyYckr6rVJ+MNiSmaUIoF8mtXxS0ieiAFo8X+lD73ZXEHwT0STSi80IKrYlce
BRe9MkeDXjfeT6mTghlIND8W7Q8F7woKUWSgOsun5fEMAUlXYS8nY/pLrVcsXwAztkvB5mi/ldrL
HK1PfXepMOOKWf+G8VYdg5SLfFZghpNgWlAfcU94RKAN0G5+Kmb9tZQCV9SjyGILCTmW2G0ZM7LO
7E5YW7WGtl+j4nvom+qqrPxvX9nkF4sv48wkc31bc8KOlJ8N9H7UI7kWNcSS/6gR0oA1bIjWGTFQ
VAuSaMos2rVO6+Y42ezn8wlYywFwq/yxX2a0KNXItqa+umKtaYDXkQm2unenDDCRoWtcfsV6r9WX
Hfd6f0u6+09wOvHFIA8yRljFZgtDrRl7cayOPaE+56602EeoAHaew8arMaVMe3vGq4un8UTxY9Q2
FE3uv/NZ7J86yvaLhjNUH6Txcy9UWVJvbO9I2ZVl9VoMLo+/59W3vqOa4kJxD87CZL72HPPTtdJv
rgwGFOZUkeKoMGrzBdufj59G+x3T3qghE/Efm0ZlF6XagsxM8gk8m7KGkwCKwmgjYKGC+IhS8uWE
UZ+vyCUTCRnTyJTX7hCPNNlyIDgEivBNXEoUDPRFNG0hLM05iPAAURMz6hvRDroPem6dOcsPuYKx
9ZEmrJHioWYyuCrPD2AaTpOIdiuxl19k+JCpuhgIVglP6VOxxUO/sqtBrzGgsXLCPQpq+qszXvJz
6Hd9b6ds4w2+YKyz/4uadhx0+ALhpO3yo92KeVYEJnRedHp/sO1g/nNDGoJIizcMRY6aKwGOxwhP
jw2w1kyb78v82aMKT4ymMSgzDsSwqtkjwzq4z/w0HllJm6OUtaQta99goTICFl0YxdqsayFsbnBN
E1fhaGky2R3SWBpuclGo8THjrOVQfzxX8YdBduK22vAOcwzvMu+Sfxtg1HYe9aWbcaTD4ObUmOJS
d/r+MrJRA3gzAZk476IeR8rRHtVxDfdrbqCnQiRuZDRrkDv6WjrD5oYGO2vKYYvoTbZtn5oIDzRy
WpeotNT9wrBxKtrTLg3Ilpw/oYahtm7R+aEA+BSLvGjRRpdw+NpXQq8QJRNMOf+gsYOAzTQA15jo
QOaXCsmiMgm4b5AWCXG+HXoJoNkAwAggNnXvxtqHaM/aeOKuWCD5YiS2pd+IQ6h/E5rzYeRRObNJ
uw2jXAHtuwRt9HXWk3ZzZxD1iffbLAG9RPt8S7Ds9p4rIm/dw4sJo837EM4oDvbYeGhkM/qIxTg/
kueHgvc/20ZJmLF6M9nQA9bd14ma9W+eYT+BskwXrDJnomYU0mf6BDcjTCxgFexEDOtZi41yfN2Y
eeIm41PutuMwrkNzppj8slVQNFb/l3+HR6llOfsV5mGbyb9QwcGJoukPnPBEsO26kT2WlwVBE2eY
iml8Seq9u3TPdS3hxLfZ19y3TIkfQF+BGJNhnDyAO1eojKWGZtSU2NBZzwxUDn/C+vNVQpWRZXdb
fLiDXKFzkYSe2AZyayXlDH0KMY6pJ55VmyAvMpSsefCToinPH3lxWkYo80Qy9cdmtwpXtUsBS106
BbY0A8M4plgBoNVFytHHec33Iso4rnXXWa4Crms2t3NCZrmOie4x2CfmgW87H9xoT8FlwDZo2bGt
smU0MM7q8ns8dkZs/H5DC+onrBgCjgKr7irBDfIh3s/ESHIzIso9kxQS29ymPwmDXCqHFaYkL6Qr
1LJetk5p7H6fFIK4wTVizAgeA9HEHKJG+Dor+3qLpFgpkVSF9fWm8jnXK8sJ3x7I4mRBM5zFmLsw
Zap8GdeeAyssVYY/AVnuLE0HKruBCTqWk1YjuL9TOQxogow3HW1WzXwGmhez2t1ulHRcei0nulby
gBCBtuc38F3j+WnozjY+Ry3/68wiyqpcu9kzWb6yjjUzd2H0ZYZR93Ju4wXrGMzo4PGL8YUKmmR+
YEZHx8o0M9AygoMidvLAqrbLF/y3OSTVG4DwBm5N6MkkjZ4cskcvnDzQX39WUAenOIdIOVCkyElM
PvXi2+dOTNwHMLRnMG1k4NPkDgRZtBCbgLnvt8X90rwiaxQ6u09BuVKtdKhwAwyveNy4Sij3mjqj
xgYYynkZfMs8y4P6R2q4NYGaXoA0RFQicOV+Nq29g7tgxM6D44Ug3aSsB0paVNl+QiroxkxPg8/8
GVBzbMSh6lkyGMO6BUhAzvpldyYvZZXxbJbIVTaZ9OjhIri5RiPzpDbpCWJD6uGlHwoqFFce5pNi
i8yeyPk0J31EFAcGjs5QGYwodFx7q3WJukZI8VUKH/p+oXLEjfwwdQncq+ALLdBhbhwvE1MH2YL4
sw/JnBWoZYXL170KG1Ty3Y88XHM6AntuoReASbYaqCNV5y4FrvWJGpNJUIG2Lmvtdap6uEN+/e6R
LniV79imeKLJiodTFZnqYAtpoi6uKWgnQ7X0XETyyQIkZ9fqz6xAh8ZtkYvxuQjMo/fTJWMLQcCO
LRdPOyV29Y52rxQB8qRS3AAW4Z6F2XtFMwEf8p0yxTWhSf7FFxK5zp+S5wJimQLf9oS/acp8IvZ5
0fB2NZK0921dkDp/sfEUQWIRH7r/b+Z9T2rSFrobchJrvfJmziMAvMmbaA8Kxaqmt96GHBX57XdY
Sh3muGbeRwCuCNSYAJvH24qP/OCrCj20jMJxAgBkWqcu/K07GRY3N9p/GzmEc6tfCcvApcGBqg+x
rUilwM7/MMhdchF3k5xPdvD8+6DJW6Z83sIxTBOj+x6eV/DU3pxn9kyvPuiTq56r1rl8CdmUy9MX
pIYPFPkpaiVn3xOOY+gZGU5M829YONfiExFPkdm3a583PJ4m88Z5e3q0l0hpW3Vn2ChoQBRBhaTP
wUaXU/DAOlqmnB57diJ0Nak7YcTZ1WtEjaODTy6Mqw0fUwSj80bigihv0wso+v7LAC3lHRvTYLck
Zua3J6ScHGS7toDqHkGBOlIiy3DuHiQJRQNane8lpZU/SBrz+KLaOcZLVmFNqFLyKg9Y5c0TinJb
dd6wP7DaJlx/nW7lvQ1diaW/tj9GMMdX2qCm2cn43w193JxZpHSwIBtPPwAY2pasHVn12NAlLArk
xWv8PDjj+0upm9AhWUe4xRiM+SbgY9+fQgQbIAUbsLjRqVF6suSQgWKZP5ej9ZMNWVy2kzSt1mu7
kHMYT6CwFKZEc6ceQ5AwN5rhg2DaEkn8mEeNjsvZqbJb7EIejXQf1q/usBGRU8sVOdPoM3ZBd84z
zUIiI8pWZk10gvOHkOysc3dgk8K/gvqG8iII8jkMWR8Q8+VyLlCGgXCRWnpa1GqTqvNIb5s0tmmD
HWTL/WmLSRSpkUY/jmEa9ogT8KcHoZ2riOXIeUU/zoNqrl+wzeFv64EDE7qINIIey7DQjEp4NcVa
J0ZxarEhBoF03h/U/+9LoDD+VSo2hHr5YDz/fE1tkYmEMOpJXRYTi0UYOE9NqKaRNp1uynAw/+7k
toQVN9yLingsr35JoYVamEn6WkdGZQXo1dy1AJ5Pane4P2LpK8ZuF1o1qtOnnKNfzKvLF5v9kR/0
inkwZOXA3uLTDryOnxS7g2QxdcXLSJGpRWWb8PhnRM7OIFjaH4KEET9ziHeZ6+DqwN0d2j3IdCkP
eNxOqcfRlJN3+5k0kDkwxkEEtWP4u9W1tV/4tKnoNOo2WmLpWMKLohfoL4H6Ak2fLZLJybLh/Hz5
DYHSjJLlw18ps2IIvb5OlHzezTap3v05bWNdRxogIW2FXc6O3gPnPz4ASPx/vMzp5rmgT7mnsxBi
KSK8IXWfQA5MLYrGf94dEP+CgwTL+4j5H9saDjInCHK/neqHWkGqEq9CHmgTxkmNpBhvM6JULqb6
zd50SvaG8+ahQ6FxA/bkYAOxvomgDSMVH2zDsnN2pAIM7OF/FLjk1/lVRFnjfDXnN419ZDtY3oDO
S/BRn2yVhSLUWHWHjlSda614Q2HUkYesTSar3QdeytYWqPHqHBEGS+wO74cGGNRR9Wj+W39RVRPS
T4njUoMJViyQ7xP/0zBDUvnvBGQrp2YDeJIxFWvo68/tS+9JD2vh6lBTUEPh4KJuTEoA+q5MxZGj
TWYRHZwvJH2czTxzQ6ibCvRQvMOtRBCFSBOMl9Y1332WDbaeRQRHkZGvmoNEPag4ZJDDEtIpoXuW
PTshW+bu/I37gj7jakB9U67YC+nf1MsPFzHp8S3LuUvWWJqvKIvuDqqjz7cn5kv6k7UY8rYma4/Z
ygDhQDm3SjDO5Wrdgb3Wot1lRkptSVBTSxMfcs2hjc9/yYNo+7jTMVJLQcl34wr8ekfAjE10ddm/
5cgLBmCf52Vq2RVpJEO0oy/pWxU33UCYh6a6KwpX5mfDBXjJ+xaQlGs7gXQhZrRDGqznebwiPxnB
Gx1jmFIJqe+9l5CL5knZSh9M4s9J/Wjh0J8y6sSoF0yCmJgb4G/lF5bDAnN+h6GaaRDntEZnirWt
kP34nU1UjWuib9Q4LuNLbEDTUP5rZeoNZEplr1ZiqD8hFoG7yow7bcf88jKoLItvoGmUnk0WM7kX
3ZJqX/qk7cgMWTZpmcrXfnWMoXUD4JK3QDhyZ//Vg+sO0KsPel6pc/V7v8rJOuH/rtd2qULZ03bq
kRZeiXQx7nB2FFlxABOeCaksRBsu4R4sZ1vnAIChjuGAixMTIQjq088q2GUzO4NYEgAD5apryIRw
MvFyWVX3pKbpZ81ZgPHI0ZsOKy13yFiF656ssEyKg7tJ+eKcTNCxl84yHY8LOKeNl5zXHKIr8H35
+bJsmbX9rVow9gPl/9rmv+tS0/9CmbMte3+Isb7RzSZ1ZsnwAyk8YrPZjr5rkgoAmLjPxhkqEySK
9JZOI0VieQg2tpq2L4V7aDy537Sn9e08WF2kXtMQWZV9w2JakX+jpUw8RgqTtlr8C5mQhNqly7gC
prAlJOjeeVIjSWz5Vf4MEaNg6rV8qJm9nvihv3mIqen/7O+dUjDsjf5rqQiw5IYrDXpWRFXftXG5
btt5KhQfAEHYHo1JAUxH/WxsN8fxvIBUumkf4+AsXaVEUBwXKb9Joh2+glgeYOzyQoOh4hxi97zv
PreFvGDy3FLtOJQ1kkH5OudLdwCbdtpngAdeSPMD9uU02y9wyvvwnOUsQu3ZDMl6MsZyjlswCpZV
GWqZGM86CC6+0NLJSaIA8sNZbBdMx/9wmUDiNpz4kWHxQLMwP5yqdrxep3nTRDZQnUmncjVd12HE
P1I5SmXERIjFCo+V6jkNvqaLW7KFKXoXsByv5pCDUw95v2rHfy0A0d32l0IK/e1vXb4Mb60Gsfqf
osKS8fQDDFbhZfe3D9qpLIRYpv2FIYrjMfcr5MFtDKpGGHxyroMIjB21funzb1WemeVZYd+bAhPf
WvJh5HF0fjudAX9Qf05IEYb3tM16Pg9bN19t+wxpeauJg4LSjhXl/0nLecxKVxrmAUrKRtpgbpi7
etbEqlTK7ZQZ7oAfRVtiHmTfTq4YE7WRSFD5j42DwIyxerRmG/dCkkSS4NJPnGLyCCY8B9NC5cLn
IUVWf0ex7yuhwW5SCFzj+YPn82EPSA4PHKweZdKfb7EqBdu4UgkbkpYoc7uvYKExtdLPHjoP4L8u
uqVp3A1H+ilL/5V2ZsHJryuz40HxX9yTJbiZIqiv153fsRiUggEbj1ZtEilVQ1Z6ulJKIrAoYRCi
06jJnq2S4tH4EbrU0q3cwlvXpU+kXVie6fldYmYFjKuGg3bA0dV/zbCJ9c174NOfjLqf38JrKtTA
LR68usQvB+Yos1feKAU88wZp79RWJONX+mk0/0ZfFK3AHKvEoJMkLqxhKK8sGEtsnAeR+tLsxadQ
+2xUPZda8KJ5SaTYLgedr/5G2SZNxRc1Xgg7IXbxeIAGVlTdlC7kBSUbG89xrB9FFwxamvHPzcLa
egT14Go/zW8EASGShbLIJLjSYNasgy+CCRkOXxmIRzVInnAFukcrpCF9MCqA03zVp0N7XzIcHmb3
hT0xukYxI2oTI/Pfhu0QTxx/yVApNHdMkAXHhnJKOVXfOpSCckF765TQ5Cjb4+NAl5fa2RE2yLOF
RuTCSbw9mso18lUmmvofjvaSFq6lad70O6zBFwjyjT8VZaXZEEF9Fq4GVPWlowSH9qd21kAWtiaX
ZmQ7pFH89t7ucGnQwEW7WcnjqJs0LvP72C2iSeDnIX6m3uyJsOi7cg602KaD7ZqCtjReiV50YzwM
6dqZmc+Gw0W0UMk0kzza0VoYncOFJodtMy3pHAy7vaKQpO1sesZ5PStsuk4pje1tN/E677RuxomH
iePpr229Uuc19q6MdlpGOkhfcPavi7VN/3b1yxPeQVHfqnI5Rq28wXPfVX5FnsNwDXumZ96S1zH7
F/s6Ckoz3xwFaIYOnMVDOY3CuYZKSK0iHV1xPalHIcUagx0qjzqKkxpM53qHyLzxT2fLQNSSYZAg
iNqtsligUnI8H38v58pcTZH1h+nz3b7Wmsi1zojwfm7e6EE4L5zcdr/zy2Hlvg8TQGhGEKvFVgb0
6OdlDCafLdHVShGw2qQH//ZNsXrRthsotyGtOPgYDSYt76q+AGb4XS6kQyKRI+fnwMlEjwDGh/sZ
b+L7OVmotbwLlYbzwQkum9J3KuN6bLwwHgknOsOWbiV8auSqSwSe734N4AqGrnHPkZ2kjmTrszAv
he95d821+lfhEvLMsCoVsKIr5YrTo73gXS5d7AtbE3SFQFRhpCJnOdH4Zzet0ssZkA8v9uKp483u
6EHXlhXmUI4lv3XwVls+fTamlTHNvVzsNH4RWjs+5hZ9wS5hzGK+XYmJahe9JM9vndkeQ0RWnRXy
UxJohvveCP9OHcpMg3Em4FVSg3YoOkT1zW1m2NqnrY6XRkK6yVFKSFDQu9YJkVHKheTH67+g2VD+
bQ4ncw5X9iIc1ys5lgpp9/5Z/PqbqTkTz1KZyBa8Ubdo142SPrL2ejen06p0zzLtktiQ0zkqc7VA
2pDEqePR49X4PXordab5oU5/07PCunkjJK1NEy/1aXswv6db5nToAS1My1dFbrEByI8xLv4S+Rgn
IELO8DT/QYiwCMq9chQQ2fQ0fi51k92o8/K9giG0gjbv0JaztMnFOb4DQB+TavDiQUSiZbnhOlWr
88E3ISRtWme37cvCFKxs4E0vRLhq2YSB0ysR21Uo5LbJ1Ghg3kBO/pu0Y5GyyhOFaQAxYawlLY1G
pGbKtcm3tVO0eWTo9DT2VYwJLiQxtoRo4HUjdcRo55pKKVlMMlWP3SRTvpLhUphr7otS03Tg7U4j
uPAc2VmlT/5v5+pICtip+NQt8JVukkfwAonlTEwm4vJGc5g5ecg0tdUrIp1+Xyxqmay0GZoKzqvP
zd3HgAsfcfMd7cQKHQ0BMTgycpGTY75vvm2nOQ42fCjGriOJSohfNzh2uvsPTNWJ1dcFrLD0vSsN
37saEFEQ+0csyNIGRlEsfzhOheYLdPZWbTzhsOtYPyH5HbB6oOsNqM+l7Ky8ubc74nrb32BnWolZ
rgCouZcJu8OTBTk1UUc+SmkTaoci9DNd4AdGjTNBW71cH9ZEHK8x2EeMApgcMpD10qlxtkUAyDNc
N0BNIMm937t5d4UHmZT+BRM3VrEVdDel9KcrS5++glU1ZpWvunX2g23fIGuneRAKCjDpTYZxtQge
6H46hcgqXpzniXoRbmjY32tw/rZl4XVkCuOA00aHMob5u8YqXuJN1rurEka0mipXBP+N0Pno5hob
02l2d9i8dn6wKnifUc2F/PMYRQC8wLJZkSdZfnHGz4M3IK3rfqH4cRxNT//ANo7byJOGsxmFFSG0
NZip3gwc2X6OK8jAGngDpTJohzRbTvtoFp5HQzLXxtuFxHR3Insheu2kY7giN2Fhyh9QVgiSodBw
ZVbhAlwGw16pfKAPZMfppOtK1qZrEtWckzr7xnzTRseFwO8PLNUtuCDz5aK3hD0CyCz5ZvH8ceoC
TQyHad7E8lGubmbAZ7+MzORrsqGGUVnWd3QQDi5wS1diG/8eXR4VGgN+IPo3QaLH6oKx93Pk8Xgq
3SX/nk+9AMbJoayE2YPHshcHXcwJoGpwvQneNvP3WwMK4MlR9TtoQhj9/EJw6fDzhkTXVteT3kwG
LXWSvZZOrHVFJygKVLvCx8WPUqbasSP2daqB5JJVarN2kerhUPIrdD+rNaDqXkMy98PAnhb/0RTI
V3Onow8OGB8bRSDZ+H8ULCSWVzwA5WnZu2M5th4MlSLIQ747na86U95NtDKCu7XNnMGxwFqmy5hQ
YsilmmSb3srSMN84oi8Nr50J7cWl+FZbeGsfnceLNNknl2lqMweOvDO+wFXSWer3PGQNF6VPeSDe
bA9YxA1aUcQepZjvsj1qieHw7wT2021sVV72YuVyytxKs8AreVbqYq9x+uDA6F6flFHW7Yp0e/6P
rBq4Fb9PQ1QozOqSPZGbNhDICaifcis5KAg3Uwp+krjw6BiNWrRfnodeWWvynTwLxrRZy1e3rWd4
iK6qswIAhMTCUmHoMKtS8Ur+NIw7Pla1mHI5HwzlG2RJTnd27fvvWgJQLZ6Jza5D8dk/w18ZqePc
XDdfK4DjOc0Wu6XNUlFbwibcXPoKAFO2hataKdFmu8V/WH/5zkNndZnF9DIZKp26vTlCfAPfP6Sn
m1vGfTQ7cDPB1fZfzdX47rVSsNaCqsF2dSKeFc8A28DOzYd0SMQs8EFtsGLyfIlGnwINJ1x1FbQf
qL8AVnLKRXCu7hpsMKmRCtifYVkD/OfOnc23iYyjMYQhsGyK5ifJ7kbHTxZH/hDaJQSg81Ycuve1
egwGeZFF+3A52TJOsuqvXq2pdGduicAeqsKFxmGRzSHODHhcL6BkGyoOdY2iu0esrPG13hJMWHtY
CfmqkR7PQheKHHzw2xXI5ylZ6C2q39T7LiSFL8Lh5YOssz+bcFmq1RZSTgGaho6UF2UxdC82IUqy
k5Gp/O3s4kUW5OSdkASOoWKHmLFNdg/MOLjjTQLyS+xEGXkVmKQTUnmrZ7F4uduyilrLSCbmpWHN
8vaWR9u2Ft5pOqs3P+Vg36l66yEqm9h9Vb0hpM8c2UwGFzrC12hHRGC+VuJ74wkFlGMuQOIIp59h
Lvloa/BnxdoHsIyep0nGuPiavlT4oqbhl+670mUYS6pXmDHp6Hdfm/TNCWCz7GkkAOWKmRBIAMrs
+8YoOdtNbZZ9JoVbht/6daOWT6cNxgIAlOynwWpENOKHVIf7EIF4iZoCCo8vl+oBUuRCdUfh9yct
Fy3VmQFBDTY4ZX/h8RSxsLTJPFjLCOyXrVaOeR/yWCKGt+eAV+tEaULjqaw8w/lOuy8y5/ayUn69
KiWogU6jRU6OsgxeCsMm6x1+LnnC893AFbtU404aqrM4D7Zv85H6IRYii+jIIGgqyEZzCBKxGaZI
gXb1blvRLjMY1vpL+P1sIxCHcK/x3j+ngeEtoUPW56wqYvRoc5KFibpl1BFD7g3RyrKpc5SIBy5B
gvzoxGd4k+D1hWoEjtdIkvWo7eXee+6obxZ0rHQztuv13kAy0tZ+1KjPIT7usOpCWrgPP5vVf9uF
anIpT68CxARc7FTOj2kng9arj7eCMikkTpG6v5OirmUNXb3+KWwJ0A3lzh7sXMSy56znSpkroyBa
qPdRLkp2GKnix07pLxEfnoLRhQgSrfwb0DWdYOUWLoTBzuk1g1YbS6SROvzUiJ6kKQEOnkyUHo0I
D4NUPzDW0NQgYxAWsXx3H5SiJvtlPQdOVEoUJAty1B3zqUsBjcgVF6j2p1rzrrxJYYQpd1C86HOR
7y56h5Fm5X289FEfIfqjuED5jm1VVkIVT6afaZcPnH+azkSj9RPHT8sbpV8Xbp2FwlNkp0CqPaMS
JTsAnYJPkvMh/c8rQjrk4Hppm76leJD+q5AuQpvB3Y8Mr+wiaUd9vuehaydKzVXnUTFs+FS9OiS2
KEVsFd8+grhmEtw4F9F7ycOufs1nq7vWKJ1S2vKKxvpQPNQS4m/syZ60PaidvzcxwcdJaBD3xFIh
vr1mWgRlRnteM+/WIpO+dFVJsiKHaLQSP6G08yu+JtSCR6Gj8sZxR0AyF8vmR1JsS6S8fUA9+crU
3Jkg4xF9Rz3UAYwiIlBVG8wQpw0Quo+urzqzRf2dfrIFjvTppB0+2sgdWQtKTeJaqVikhT5YIxAR
3Nh42swzz6SWSC4ALSZOaKrJWBzWhUf7CVd+AKLqoeMasrcbxhd8pODLgLkFIKA+s7joN3RqXhsf
AMB6xQtESeidOIZ0++GBXGKjMgR+kFg2UIjjJD7jmKpKQ6QR4elqJqmXUkg5c+lPA3vdZWZXekF6
9u1N4B5OKZnnUzxu5tr206GHZHYgldUvzWX149E0W+tK13Z4hwd20Ja1Hehzl0520RX/TkxkrjsJ
CvJSQGeEE8IjH3x0+EC1UdMdcicJMydbW9yHFI9p/7/6tZSmpARn0Z+dgxFg5TFaN6dv2TNNFwyN
SPup2EWN9JQT2ufU8gVaNsZHisWSplOUpoEb2GANqy6YimCNjnvHqPYWCCZHU2w+SpjSZ+e9Ilji
LxqswQM9omQTJUD5NkvRRVp0YZ5MQmaaOeI/xJez4A7n5lXR8myMYS31Y3zFwYns7tjH6Op4t0mf
BII+f2gKrf4kPC08raPIwSKCjepXRovQ+gTVP6LrPrOmKFuqdlLygNbJtSLZqYHEiLWc7VTTcjG1
G7Hi/iczzO7gypXATeYOD41GdmMgzw6IiydiOhvZ5TjqAYMmfLzrGU14uw4QU17HXRzXM9SQ7GBA
DnmOJEtWrbxGZ3jVdBPnoBM6HOroBq+Tr+Fy1skeEBD3GyvF//x6zJYUb+kaenYag7sEx2uiB0TD
Gagsr1I4am0ikMTCgUGfntYqFmFXoxUsFQsF9l25/f6BIh5FnCu8b2nExaCkB/WyofO/oQ1mLKg7
4uIaCRMUyFF3SN+5CNeJlWUt0nafvKTl9UfPGvryipYD3LAtZwb9/ODljLY4fRy3jJvBabW098Jl
4cFgTnTP60lMccbnYHO2nWzqYSjeD2Mkwt9nThxmksuhYgm0mGU8fkXfnAcwtj46WjPo/Vj6xt/+
Ufb005ayqedGgbhxKtdHUJ41DMNu+1qhCY6Oory55VWpMJwBDGoy2mPGMe5RMk4MDNx6+pzyx4t5
qsq9Ti9N0AnQYzXYzTdhtd2OW3Y6g5zCQcTjfQAqcvGjm+8ALPLRdAX8Fy/znvnArYSL6APNEfdZ
5hWEFVahYZeY4dp17sylK5aGoWQQsA2/VgQj2mD2N59Luoxc9k5gfMuHj6QCdOU8lBmh5nvcmFwA
9t7wWb0ICMgfAszhK0FQJb3eA5SXSJQplOlz4RcJHEQB3bjIeXa5O7vTcDVZtDWrY9U3sAdHinLu
GIuH9OJASl0mqfdsdl6BQYrLbYPRLRyKwg7jE1UG0cERGwfZCDMWCnvheETnaZgjvArgQnFBtsqQ
Oavfooqj8ECZKJkxa28B1Rp9QnIdCHFoyd0MFI9yVOIrq+iyV7X/oAzGrYoR5Tun6y3Nhuuheka1
YNaL0rg2qdqbSZSDvC8RZofhmzZjtzGwNkb0VRz03r7jvp0jerbvAmtffI93WCWugolLZ8Xboumf
z1sSXkkVoBrm6Kg23AtMfKIEfSVhn/5xzeZPJhY0pd5S9xuVqd4ndW7VtatLsREPHX/vJw6TwlzQ
si/IabSXGwDXgMZcjeSq2OU1N+IWz/pvKHoMas+TiKgjwB2QJY/7vbKI0qpOLDJArM938TwqzzSm
OhfsHMR3EH7H79K7FFGpFplPZigO9SrGY7AKIPEIdBLT/7bbfk80SrgC6XukqWh9npUEFXZOi3HW
DpjkIhHoSqQZVe4NqOvac0RGHWGDyvytyHlx5yBXiwmP0oz7g9pRM7S6/5dICvNXOHdBlJUwaRyA
2fc9fc55UODc/Mr1wQt6q9k7EE9q3M2AbC5X5tMenonScJ2R1Xsw2FcKwGJ6mkD2BLMZVWiPbus2
FA20+RdLPva8slMvW8VkVnbw1zNsETpY9JMuQWdutpdBCMxT7YlqYrwKskoQxD/BO72uz3CL/xdz
Tics0oXyCQdO/is70MOB2JHh4AzoyC9Ss4Rku3plRQn0zi6qkltHi1dVnaYIOStV/xc5eYiSEgKm
9e/P34NzoTviI60p7rCQWS5hS/CA4LCYkf53gaN6/i7TVAUccsvBrXgzRPWnmTsrC/9FIfK6pZOE
6mLTHl1xmM8Tv4H/6aw/3+4I33Kd5eQwnFnufhTD3/Xc1A9ZYzn+86AuJ5hTSq2PdZ49Vz1uHthg
NVvuEDZegcKwJShOZs7M7PxEoHVuVlq/T8Qmp3V9k0Ob99YMDJRix7+jaBSjV3ez9c3+w/vAsotu
7UDvFAljzI2Ahx5L9aCqgf3BMvBTMfyqBEqI8+F0hHTR/0GDkmAdwjgOXo4OzgL4malYlqSU3trV
oCpmB+R5jI6arMELFYkylCEuyktDlMpxB3nOYJeryAobNSIBKFMEgxpcj/gU3cSios7FWKS1xpnc
yXvtBgPOvtcF9kUsro99Yc7rLJKjVVJKoKTK3crJjECcXFyXFoWRDk7eKNzRur3gUtNulSq4lpx5
uskDgiAtKUISV2QJA91IiO9e0EP4WCuXoECoYg+y5Rcv/jIfAlNNrXUWGYWW2qrlGDKTI/MZK0Wx
VF/jAFZFMN2G3Qi4sdkYqRITpJjJ2eGKSgGmrKzI9a4SuMbmd/eFW0OeatK4U1uWy7fAc5i8imdB
A1ZBfohemVQe6fYyVhOEjOlTRztSeXjd/v2i0Y+tRpfeoAvtiW77JCRc8rwmN4eezL1vXRlrDBwe
4dwpp33kLsuUWiWz075AZzURATvZqO40RcBo/pJdCu+dilIYJUj98RCiIfH5+4qXLysqRwYyFKl7
H6Kn6uUZqzXY1PRVDqs3dtLOm4a+c9Jx+MBFAVFzk3r1B7dwBweVG9FG5DclLsSbkpSK1wnymJnj
tfXIhqe9b7SvqeWwb2rYDB+++ROhUpHunRHVkT2LD5oJbBJClYD1rQ3himf1zqof+9KMEXs6lsJW
qEnMdPm4wEZGqCgf6U8fUFoL8chIiSGIFdbQYzaQzZK0UvQKsWyU6AapTFn1o30VchuUSK5Fvbfs
qZ3J37BoaxhvB6UyOxzfi3APBBEgJ/upMscmfCsfV2kzqk5Z7hu8YRBZtVVnmggzWnpM5wT+QexW
xZjKOGpDH3VEp1swvY6wlHh0e1z3iu1rPgqLJMEKFJIy2nlyuuuiNMk91bbu/CStVHIrof4tsdxJ
102bBjp4KcA9MVq2/1HeWJGgG1yQxMXepHNva6UpfIAW6d40bDcuCUD3byqZy8KE2HYYOWEK2aIA
jZy4FeJ4QqEX2HyuK1rLJI4PgWHE6VG6+v5KtKE/y4y6xyl4eg/SmYofux4ROzFzlxNnhPU+/Z2u
ADzcdAyVSpBEbd+zZ/2/oEkDrrqsvr3Sv3PjlrDVf7JZU0CgxIEKASwXa4oL3uYKs3AG1Kj/w6fm
BzESibQOJ+HmkMIqat7A3UiqatWKTMilrBOvMxZQNRo/Fzq0qbyNbqk7mEfky3CKNWwR0ZsWW//K
u3U+8a81faHjVuEc61D3J7eSaOeDTkqSoNaeO926wjNj7Z5cydZ6zhysKzm8SSrCG37h2uci1EYm
7jNX8D6Bazcy5zVc3U58BhZZzcqIkntiJJ6DwPbUVo9jGU+Qy06UrAWBsOhoxJujc17sL/bCXmtL
fysnKOkkGPBBpV5mBAaVAEh615g3HT2/BHJScGdxujh/3xAomY4CcRyf3VHXrjeyZbKownv3ejRP
N3nMA69v98jiJ70oVpzgAhDmvIXAuzR/Vf5ww8aWKjIo7yvUlxEpP1gRabvQxKipUd0vOXDNMjgU
w2kSaF323HOadLrnLKfXX2yDHnFUHwYt49s+/JMam9FjQexFXhnWG+8oUYvhg7sYmwfQ2XllK613
tkhAgfgDlC2SUShrmMiwbYSf29AsR5FsGu+MzzDhwzW7QwGJWAg76AOwFxnA2C15DidfwXqlP+6s
nHblLPDeFDK5eufDH+ScFllI5Ey5pGbDIVnaXU3STG+HF9MO5D+hB0tLg6tqb7iVePdahpSv4Kys
uIN6TOqvJSMU4S61Dg4ya7AZc+IVShpofUTqXLAx/bv+SJHlmSSRiGNkSlki/++7OfeAR+/lxSln
cG4qLaWhyQliXYDWW1uWXqJcnEIZeK/zqZflU7LDZ0vlAu8/STlCvUk2PBammUtbBWlYnT27QHdT
CxZHVTP+UodYxiNN7VJ4tq3lSZsdAHSez0y1IicL0XwmXl6ITILAhqvrPNPc76eF7RxMydv0Gj1w
Ogbt4kVievLdUzJlFIvPrCGB8UJYiBMsJUCkc+aHYIsdqnA3+MnGHiUGpla+qMrJScLwb2t+i8wQ
9yy+N1feSQ/S8nMjZ87iL8kQRPSm0tlCUblxZiaPS3mnGzP0BTke44EInigW2zFKFcrREaYgTVwC
3safbq5oFtjf1cRKyl1gz98M1NJngu+n+LakKhTq/OoM66bm+9yeQjACYSbg2f2yyWUZF/gVKt9x
A7tpNL9ur0i3Kclh2TGZJOgdQKGdsAOeDuRwv+Mowogqyu1ebOK2BGWeDG8d+tbr7UPHv8C3jY0K
DTBbfwMOyrdn+XDQllUruqv+xTqnm2+DeiA/VjQiIKNYJu139J2cb3NXnkhx9IqgFAOsBhxnjFXm
fmXKB/Y4wzjRPrPk7IGsNAWHHIYQKAw+cowXuucMIFr2pfzRwKb/fK48vCGVmWFln2aeTYRALxiK
/3rmukZCT6PKrpE3IhTIpbecolPVBzxPgD5VRNoq1i5zBiUGAPC0B7oGADF+8FgsxptIDE4fWCBv
0XPoDFzJaCYEgtqBvTjx9xhVSJ4Vs0M6lyx8/SBLgEz712q6NLpnhsWe9lQqS78o1coAAX1HECEj
Xxg54Fpo61Tr8CoFYTZD69iBtOozQxXiEhQVossIfXkw4NOlef39uHv7Y4HZ5jG/PlkixsSTIfIg
5hms/Nc/uUxy9mOyLUBOd4VSBOqFu/iYNS3NgEw9Zn475mcIlQBOdqLLbYSmpy623y/nZYmGWB6w
2LbBGWcEt0aJHZFqVieDYpBWrx2bBfv6kFo9sr3eehYO4IoIhlPz3lQmV4zJS5/wgXZEQrRYPVhy
SQH8Z21dMnMd4NLBy1gZYYV2e9dixNB6lOjUHlJ+q/0Ot1FlEAOjR/QDUdPJh3XbHuezVDnOstv5
zyX2vib56cd+f1YmYtdZ6bCP0lb1XnjPgZncTplzhOFQD06647ZPQjlpdCfATYbUuwLFFC6Kzg5s
iWBrdUGIcK8cSdhE1l7rl5tASUiJNrc3QGVmi/rCMkpnUzPfxC7OFLnE+8YjtxdzlSbARi30IEF5
ujbaccRj5yVHEivA8mAE4Zjla8Kdv1RwM1u1LLcnBNxuoUs0Gom4hx41vztHCOiDEqVZkGJbZKtD
7/ex9L1A8ur0PSoaLVA86FMl7LAyRZyv1IChaksb2mDrkuM3eIJVl0gCyfkJa3ZHkSjVFaxj8w2c
41yp+Mal9BLLJrh7BbCwmENoI2lJ/8rzzGeS43wBnbXGQjZB4RGTS+adWlnrnqJLvTx6nh5hMjx9
GOFmUiCxPtUqpEYAgcs3UjuV060B4l/dLfAD5c46w/BXgVb5VK9h3LRROWfGwSyEa0gXhoKwfmnl
jfxaKrQZroMTikwTc8E2ucT4EVtpze9IV1isrlC65gSwMeP3xTSJQO2o2nSv/1zTe4MsMKKeIHaf
dyy/1nXj2HzJMSsW9GU/CHRzX7eYRDeAA7pM1/aX8W5Ojx2dW05dE77lSiXJXtMnGfA4fq9o0zrE
Im/oWsGophegE//IhqSQqg2Ttx7/9dvjXhraR0VbrDbd4teKKQiD8O3NYbQ7bplM8y/7CvmJwJh+
WFJKFvG/4rgYrX8zIZgYplnC4LviCJjwLeN1gEvVDlfN2kQIzmnnCCri/l69ePrsd/kxAY3z2Bu3
QA1AJZrR4ZXm53AP4GI5X5NqQh9+qxZlGnWNlHndhPP4jpTmnZoJI0YqEiagaI1mLRyBwf3me1nv
W9z76Uazs9aHeFtR93VTv3Eh5Wwyn0NqZBFo0vwkoLgq+1hngnmWopB2qOrO8nflF2zPHZ8+yKuo
tjIVye339+A5q2O7J48d2+pdEVId5YqGluPMkVtfgNBFoAPXCUiPa2eslBFQ3FDGXr/IVMby6SXu
d/7KLRXRG9Bk4lh+jj7HieGBkf9eLl1m53x83bqi7vYILsKeA0mbD+fnSAHKX12uD+ckRMXfDsiV
QJiR3SqwpctHB8D75/Noxai+U0nIislIOIjd4O1Ork90E8nDBHtgPM+f5pb5LliBnriL1I0woBGN
qMFrezcFypbv5ATVRRA2OC9f9ZWfv7XESScjKW7vyGlsRIYzFeUDHwdCkCw4WKvfssNhXHFgDfnG
4JSteLaelkXlMBnCRBLBoD0R5VHD2kCALyNNeTne3Vr9nN5RvjwQ61kyjaGAQIHqh391U5x1Ov0Q
fdwoKlkVeQwyi7eN3yq0RadKK4QfJ4vFdTeTi6ex3u3RNntk/H60bwlcQ8Nsa3Mqgq2PFq75MUEW
/kGK7JEiNdSYfaWtBwwxcFAH3ekWikMcHODWDZymuHBh6gy8cj9TXn8P6AS332Scj5/8j4k1ojD4
hhwaGPgTyXBz7dkMiYoH4S1X0Ee1vmP7B61pUD6jGy20SXozybUbtwnlfTNkCZy4DzTo/ObM82mG
YCaKmXUfqePwTDt9kfB1FtKtvVBG88fGHDRnznZOGkmRf0OK9v2u3oTuRRfSXEzYjfOsH2mSZmLH
pjzEQYcq+IofAnfB6TaEm3CEyfhkssjf5jt72BorpvjlJRJFRLeHUlxV447kvejuJfyOWBLcMgSV
HVlEkr9jqZIn4wi3lL6otlZPdPTrhFUu6g0rCbpilw5QPcm8CuSoS+iqDuRG3gms94OweIn51Bip
L3Cl8P4n5LFbl90XIqJ16kX0puS0RVF/nKOe1z/pz2LDtvBNfkh7PaCp9ycv9ZhxWAAgOtbuS4yc
thtX6uM1NymE9EY9piakJz0ZIMfPRhFUw0AGwvEnZ+RbYmyrXq0+LgSBFNR/wHPYN8HIMCOFk9g2
LtV7E2CBaBuZuC5syC/WnVIjdTxchDjE6/5qA2mAM9AcMV20ftg8YA7Frg18uYZHpLkhFQvLg4H3
R2fQhUS9DWWmtlX/VzYehZkYZzrOxTK/KLWameRoTLgptbiuueEkdMIBvfSO0cWwOr+tLbQjYkn0
gTH1ZN4qS1Gd0aOo3TgI5IN7T4T5QA+dpbTcDh0I33kHYkctCxgCYVsDkWFvEoCwl7Sq5wq4z1Bm
UUt3718jVEaZfBn5ZtuGyVHFgcD96LOpiJtL+NuevhddwCOuF9IbZvFsdcUErL6tB/o7aAqEqIrD
7qjntWGkJ0uaxkG5sDgCAPg2QgCxADGU4Frn8v8VV6sILKJC5ymNQ2L8wBei4/Zk7AlkxDZUTiCq
C4CVhNKSE924de5qgYu6ep8Et06gWSquuOwxHGCH3Ar4/c99PZQIm7iu1VYZDXvu+2dc+eldbo2U
Zz56Fk49JSPygcaW279FPGZ4QXNbgRtjbLRCl83aQ6MN35h/Gqb7Y0ObfBv9W7k0ZE1S1cwTQQvL
4x3t1lryXR0TUQkg4RGgayLDTTSNUFk2lFupvvBbYAvbDfra5t5ENF32hkD5Yi3M2pmKcoxojFX+
qvv3UpBlGs2N9I2HjrqFYeo8zXSU64vH2nyFIxxSPVBIm+n/CNkaS4zLdSiysAelZRlNaMgkPf3T
TITd5tO+Szh458CHSZ5oPo+z5MvdEhk78LBzBsmMVs+Unjhbj/PrwsSrl61US8otDnA/4RTgJE5R
cbtWvHY6R8dAr/0erIKfIvKPVyMwSRIv3yNh4jaSdgFXSX5d7pTo3pEvvrSMWvXE8lTV58HlsSEy
UwlXVH+KSFUwhbng5nYnlkcJULDZ+d6wvMmzPVdl8Z3ySlHYvzul35zyZJN/WYaNO0r9+MnVhhc2
JIzU+Oi1VMSQ/L9o/LQHP9hIP5ZFihvgf1BWoQiZiq0PAkPy9XXTcZVf12N35NbL7RnHyFUl/iPE
In6ODUT14QnD0q81iwX23mx1KR+JxyWZVSqBRwL/Bm3n8gjtStd38O0Rrqh9kjb1WykMbueQvsIL
XkaM11/uWtGOc8WJyN/355Ajb28jynFaH+zInHR+J5QdC6xL4dLEno92/bWnvbqnjY2XaB7kBq3i
VgBTIUMMcB+cwxnR6pUx32C7OBphPl+ktMB7Jgcak02NVYOer5+u7jOJkYYbSmPEzXDxw9BCsNjT
n0Lmxo2uquGpmBx192DqI4IZ3l4sBoJ6F38gopujSmvx2lVG62zHxM9o5i+fegjpSs72QTtOrwh9
mOeRmYPKvkEWffwkdvPUC5UCWNVG5tr11geWk5X3ldM0wS1YMdtq4DNr8w+1cSv6Y+PWvl/PLVVs
moZmYv0uTZg6bMOZVidciTRitHxhs43kxua3zdHveKNkrjfH6yVTa2KXd2XDptVpdLYa9EFpuKtX
ubjb0XXziMtSGL733iWpsiD1mgNmUauzgvFe0JQLmQZ/SpJ1GXJvHUVBeSVehhHwUWxZ1yT7vWu7
P/GKpyjmzrAQjIU4ajCig9oTRCwBLbeNNhR1+GodQUfXuOcBXOyUcZ87GKkrKepaxYrAbFdleSli
mr6taExtL2YzfjJn+rEEbRkT+jRQZX0ttiFN6aUI178Pnj3yHU4DjoQum2D2KCDcU+RvqtPn+Mob
iajZgX9itPI5Pt4g45h8A7U3zgFFU02tXL7L6YbaMYV9xyA3f0Oy4gMYLkg+zBkm04GFGfrFZYY+
b5D9KCZxYXrLGMYD8MMQmsrKd5di/4B4hyqATawFZDqW4LWedZS15GMbxQF0QN2PqJh46tbiq4Gm
GcvddOu7TlRRSCAStJS4L9oLKp3nBcJ/PS6fbGuRcIUJVTsKDMDJy5p37obvoA7uVmo+x71CcWG5
vF6zRXfFUE1BHQO8rFH4YTzlL3lEDLmKYUFoAAokl1vdF5xxks+EoUv91LuTXz+cx/fB7Cf8yzxB
ZjtWBR0TI0LI1XZ3f+a/OeNHsKqrIY7IhhjSVxKxEhTVxD3nPbRCrEbvNPYBB37DWX2w0iPFx9lg
FdqFIVc6j/NC+D2YP61O3GP97yLXxmd0qaaQ+dzzvzr0Nvxx/ppTGqao8Rc7kTT1m2wyd29xIIba
nIASQ+SX5bof4ruvKe8He9uaA+1Dm3hiZ3N696GNABBV7n/viJoC2J65cuye7boIGTWeThJRqpvy
1odJ8IZaPVQF5jMO5gq4SGyVh1n9lvr/nKFwUPs+XXZq/7RZ6nWNDIU8N0U4urEUGv8xBB+iUT0U
PTnznewtHz9x8ZsJYQ5EFc2fkYFY19YiX4fM/BMoMxIewHpne0+AWBPZu4tLg5S6ifPl2lu/CuR4
DABkvCBXRh/7Fp44TINw9WB4Kw+rMSlc7Uz0jU+VjY6TIWXfVfy6LcMP7s/IK4B+ZFYPRG1LcPDe
juv3dSusxIJnxEN0PeKIGmpE8lKJSWTuh2Chm0a5hWp27OWUNQstVQrPH8bM3wcSlxJ33KoaTpLF
P9juCyHP7+VEzw1uSyPj8G71A9zGUlWgPx9nO9IMTZaFCwoEEv2a16AiHX9uFcdI6FKnTMyuXwf0
+MBy7j/0o7tmcntGy/cpYOyQNR1pHYb5sZajXcGYtebwhQ3tuh/SBMXvzSYjshQZIONtwbwaC2ji
ZaiHC0Pt0xZwZ84+5WwWKPdJkhsTxvecMb2kESwwlyrGrWmhXRwyzAebK9nTdhNKugV8K/ojchEl
w6fnL5xMmQBiB5mzPZvJKrnIIaEVN9Zh3rgPeF1M/yvIyuex+X2qERk0wLM5qsBsIrn5nYI7LAU6
Z34aVh/NQ1SMen53siia4wMkMz3y2l28TNZjd6Fcz/Fsgp/YcRlu9eaGs5tLflLXVCPhI6Oo6cnJ
t21nnAIMR6gAjowDinPw0pQiophmelsUfJC3NvNTt7COLN5HkC5OUFKnL+42hgLjItjhzS+IFlZl
E9PqT4JEVxlgw2gNkhqmTdYrXZEIdr3ZeXczFxCLEaODFRMVLvQZ1EHJO6Fs+jCvY8RqPuKta/hB
pPdNwYvPiH+5AMWPLr77ZpxMfFqluJ0DIKKOBmsy+i3jIzqmmegXTYW8qhrmOGCLiDGksXI27bqP
xmXJDGy1Kc5U1IaiUbnnvd6RK18F/DTnKhXsI/1Q0MHV3Ozc3p4JjrVuNmRncFKrTORaYqMfzB3/
y+iOZdduT/goJQah4G45gCCxI3y1pkBBkhdxUEpaUNxGWQsxxh3rWrj3ng/eL27NG83YV7/a5Qdi
JKXruEDwwO6xgqxAU2ClRAyn24lAlgCwnn8E8hDQguHuz8dD0zMHtZ3xTUXLI6Tcye/Tt9YbaOPA
SYdNG+PeivzPMEwOq3GXEX6U9Z82ZDZRSNlD077ObEDTq1Jn1QbLOtgBv5/oPo/7EBTD6LnPmwNU
i+Eto9OGlkgR1xLpVjVnXgkwNekT3JS2/IUHaZiYCZLHwG4Knt8fN6OaTXxldGuzv0CtzjKZLIAm
aXhnaVNgkjyw+kTbqTcAd7FZSl3fuiZdJDIumHVedcSYypGT4EAX7kWx5j95HNvHGc5eDQC0uHdY
K4mP7vWIrRTECbKp3wfFskFmR0EOQf+CDRiWU1zgtMVidevfCIBgX6zErSrfPBKj3Gd01qqFsRrp
E1576czEUYT2bm/KV5B/DQ5n5J1sIJmQgth4wHPqeEyIUSeRFiXeof2QC2EW/2LEdkCQyuVfI6pu
Z+VfABvAwQsgaFgupQmvAacz6preNVpLP1sj0AtPmOxRdlTWt/en8A5n+lVSrYVJub4Ylvdjo7VB
bp1dC7DVlPinzzjztcAUKH1V5fwlNIRfQj9Pzv7HM3HK00+TednTcJlCrl7ZUeoh2E/r8LcUU7Ky
jfxM70Sv5amdE5zq1/nt3VIKrpGqzW2rA2FJn59RAA8bhTWXTPq2YELhX/J57/v356GKHDxqJMWT
l7rPNzIUW7BqwGVwyEnYS4nQHlACHAnMC0ooz0FUPK8jiP8jjEd1T3vXNt15OWX9bDDHihLCW3hZ
yAZFIroic+Gk22lNmOpq6EMyBSKfp5VkXHjE9dwuNTtUjq0ZgpJbXfoM6aT51Q7HHAUFSTBDHU53
tnNoNOKcniznWadxHWL24w1hU9thPljt76kOmFCXjcWeZq0A3xLZowx7LR2Tz4DdhjuVXDLiFMhr
o4Sko8gUt5G0aUVHWYqSbinYgtmLeOX9UeHRUUumWVSd/70L7Kl1zOVqUDvpgMjVh9w/4Fwc609c
AFxOBgT8cQJevKPvExL35iaVJrWP/dAHBrg5F7y0T/PD3uDMSeMZ2NmqGP0Irhs+hITi5ZZFAPdC
jtaWAmVOesu3EwSO/8nW4x1kv2n/CypRopeYXynlee5Vx0cqb5Sb/0nPY3LoaNR0aHu+pr5EH6lp
lM8bGp8OEo4W3wkzfZ9o+/NM/Ojaf1mj0muJ+hF2AOMdElZmxne26x9++GFveZwz934AQP9JLm6H
2xKKalzoy6RLEkpTJNjc2HCKJDU+uHb07dol6CjNeIW9puERkWyKCLAT0NHgfmgtNj1gYAfiJGB9
aPCp6OspibscUUmSxvZEx+m6cqzcKfjCqoRZ/0E4x2Es+Xi4Lw/fForo7Pbib/JV//Jsv1/6PR0a
xRg7sIw5vEydMS/amlwPNbiyIF08xmq1yYVnhXBs4WzOq7DWs2GZ2uFu3O6kyaH66h2yJfSVuMwI
QqVgM2DINQCJcEsSo6uyiUIwkGldTc9kEsCfpeMo5Jb2u81UVBQY22OmT/HRvtkB/afCPROWuVHM
Vlr79ZmaOFirjDHC5P0b/v5M82DRS1slP7oE5XE2+wwsg+mpS55yHFx47W6IzSVKlj50bbrIsw61
CXv3YZeYu7iESOze6bggYRi0JjG+gFkklWAJhg/KM1OR96B15Hw3U6g1VB4s3oSbjaUCilMpar4S
rP0e3w+c8IWvAVXGxXDxLe0pgh809sIrqUNYMVzUQPEgal+PG0Y7cSuVV2Y1rxWaAf+3EJY51x/d
EJs3zaIoFtomrK1Z08T7mu/mgdRUREtuB8BUsXoFIoqHHWKSV/qS9fQN764LOhNQp9p9pfHqs8GF
oaA4iGhMXTBEihIFpTf72VMUlltFUurszgBFCd/OpfSS0a1H0Se9nvmcpDUFzdQJEQSxnwO9UpNt
IJdPmTkDekIuI7yBMg+GSlkOvG/CaqRlBoPuAgvadBKKodYKjCeAXQY0iO2JLp4mX2Giiz7hbYNH
73IxduBvOHML5IR5YPufpKr63PUHdEz/B6w63L25TQPr/kNZ8hEkUzLejLO7w+FYrE3e6JbTfOfP
NII2csAqn9xafYZs157xXHYC13EqW3vu93xdwIIWBBRHIKsfYYe98YZHDKCUIPKEaX1y9ypJiDA0
L4wWmiYSbiDykssnWM8cG8j6avdM//vF7GSPu/nEoqiwFXcB015RIL4lqagmPoBMXPOO0pgYh4a5
RhbWO0xBZFZAVU2eVmHkc/cTQi4jjz54/P+UbJG+n8LKGzU2gnMO3midBHTMXLziCx2m0iJvxIqr
fD0a1+7Xwq3ZenGNKyVBxgPGpjczYa9E5GMpNXUSEb5YEyDKuVHad80LZvfHj0fhWojVQqHdGheP
Jka7ISp5wsxYaYys9L28e3zwx76hmf7kXQnLyzTmPLqehO8dAXtI1tpOHzAGZXHTJxj2jCL0sFlR
YQty+vrRc07YJdzjqPLyo4auUd6RyvIZa95URTYvZeXDWyeV0Me+JDru3c8cldodvQigJVflMCiS
ba4DiGOCHxwhbiPSpp4M8TarZ3VoaUG5LviG/QWoJ9JOdE4bC1wDq89fNauvSjzkgx9x/HFH4N0Z
7EoT3uBGvgWTcCN5GIpa1e4V4PdFKQJmUW2p0hBNKyIfUtLZGEcbF8KV6eAjI+nmyo07vQMrKadV
6BcWijzLaixo4jhEwd7OivKHmBEzNOwjt0YjPmsICJ20QOEUzxVENiWNquFezyCgnAQlEkTXgixY
ZqF4Q4vSM3Gq2Jabag7vTI1UowJpXiIdNe9dB/HOMRrlxD0p+DCv+HRc0Bo6RzfCye/XP8bIqgRb
loUVA1u/wmKNm+PIdCpMID+wYWgtAh7Izg6VlfXTd9+xFazRr27iJiO+PSHcRc7Evx+PPdqp5rh6
d5AQQ6+PEARODBQ/N1s1FzJc+n9WRDlFzuZtfDdzqM/ViACMSwYj3RSXBZV0ffYfhIDvNhajfPpG
XnKiuuu2CHSuCvjx+v1YDffJFwiA+nl5+mHDrnZqVW9CQnPQQnV3HXstBQadszFbqzeIq+0IKuro
vvHqleJFaKFW9fplPKiXXrkqV0kvHYIrsVI90Yk51/QMvKM4FxgLQhe63qnYr2wguZOWafM05t2I
/E7WErRGVjXYuo4XjacIbFCCljFuNxy51y7Q9qTWbScAQ8uLGnIPrREGDeJzYM1TbJPl3usFfqxt
N1xm7bz748nT7d3oOdFGT1LwfT8/sp5GI2uzTpSONp+FOGp6YUfXQQ02AYA5tjMwTnZHhwcmHrq7
GOEJ/Dgne83uxWWy2evKjmBiGzC/DF897ZlMf9+ysXmvkYgY2EfrDX+yRYahzItqYqrXesszG7s2
iRZbop5+rrPxKzyFIMlPDoYkCyM0IrbEbsW10LYEvCTdEJ26BPF9q4qtgFi/Umbabrg6cl/eq73y
MPz5l72ADCVBiTQfeFiGQ/83YxqJPWH+zpCAgEwqconhnBf95uwpPgZQLDb33cxghBOwXEIcwBVR
cZyQLDwgKJjsNL/PxgJ3CThq7t3r62wUfblB6xTZv+B77JkbU4aslTb267x9KlApc5f1Ye63qcy4
YrkEJELhlyzvAKFb6jBZSIWmxu+71Uxp3lALef6Tu1BX530jGGZJ+05IDgvBiy/3h6hruCr2Y7Jl
7JKXGvgokO+nAiBeopyFfn3CR7dR8kicbtqqnu/WuWxP89bzh5XipgMNfFWSv8jI+UIbXkk3/RVi
raioRcUmPJAVXiTFvAPqRk9ME7sWdk0swj+4GxgkPcw83i6LeBl0jm7PLO4x+qM9gf/laWQ4AL2f
gnJBEgb0sJbj9WzJTIB2WMWoPoN5NAVDKd8txwoPG2PGw6jeI8aXpbsN34470GTEfuTEoQeWXbiy
u3Lw1NBDWlc29SBEfwH5ETON7fet3tk4VoIWrbpvuxnrj7uTwFRTZLnOeD+njsJelDp924USZN0w
t/NVc87oo7EmWmRVe5+kriUnt5qj5iNjqo4osiEEoQu7fluxuUuxOF+O+k6pB7UDkll6Wmp76MyT
7NST2bqrzhUNkFN0XrSVVnMhEavSXLxMqSx405Q+tl1bHVsDSzMfe65RsOpuaeUgweV8sr9FukqT
l4fLsloYrNFChrrlSvlcPFEsuAdp9FBjjVOB3CHbVgWRd1sJTMQMibeVf0Uh24AkzfEOOsPZbSO2
VV+14tPRTyEvU0VQDJLBlNyBK3OqyuOOc8GDdu8nvCned+shlDlYnhTEOXL1lw9hHttYzvZyshn8
FyFbwec/k39hyrwBMVK6lye5Z8YvgjuXBAWHrQ7QFfnO9fZvuDRRsG4hqUo95fA47GLtR3nw54Ew
V3Q0WjvOF+7nu1zQ+yJedXIm/s4uj2M7QxLXIDcCVPtPIGxNPhOM4O5hJAQ/GvvnhW7xZDagwcUN
dB5EfIheD1IMfsbk78z66EOOTNzqm0HhJutMguBlA5zpSGp145Tlr24ULnK7OD/OJn8cZMhpvlV8
6Ci672qYH4hgOFs4jtp1HUBpRcqFyGfynaMHXmAtKr8Z8lpIJxLgrc2xEHMEU2LqQsaKUfKgy7px
9cL2OvM0SS4aL0iaYkB0Ze0QQBHWWdc1nKkkxZQ79W1HODQP5Z5dl/v38PHosTyrcilulL+uSSQt
i3yKmGzj4yo20dPJI+yvdUFqeffD594C/otQqE/IZfdyzDDC3o/uGfjQI3dIgq3uAkh29XodBgsi
VdyDjI6nW0ZoWT3h7Uy0KtvBIT7RHXGUYEjrVdVnZGdgOc3z/6ZRXWjXmk0NjqIyCjGq2SH+APNB
/m2ZwoDAAD0UhJ/naHNw+uhCTU70YgeHyCEH4AcsRgpWgO9f4FJ9tkQOkBJUbdvE3Kw7eEvQM1lI
lssmL2lAu4TXOolj9lrjVZzqtQ1Np08S0RaKTOK4qrL26K4ExmERzBBI406soYjqk92Qo8C0UHvv
brZDAulDckT9eU16RmAuFvt9tq0Q+B0jSrLnDRCsUokjFQdYDUk+01ZadHn0eD5Y6GKOsdXz3TXw
YcgshRoJxltKVJIUUZZYt3sD6ErashTNarmUsKsUVhP5gSxvO1QIoq/NU2qrnyzcrIL6KUHcts+W
hg0UGD4LwghC309jopLsnVzy13csScmySicKEMe1VJ/hhPRdjTeiFBV34mTZ1JEfvStXqkRVFyH6
HoikhyrAoLahfu5/biLSh5LCAEF6MyI08OVQAVJ0p+YXa0Q5IfpywXBPWzSCJA7SQLw9ZJO1qdbI
5fdnK5jggsdBOZlzqDJpnBSC1aAJ7HXd9Mb3DLlnoehwZHG1AqE+S+2kss9+ETXqHbkSbnYnaCjQ
RpVDcQiQ+qJ88Vu84hSNoNyC3TAGswgbIgjAnViRsvyvKVQpYdsNi8MhAcNR0AUWiwO8C+Zalbtw
Rob22/l1b8rVVQ1TyhxRCh3EgicwUBqXnjjlx9rKJvCY8F7vc/BjFmzOomsUExxnJ7m84LCESB9a
Q24PoexSLWzcIOWNX/R15FCaEXW6qH76JW3QiAUBvlrRi9ApPGRtB/fEp7tO66qrHLmjf0nqkTXX
Vbniwfc7xVQqP6bH6+yphaKauaLh1ZiCZ7GWc+/y7sZ1dIeynXFS9bTeOaLN/mLcB/gYetuZ6OZu
VrU8Q8bNLoFNWDQ3fBj9sTrHnyQ4KaFTzQ54RnCzdGd4ngQJGwhCesDk2O7K77OBDDzNRMR5CoEZ
0BEmN5/vuXb21XjsbmCAaRconaBorbU0q7iybb3+ES7uwTZHc4nRP2lMIYoYsYb4PyeR4sgAMs4F
Bit82VFGyCFU+vNZHqd0XVW7HctRZo4MZeRAixIWNkaFTEKB3gbYg1w2T7PmL5Njli38FDMqnReO
Rr0LXtC1pTrCCMQ5K/n3ovLJL4NQbQDqVfdeBwR13aERPfxmjerDbuh4KZfUev+AjJGMjb0vJvjv
QlOQeyl8WifdSc+fDCzkXgRn1iVuOBuyxGTlnjYHZJg8IDoRY1ovRRs3CGoEx8dzV2IRBGfJ8g4g
ZvHZx1JNUYst4PQT0mTzQiAGgMjeeREWV2M3A9l6eIBMtBsTT0zy2osGyt20YblH2lFQPLU2ekDX
O3QvZkb/SUr7xEFyIP4EHulDHHzZFKluOmcR/Zx2zmR1QuHRXJWmIddp8XEnZ4ou2XoiZ7lsEPNF
mSh4vO2vV8SYMoc+shfLk0o07ekXOJkXFCOMxLhd0I0ydwKnxV93IDU5d4ArpYMpeEzv6pX63Jpu
AFRQ0pkQko4Lz9/cDxFiV18A1PZMC9JsLg/nZPdo0mpKxeKyYRrW9+vYbnNBb8yAywqeX6Z+M0sG
oIfaUX4yohW0AHRdW5YIyzKdQlzwuzvKR6zL9KMJnw0bwvPbfs9sYfLvgR9NVmKlpqADsK3TcA/j
WFnlO7tmrgJROGhVJLcDWMqtZ2p/CchDdmCTksgtswgs60Prsxo4nXmjtSJVuNGH89T9he61LTAi
rQyfMngy6ol1Wa7W7gtImnzTreZ/bDx4HPXkSIYCR7GnN78OcW5dTiR/D0lrvU1jXcoYXy0X6zhh
yBwYEgHpo4FjThyB08StxgENUSVrYZk7f9LQU+u0Ahyib0X5AhWOVfqWiD+OBr++7PatGAnhKZY9
H11mW/x4UipeRw8Hmaxxwj/0G6MXDGfboST/MrrVTR1m4mE9vOiXiFhzGwem6IUMTES5zGdyRiH2
fnOLjY4Ebz4b/ura5DD/zvDesU5Wk8nA0qp5qTccLqkDWV1pnzeJ7MRxhQ55H7dfuIGy3LKJocVR
t91GmQ2AdvYF2nYP9CU40dcY6YScYmRWOznh2537tvj4CrD2bT7t9i6ShnBkGqbrTTy+RtX2yyAo
kqlHpbOGj4cYDEPrdQiQdPBnIXHnyRulCHqMzJaA+EcBOmMlrYK16bGt2j5YwusprP2tbdzuTO2H
n9FM5b3iFwHksWx1LtYI5YYyQCZZOfu/3VdaLezn4drAdsJPb5Yor+FkfKEyBhMl/mgQqtUkUNqa
bOx/sLF59xd0FQeytnMMPSbM0/B+K39xLRvm2SnNQ1dieSvYIv/7PcFPbA3n/h44F9txX1RRX4K+
IkSvBZfNtu+Dm0HzKMbuwNMyYwJAL7Y2bE3K3uVByA7ly9VDU4nvd0+YQDViQ9PTHFN643SCr9gc
qRDiZvpJevCp29pCPZLHdj/rUJoMWZ8htQT8gfED/2IZP8wS7SV3gU+hHtLPSRB1wGlgZ3D1obSX
YXCv08Ww7dSoO9+jvYjOXO22OaX2SNfU3Gyk1vMwfJrgSv4A7y/FiAJdFaelYK2IRJeKSTkIgawJ
OKnTD3UTq0X/742VVfiPtux4jgYFUAYcREiRcc5j/98Dzq6yfviOgwy79NhijrvczKox1aKy3vWU
EsMp6Nn8huQyWuf9ZRLy6rMcT5dhfK5gAb1C8NWDq/QqqlHQXNMxxGT68reykTEhzDeA9p8cDZ/T
c81zrByAn31T7BtTTWWOhzDneb2XKS0lZMtUcLjTpEv+BwUwmeJZvSqxKZuk6OeVebPWJh702ZZd
0Mpo0VHVIkds8X8jsmWsbSIyKVNdC+NOk9d5Vm84EDrJRYohiPvr8wPiZEW5z3er9nIxhdZxAxmT
5O0dg9cpyWOJy1pq4yU3j2B81vLhwlsByKdjSVe6XpsABbGob75M//be61krvwJLT7urzAXtc2jC
FWTS7ywQ1oDBImnaM6vtqQCyTCQFQZuc0l2ghStRZ8W6jS7wOu51mFUb18vRJSndjgpDybrr/FE+
1H5sigBfg8WmDz2/zvDnA8yP9Q3eSeyMN5mAn529cvHBCsl2KbYWo1Sg6gEni4Lv7khAGyCdEwBl
iVWQ4rBxGES/jLcyNDkgnYpJ4HLwExAJqxhQhT9IdllrXe/0leY2E4gCcRFGzOjMFUk6/B4kgvTS
GktfOr36kq98jRHQy89BcFonDiiiAqp3rzdSePOrbDL+cqJdA9qrEG0QguHhqWtxfd29mJRpKHev
H3uVAFe1PdzdLqFN9AVTUTZ1Sgj06nkeLjexVfhq468VlzQIUhvCCM+RwyjNbSl5ywP9VVmNE24e
EhrJNT1CCFqkry3GobZDkkBGNHdvH0fUzhuHCuj5WGXAd4/xQthcGkfRfHP7KFG+sPlD87xjG1if
4FbQkkBNN/q0h3Ge/dFOaA030BhTAcc+Ul0LAQyamHQVh8vKBE0tPLl2DhzTBxvcxJYOR/dvPZbS
9lXU+qW6d9ry2qnfpA3L1QagLmYEXAMxbsl2fIc2xAuFPz8Ko93YUeYRFCPsW0MBPMjGd4C+piiV
FnagHo5gT4mhVrBqC//AeQj4AVUrqhsFuhOYuTmU5vkrfkhLHRe9ctkRIDk10uBm7ExaZFi5fbhb
fg2COxKVbykKaMlBb+sM3LwiLrHSZ3DNuRuxqsSUDK956xlANTJqYCLAb1X1OTsqEy2h5W9yuJyD
B+/MTPbsWQNNHQehe62R6FMuhNpK62dUdBuykyennJ4etBO6Jaz+PXa29sZrfg4i/KoX2kiNhSlY
g/Pe0D8e5MoBgqFCOT5SVcMKuM3iwHVartJNjR/1mbNUFPAC2E3v8fFRQdcHP9mwSVp7LBaoE3p0
1xUCUaPGTduwUDkXr1V4grG5WfyUzihpzISto2+eoHvH3ChIXd4ezL16mEmiAVkAvmecVyiNfWHE
RxByUxpHt9ZY7xEB23KTugvRgKvPZtX9x7Gm8yTlL8futWkOd64vLDGNkqaTnZ5ALjuSskJI/f5l
CXPYBxO57oomCzWjZaXlw6kJhuLy9LM1J0ey1pAGSNpsT57Vvz2wKyExzs1nrQO4OI+3Vx+zjJ2+
FwIlsjXxKFiHYQJ6dREyiLhXFdojAc9kMfFuWS20Pfd2s8/lGp55WBhKwAbijbO/o3KmdciQVQRt
yxtx4guvUTejbYtt5Gd2Wc3IFXxIKAswNc+3XuA/ebrvRdQ4yAugCTKrL6SNdEK6d0XjGQC4pfl7
JDWTqU2pfxLDsdXWItx4Rt4QMb0qdWDw62pOsIpmcWNGhJHECeTl9h3wvZRBrLsQnLMHT5pli4WM
zCMorvJLKedgbX3is69upbsGl6R9lP07cXZSxntsuB1EWkyV4fKNDE1W+wIooWLvfoSNX7m47RxE
dGj9bs0PYQFlAAlVy3yVwuZ+vIn3inAYKBdXuwRW6GXd/1nFOn0A5JwKQH9Qz83M+eV7gZIuBpcE
+f6hp2I9SFruE89s2RF4i19osfwFkWxLwTBq/4kgAhvjXUl5j81s0+2V0DVqEMADb7LjUhE6bIFs
Tz8+BASshM5cnvoFcpy+9VT00E4hyh7MrZMuG2WNXWMWmb1wNOv0iRdLqZRynXxlR6+Fr5lWlyRo
uHltrL45Y1EEKGyCGb1QmfBHbPyAigVRBPioTmSPgsLe4ybZ1cdEZHbW6GfZuxLIOJDieGnd3L7i
hv2tZJHUaLYI369pMjeo0Rmt+Ug0foZ0yvxu2NZgwJ7lMyv/+q7fXBrzpm2WOqHp1NclMyT10GCy
irVWDe6OgXTHJ20Mp0EooETnBr39Lv7VnCsD2Ca3RRJGfQC9+ZEfiJbhCpPmO+OZ5Hl8Ab0diuZg
ll0ln6q4VMLYNzrXJ35nqFBhwHhnnoD3xWaFLR1sUtZ8BPI6n+27E786B1nCFgO5sqelVEW7GoJ/
PQN65GYZZSwfUZAAI735Wz+kfg3lxetVS7w+f3ZvijgSVo0rOi7jglagMykFYE5z0L/ziKS7Lahq
pkokv63qvKC3W80ceMmauyMgdsIO8Y6Ey9C3gCXoXnqZfLNdmo1Jrd0FdEBB6fOqN0W4NmDBsR1m
+7c5CcpZP7OfGSjvQi5TUQkn9arXOGLG0UPqUcQyub/g/1AC6TFs9CstkdJfkfSyabS/wXzXWQfC
Tta+PcevE9hBAFDsOfHEP7mWhMKBmPnDxGIrmJgLDpFCP4csMJ7L30PqhezZ+j+FOKT3rKSzWYMv
pRbfC5MO9uiaN5Opm0IQuWvw2GeVbEhNQDrQdvGoZCSL7LpTjLV/z7DMKRaVecu66SbC7JM5kec0
ekGyZh+o/P5grPWXo68UZSRkLbUYPedwv2va7tPJsiy93bRvEtod4yXCayPEv5xq6K1Jly0jVJqL
k3cGMm6e1aVW4tKDh6TsKg8oTHjBnibdozCbf+lWjGnbhAWidEIlxPpRfXkETMl1u+Y0Ws+VVK1m
Cp2PPrwtgvKuAMC8aLd/C8SqNrcxLxwBmu+26KKmTomA858vF202G83f009F2LhoL0nC3CMSww46
OabBXZbJwaVcTdp1TOAXnRyfXHgOykFNzUv7youpMfsITZSPoe8KY5ulbkQeG2DHh7QBGfuI3sN5
wjF9Y3biQ/GSn5q72K56Ov4TfE3L4+Tmu+oEIrLL1HbD2y8GAqZ8XGM72dBFqCOpVUDwpLyfUn5g
OfuVRi30/thbcmT8km8WgTAh9fLpaR/VZE+Oeg1qKpCGxZ8g05Pkr+UnRv5sxv7Bfzkb6agRz5oc
uQ/0FhVVPHtmdLqr0NEYXETQAaws/C9U21jdUh8m843uWjiv/aPsnbL6fqFsKIweSnAGzQuYwK+w
H2MeSR8eNenzlhvULyBKDpVTC27xRaGPoEcmIJFWEyjQzkwpaP5DcIBDUACmlWzEuLpv08GHgZaN
VBQNJK5AikvK1ozfFdtCMuQA+PKhm9Zpnfa6GC8n5B+xvIz8pjT2aoBKJL5sOEuPp17wLLLXD1CV
fCf/FRE7a8ZNhUDFanFpsIQ5vlOWsWNeKIhW2GM2TKwZ/KMazuOSygGtmvdSTLl+csiJljsuaohL
lACzRnwVlRhc5EI089gNwL1PYWfkDewrz5kKcqhlByOAHgv6BUu7+Y49PcOr4Yd0rW80AOKS1MmW
KgchO77SLPlccLTRoMMtzmB3GMsWGe8PTcJ4+kxg21mT+G6DfHusCIeCIupa3Xw5IvzdsbLYG8E3
fklAlbZ71R1jgO+hbL7mnWF5b3EKQq9FZUYvDvM3TtEr0+uzsncoVObmINiDyGh0cdOJQTHCTKvO
n18rmme44cp5D4/bqe+DdkAF5MbolLaJjpwyvsjo7w3fJSW+bfqFwr0s1zdRQzZVAswAEf0uNKyx
z4Ym33i5+gs+30snT+aMvKFgUb7+n0lCmZprUl9XlgRcWDh3p3gjwzbpKjLotUqkJEeuAkUUNjiJ
hne8elly7Jf0WGtWZGplCi56OuSlYObZ61TkvfL+F2YldLpYtDhaQI5QrxHzIMulIeL14QQhlC2a
RC5HoOcEaRQUXrRjk9SvG70Y9qGMvHRtwi2O62kmMau//WyHWwOPYyy8BhQDDhj0cLEFBca71e+4
uDaTohG1q1xaaJ5qBWbjUShaJFY8yXdxIhSOaSALlNZS4cFhivvZhDVFnMsL0vNEXohAFbz3o04d
h3AB7RdtuEQ22pdb9Idob7xDWI9Xx1rOPPh3WZR8DbVBFqUkh/r0+W4Xbqlfhmd7CFA5dnL+SCYC
zzK2kSEWH8m4mJ4ecNWwQ76G4SPnIKfJfIJqfGEe0EqEXedNtG3gKviRSvOe5ZEsRpyQa1MSqBLA
Nk/GmeGXfQBNW4WPYCgpTosElIfFwvHmuZtSh+97XlxRiCE46KmbEgeogmSv/qvjx3Yeq1SAoGjY
qIZC5z11EbqIO4+EfDvds1349eXi+eTBdKCiXEskTWSW6FR+Q028pbBznfu21PaRlY4nfwDGHEBq
WX3dYXbXeIEvO/H9qJTwa/MIbQm+Y79Mf5HoxOiPIO+Z2nJFypg6bmOqccnCeGt5KjUHPTllBoqo
YdPRsINp3T5e9wb0wq8Deh9OPy8vBWLKeQ9601WgEsUs0PN5ayXfcy6wmkVj1TDINu9W3tDn+lp7
LXeIN5L/54T/x1L0hyt2K+mMLDrrcU5Wl2GNwVQzcgjksdQHqdOWa0hLcxVR7Zcu2TgPV3snP2RX
zgoCLmjMMYqpakC5N8FeRIgBZ19Md/en/KN8F1xkVv95NNQJVSLp2nFqiZavQa9LIsutYsDqg3D6
IarPqD5JXto9HPDZX5y/I24ObS+cJ8JzkNbAWkuZeE9tu57mravWWXrYWifLYFk0szV1fM9Dsy0K
k5Qq/hjzYzVwVly7pacIu5te1yeG8rLfbw4Pd9Yd4PGBGQrZpD9m2Lv09a0juR5bMgC6LCA4Epxp
9u3L8rxXq23VvMVx0D8ddw4hzmmyLeEwBYlLWEq+5DRrIZUD4lNvJcvXLf9xMBa2HJ1e9MKe3Laf
LX5TiQNIF2Oyf46xnWvzQ0BgZ6cgGd4hAu/zgbPth6YZli69Agcpw+tUGmQa/Pcq7Mw0uajs9YV6
3/+gkeSVn3v0dhvF0bWI5hfyleIoD+9XwCAEwromzoHMSD+KXgz1r0pe9qejAx4y6L3y+GP1wf5j
BLLDzyhm0aka8mbm/tMWL+CQGpqIEpCTC9g6PquP+SJ2p+exlz3zius20tzW4CzaY4T6GWeevXco
DL4XrGC5fGJqLwjkb/967IR4YvpPycDMAiteGxJ5h5Grm/neTdkfKw0biLQ5s2+vwy9ZEHSepDoy
+Sy11/mRmEBmC+OmN4cKRs6F9v6AqU3z+EjldLGMF1Vkhl8CC/bSlvwgT+FTQ0PmPA+FW0unAx+F
a3KNc/A6VSTn7DSckwh5FzuxGwuZ16y1XssIW47GTRoTKhF0nvojNuT6CjjOWjErMERm4V+QyUmb
Bi+ORgTw7y0H2hmz77ERhJoablDqxegMs2bLlnfSGO3TTdVU+PHjtC4lO7010z98ndkuruqebdmx
6Vh6ii9c4/MHWzCHnHxk81XK5aU+Eh4jTsoji6Jm0+k58Hy0J7YBTxmpkYNaovaHqCoA7PTHZccT
ER2DXI9moCy9NUwWUvDzyNZYD95MZ8h6h48vfwp9rPJTD2ywUBEuI3OXbNFa49StajNeZImlaZjc
pkHG7y4w56fEz4DvypNyPyxEGNriZFFMVnk36Sbo2GYXKWI0evZRSo3buc/Ewic6qFCLOCm2NJlu
46lk4LTaRIhj0cmEstXUeTQQjTStRONejtGwdnfDUceayNfdnjjxoOfNUqB2vOgeYy6GJGPda9Hc
6lNheTWpHHGRcQ63K9G32qf3eZ26dVWqJgWeXgo/VCzkLrVsAFSjyrRO4E7RrjH3dXW0Jcxz4q/X
eA6yLcNnj9eSRp4itsSYaPilKGmgWz8PrzODsgB8LJJRuOuwG4vU9biUjOj+So+0i/CVJKy4rH9U
+2N28sxxB3G3SpUQ5KmrEFzlDPjqcn/pqQvuRy3l0ulWLSuKRq/KCCFaN2u4AmZJYPgeHApi4K0Z
mjC/1OfUukCpbi+Xoo8MyeeCcWlBvg3FI4/VG72mcU0IbVHo49aUUUHc//UWOe8scX4zV0Rq9AQw
vWW1OtSD3aJ5HfDjGlOOFLZpX6eWWQp8Qqhww1+fMrPh2Qzyzfyg4ES+kCEr97rQDfKKEiqJLb20
q+OyjhZHzbywBczXQrcVF400P9gCDv2O6T+EaGepX4zqXQ+3fnPcdcQguugYgj5GgS4d1kEOkXxx
EoaJQ2Yp5Pppv5kjLVqdzNTJm5Bb23wNojH1lGooWTXp1+DiZJDJoRRFT9TcwmtpLNKhUY7OwxI3
eIMLKkICk9IkTOriL1dNQ2AtMCAsoClh1Yoca9m800Qpm1EDAWiJB0nUGSiVcA1aWPSXdQyX2L4N
t0JLVFXjrsTvJrGU+br7LvwlMTSECylAXnt3HyNcqWVRDLFiuxzwXrlUdScSlmZbztkTPGlCaSvi
5XOjN9qW2FL9I7Cg5iZrqtpP5Nl7mZiXuq6gcIP/vxydRlC3/KHJiJd36n9SaUbp8HSQUcDTh/mI
fDbqQbXEbaCwc6JWobgXXJ8M2dQ7CXIttk3d66JGf6fHhPEdTnH6t3LzBJVojYzSLgvZBCRBnHOa
7wvjq23kdi2Cw4GWGvWT/IFdwVoW2Jd+puJR5VAF6dXb91zSZIj54TBSOuIdhaCr8QskJ/IhIk6R
6svKf58VSyDcemzRhLPV8IeBzDDVxo8TxXZKVHpBjWAhWuAu7pLNbO7DdEjyFpq8ZDCymVFUu0Lj
h/a77rZuLjX+DJ5r8hi1JjYERXvu8rpfX3wSlbW2JReGyXoxcEr/sP4M0+99jT26bL+Uyv8rNWyS
39mOpfE4gzlYIZqdOqm0WG8W/SrO0aKBmg38bPhPCDIcuvDExdJ90cyDJM7jW6aUxQT4HHGUJdtw
JlEYSAISFO1oZb3OByVZD+rfDIEQJ8uQHDUmnIJy7J6/JlbAxwe90flv1RSntdTxfogMClNfKecc
f3ndH9RH/e/pP417K0yTJ2P51kncasWUKwvthnRgceVebk6k+fvZT4E0uNPaWmt0GhUqi7UkBgi5
GekTt7gJQDNX/WcICHcEhWU8as8qravLUozxRo0ubMFQCs0EkUiYG4gw1Hqgzv2ZP9oKsSL7O8VL
scKuXNHP7b9U8mZ0MoJKoHGaccVn/m9MzRps+osDtiPVuX+k3McrObp3RUMhbT/qTkAKtMR7TAAQ
yIOeRCoCSFIzuWbNJz3H7KKdhU6qII6aKPdmCqSVt7UkYXBR4yAqNTRw99c77ulTP5fQH6CGej4S
2t67jke9DPponKg+0CfBETapf4SIJQ9OW/9dII0n3eigl02HY5HIEuWXrwWRedh5KPGoD4BoAGG8
UuvFSay62rIedoI/MoFCGlSAHaASjrDYOdd1qCyG8LhLQ3lZoZtZmqw8wERIfwkgOk0Jhmwb1+Z6
r8PJY8lgAy4iNgTrzNsp689Vuvz+TxsASN4lXoocyJlbt/tfDyv5T290py66tYxyixgNmfOtvAsy
342lXdPcnCAY+W/uDqNldIPVaQI0o1Lq4PtqGANG1I+Y0XoRdgu1YlkLpwGJ4LDzff022VlrbUYL
r7ipaZcLlHhVRACF6pxIFzTqs/Zy5QtN0EghyK1/FAu+j8j9qs4Wq1nJVv8mJ3AIe28ayuLmnM7g
+B6uIXed/So+DaAM0X7T3NWKOZa1uGxWcNpGKs5jThA7ptg5lIw3E+4RN0g0Bu2Whde7dw+cirmV
orFjTvGUsc0vZ9Ig5LrgNR8m0X/m0E8tzlET94VcyP7TsHPP+sMGVsJ8QQAhmVsOBk28SwtKoGe0
ZniIcaunlCgxP/e701XkI7lGaCe5BosGkiWVHu4cK8+QjgFNsTzEldYqer59VvBTQijskdZtLs2C
J/VEBWzRe+ghPi7Cp/0tA96jn/u9P4R01dvM8Zsw0OlKMlg27VA2b+5kR5CQtjZ6S9379sHdAXyk
vLPkINV1wY1jAWel2UqQQOP+tKlJhKkJ5xBix4WxWAvNK93yL/r7ghsrlM3zgHrpOMPmPgo9S2/Q
KILNvKjs/iAH5rQMiJLDSoq6P8ADX6CM/k0aH1CMu5lIk/qhmLLP/Q0aVnxvtZaMlGvtjc7N5fA/
sQQr4vWp0KaJfMh+TWmQVNrC+7zpds2+fRWyrLvg5KPq2uyDhOsr3dwT+fuy69hn3Ia6YzNu9UfC
ZbEfL3Gr/RSIdhB331LnH2dVSNiId/7MvdPNdCfRW85Lq56qcBQH02hmSWIu+j8puFSzn/VHSLzP
iWxNPdKoRUbnQbUovpjSjMPIZR1GI2xgDuMCKE60QSyqc5OxvDYE63A0mNJ/IDAgKZpJIYOYAv1F
pRO+4zJMTi+lewr8ik3avOoA6X4qihvdKgk7Qot5DIIvZgm4ZpQ6NzJL+GhkeupQYOaJfraz5CNb
NuG/akN0aC531lLNq2UPxoV4EG8S7LfsrYhqQkDM56EwRyHewSoIO3wmjoETkCw9CNjLhUR2RM9Q
M2YJK6My7l2gVPt0AJgg/ohWratt1m6VhF8PHr4dlYgTzOxTrIUfaiE+Pdob7okuay01T1Y2akQG
Q6OVOd1BSoQkznO1Blnoe9dhAq9UPy3TZ/fi2slgbH39MyGj5W89HAhekJNOUL9WuwPJD6KhoUPu
u3wp5gXVUqhjWqaN5fPCQ9M9FzcKMKPO8nOLdmK1lSV4bTL/L8pn04Li1Sqe4MWSWzCR4kV7UTAp
c8f5bMcsFjd2wQsBGPlI1WO0EiZz+ciro/txv/VFDmrLfZ6QPbpHSFkifOLX7qn08ccbo8X/A1R8
cDcguxF4/3fGSo8qsZKJa+qiIVfRb5D11R0/Nu3IBanRCJRXaFfZq+xvvndT0AVY0QZ1drAVnr7Q
15ptaZ/j4plLN2veW8a2Yxe8xMdyKhQVW66580N71FQgaTOzFmzYqqupPsyTaqTKmNiBus9dqkLk
lxBvaPEQrd4Vltytq8tCFl64buDCtNpisMzoS6G34iUxIVslgH3Neul+mJgAo4omaoZFwmoE8up0
AVlYy2730COTn2h30984P3NwwTo54Eeh3C9Mt0Ew6r0yrdaGQmOszhWfkzm213/SE3h7dij9/kdc
4mhyqb7VGUkhDvGRjtktKkkdTMwgp5s+2CDE8X/k2k6zcUwng9lVwnI6iElV7NSBfr7Xvn9LdgXh
/1eDmJ3MRq8ZdjEOpFW1RXpfGxFlnsQza+mxm8KbHiZY5MftA8sxFqf9KEa7tM9LgHCOD/r5SHLA
HsxTQX0/d63Hozw2mpNY7TCFjC/yqYuS/10WtMAOQQY92uFE0tLndmI7HbG+6DxGS8ri2XnucAEp
wthme+grr/mWG5pG/tJEALiWBHQFqSKA6y/oFYt81qHn01OFwDPqyKSX7+nTxn9lM/0rDkzo2j4H
HxVL+KGbCpUz2SFifydEfdLCyJeYj67m9lKVXIOJve/0bWBH5D83ImrjL0fczKXlTtbjiaX8AsR7
Ilped+d04KIq1nKJcyeljUulniQZMjaHgeSZArx5tXbfW9j7X3RQ4uHLks5fCe+afuHWBnvGQTft
7QJhosyvdC27FQrK/iF/P6YlQIVYbHO3wDpqpnr9GCLoovHWtJ5p2PKgQAOAnxbpngpVvCu7HEkp
MJ05fJPVid7FeM9s/xJlln71IGYXFQMxJYkaa9PYareq8HYZjDOyJ7MHMJJACG203JEmxysxWe4I
kpMs6X2DmgfuZ2+gDlTvUVIPOcjhAmizxVHZMdeC8sK3j34pO2f+pfBKznAoYPPpN6/Wv0JAH8SE
YyRRNWFwKaKZODb57qOfGa62DdwK885moHJ4k7u/j3DdX80u43a4TR6FFR6EHweQHby1xHXmvGqU
YhN8rTQVWAPI5Y5c+3YJd7rf+vzamARX+TzUmEt8CbXMwQOD8igN7EEDKR0SwXgd/iV7YWx8onHU
Ub/Kw5Nt/D4CSPYzSjCXV+5YMwnGFYCmhI8l7l+E6xkWN6MbxieebsGPlhZnlrMQx1QSw0nctZ4/
iq9E0qqUKKQ4UlvKm3VdsY/2jOL4sI5hm/nXdK15g7tUb9ezEkK/4lNnp6FWx273+KFYnwUF4hhq
uSFF98OPUwzd8P9HQky3bdHg5YY7BCLXLribvZlFEVUaNXb+Lle3LT9jVcKUIPmj1ypDpzh9n3If
cAHVYv8nseVR5vJyOO4SApSOFoAu+VrMz1EzDCLAQ516SUF884pWNkWh6/IKxU0nbe7BLkG76uCQ
hTZrOmLcyC1vscAUkYa9Ikh9EoN4TlDTPewI+DQpTni+f05Q5QNjLiShM6YShMr5HbYOD6gRa4MJ
Z1M9miMzwd28nzxpYkghoiMjlc7FtpDWH3WfF26r1HXXzfGRCkYHkhFuZVji9flNywNp3/cR7tpI
o+m3jpxqmdKm+dP03kZgfrRKZgGKRNzYUQLPswyEqtp6r91GkynfUDTJG9KkuM1jKkgcyOgGy4el
repwjQYft+hDErkQXurF7F/ohQgYTBaiq2bU2iAtyAlvPXJLfpz1B0IJ5zKoQL4/J9A+YQ/XCGBv
lZggQgoMviYMPwO37GcrCy2mLfyVRZD2lxwuhK16wNIT78omog9qwl1/di62qGu0onTIR875Y3e6
pCEPxsg7MVOoV+v5nhvHruY9bCZ0bZqfvB7jOUjxK29MIlVjyF+iFD0/2A6XJYZTdXfoSLW47EcQ
YQkoOqok9yElhhcUWWYzIOhdSt7zIy3vzSJpVvkK60T5wwIIh/Gy9pDDvi0ZIpv1UvYIc/bnk3iH
SqWvLthyTE92VBC3gksjEcwiYZvuLu523HgZPv6xfb9UfAlZx4qy7mSvbFnMd53zM3YBhyLjg++x
F25J6LqLS1pDGVkOU95FC7eg/dDZh9HCGlM6UeGLVwbrOiA3IpqjztmslZPwBEMJvMr0nFyPibdr
X7n5qurgQcuTLlmlQi4kv5gD4Pl3vmHV5Yr9ofloXcKL/10SGnea0SOJC5fw7VADs3pcSAd9y4xf
GIaqUShVN5u8BIcNHSqXn2Z2LFQlvhI3NeS969R0UoRiwREdlvmoZ0hKFm7nNmwz/8ylboRhVYHV
iKlUcRZ5escPCE5zXnd3nf0CrVfKYW50vys+rrVVuLo7GuJpxf9JAaC1eNdayRawke4C+wSVxnu4
OH/GCg6+lZ2Io8mt3JpE/aRyEX9hgcKEbVMmP++xRybfalfUTa7w5lTDI1RXMGV4urwqNWnvv6oU
q8Go7JaEQ7ZFD9SR48KzSpHrcz1djGfX47yCuhL0dB+DTmCYL5WkimE7SgvFIaEDrtOAO87k/ntI
1FUPjQg3os7+ul1Atnxon/8QL76sb1gA/VhgYcTpGMKDYdMVJzce5gEI4Jti0mBVDBD+KGRHpPTe
OX7joHJQGUnqj1iLk7RbNIdyfw8HhHpJz4MeQgsnCfoG+Fmf00kIzzQa+4APNsfd/kh54Xjpri7O
c/l/TYIIFY4HWkaVJyN1k2eOXp700PNl2lUSt6D45/k3ZdDhcS+x3mt9meE54lj0z9VndmC9o+B5
eWfV59OxSzTCOn3IqP00XStMgg8ldCTpkolLs9Qytb9l642/TvGHCwQ6Bw8r/VW/6O0eiXle6UY2
6KdoDnJpQ1SJhIVIRptFhmf6gJpnWVhrbGU7okRicUiAJ+6wQhDx++KZ1k5tZB6iV94hSoy9Wddl
HEM+gAFKIFdM8yO7z3bGxakIPQFIHVkeKZJrb1EH0ZlWHi7s4UpbljEQS+KOMfFzK42pRw0d+SOc
v9R8oxLwBTuHwv5sO/0LJ0WPYxRXA+dNYVZJHMPVSnz/daPLwTO7Wy1Dw9Mad3XTDtx00E13cQ12
hBCKkEBBc2bomf0SpkrSp7oZZIq1yUys2COqYVosNQ5SJ656T2fGld/lnymDVuaeOUnZBEEJH43L
KLNj3jNh3q6PlWfb2eFkW5D76NQq16sKVD7aqivz+XBQiddKdEVmB/AKr0cXUFZgiRkJwk8oXUKF
S6yafPL1lHEhsEuL7Gmk9OY77e9XcVv/HmnTxqDX5GWSgBAsbnS/H8ak2EnmyX1CWkWyIr3vLPWs
ckiRg9PTo/Ocbuw1F83reK04diUzKu8XK0IWiZ9bSqMM3Ki1WDbOTEPqpRFKdAtDsExW8jqGf+36
iBtu1lgI1gsM40pJkFRU+Q9AZ5Cc5i+zNsEZpuUr7xYaVXlRqAkZBpNm/zdAr9Q87SllarDDbeXv
1piJxq+kFTsc/TGulRwxTOja8AcjR3GvbZvbWW0ewnHUd6zUOLUFYTWCpjeV7MN12S5ilWM32CHq
6jhJNoKP6ZWDuLwBSLKby0FKWGPP9CVCk/Yb40V08a4/WCw5+iM+2L0+Q5TEGNC9QVSyPlV5+fIK
UupdT8tuj/cYT3yx9BMCkdvTEOlmNB2nUD+brXrXxyBxhitE0eP+cOFCAupJ0gemKWglxWf0RT6B
zAL+UxOnwbNmUa+bnYVJxof9NyMPRTo4LMpfbg7ECmlASW3u13ERAKAATiGKVU4kK/okDc5HtUGe
4Ht0pe0rctF2i9IJKRXRjC8G5nYBkars07GXVcIyLSpiZEvpfVO6B0B7pMl4mJoX6Dx4+o0bZTqq
4SZjHULnBGh4OIpEf5378cpTjvaTHgc0J6ODJXrIpxldYD4lBaFSolv5dgRZw8SB6QTqAipmDld8
XW9O+/RIz+hYqcQeiJWvkPjOa463CvEjMVufIxA48UnkrL40UVUCqBUJQRtYPmQ1o2X6DTtbdWbc
sGAjzzQZOMd+eUu24OErmx+fn77oLKIAp7G1rOTOm0vvbMtAs0BJ1jG0hwGPq0bsPgQPHqWKqOlT
qiFF1QKRlkyXZGlSiqVNojkXIZwrK0C2OmuCKXHTqNGYD9wn23iJJau0DzDwK0sPvE1J0xNoI4SH
nklcD4ny4/5u0z6PxTF1lqATWGblsBeZmsedWuyJH8y87A4/rC5NbvQ03ggR8tHncJ/Iu50b/nca
eC49q466S+EpjtNY4AANAjOKKv/u7Lw4hdvx0tglR6FFmFsW2oQG2Pbs5uZCSaNjVyqREaSYIpMt
QSsiuhEyXv+WFsa3JAVeuQp8ZQ5kvB5hi9B9kXYlT1i20xC2soxTKBnj6616EMtRuvS82+WMohhj
JqBR1eHfV6+9o9tNzZPu9HOpGgfdRU7K4zmKXAXSwFwYH2e4hueGhZohIhk/FuslzmVxRm2N1Oob
RNFBL5MvxN0wWDrLlutEQyEz0Y0IBU4+Cage8sr0ixFqCbxsk/HvlXpZnqdwF4xim8Luy2w+fXvx
RWFQzNs5++3RGbJVig+M5Y/ZIqeNmVIlEKsJ39WtCnjIeYMcn3xJOpAGM4yIqhF/aYBdzOlHHgu6
LzTBuK6sPZ9cnGe0BgZGGWKWd8WC3h2YpVG83aK5IHLp1FzzQbg7kSrg+JAF4nm17/20YiiGskQ0
CB1VWkdLs36eDlijR3Wj5UUv4lcd1VGhvH6NzI8Me5+jts/j8Pjtd5uMVjSdyT/Rw6z5AHe9ev3t
rou6FWe48hQ6V8sHTCDcywN5W7Y/LagmmdXD+7WnvZ5A6+NJ74AKgeFABgqn7rv9IgFQwoH9mnfY
Knv/XqInizmDgl3HWL5MZyK+0Wul4tfhL6LIU83fgASwBZPM/dW15dFcIRStyTfi+/dIAk0F80nT
TtFjvHNcfx4QCuv0kjrVMH9nBrXhGjssnBk7xu5HVp3t7EiUS/ykCMb43PEb+wuSc8tbQmN8rVTJ
n6cjguxOrnf0NwnJCtFJlA3GNgXeU/FJhRt/KIOgwF/OWbTjctF0Imj9gSPUzUPhw+tNc+H5bFEu
Fcdk1za5TU/a7nxccHe+JbvRDtvVXqSVuaNl6WkpopiyneK9B8IvMmLFmENNLpMp0BCwhrkpFlNG
WRjTGMQPn1v09S9zUB9uH7iNRi1+6iboGtxP00C90aTC5QYB65dhS6ObMOn8MnyTlDt67/ipSbxs
AOtarm4b9/F0G2FxztuhoBmEjWjCA8FSQhW8HbTKRwEfoCigeJbWHNzUkkgClN7GeUQExzkSol3t
Ik1lgk+mbHroJVo2pzYEB/EeltnLwYVCFHM0m9l/WAteOSqeiOcaNrh95hnb+J5lc6c5nxMiF97Z
RzyRuWL9DAWPgUA8fxVMQvEpxlltZ0wfNVHfAFfRjfy2XfMzndTgPGg7xGXbj3cTmpmYSqr7VDyZ
e1BMOHxw9i2jNoEHZNqFmke/0020SQzxgptZfuqBHndZ1H2CCKXKtkSoTyCcWPM8VEkn3FXudI0W
OwUnBRAzTh3hqDM+uQjXx4AYe2rYDK1BYJZ8fGIelbzK4ugPqz65ZSz+wGQLC65bMcddN74vyeGe
G6R6ZjiTLNCrDLGKm+/6ySccYpgu4iAMdfEbK8tgs4VbUNARDKytFqsf3p2v8S7TPBlyBP3sUYhy
ARexlcleYxlWEf4G/0dC1DRWyRUEHVm9najTJMmwzbuTG3+Skx+WgwgMSZt7ErFRSboiOZf0AEJu
foCakoQFsUFWsZA3h2U9GBhCWjZDRQHq8hYr5Z4CLh6N76+UJXykK1lI7t8Fqf0JvbhD2FgfXAEm
8Js8T5GFEZ6vp9WElYsOEGZdxOamV/z6WIml2r1vn7tiGR0N0r7zDNWAF9BC6FwV/s0lnEiF6l7n
d1c4vbJ+t2k1SrtxFiz5rtuu/C7bf+E67dyOOqhpMX/+E2n6aXysuWRhYfsMhMx3J4Ed1rlK6G/n
mhWYdaVHYx/eLr115DEnU6AguS5Z6VoY5vInRIHkwNIm9/5aP/zMMMeb5Rz6nVbt5i3i8gaARMxH
YDArcW1+nmBBjKwLEwdTq5w+QnC6HC/lmdHqPaBeZZ5Nv0sZ6skrUZB1KSt61iiczj9OgMI/IT3I
ZTyvAun3JTc09wA0LRSugWJYa7HPuQD3G0yXf1qRp82Hju13VAzUuR3P7A0JiS4jGoaoJRRXiEFu
gV9CGBoa8W7/lNH/CxeissTpHKesJso+/4KHkDmf78qWW/lcmUk2w/dOhTHGf+7mQD1INji6sYs/
6O/DcJOnytcufzSsO+/F21qU+7DJ/mPrfGK9xzLWkUBvRK2NhSoF1fr7/b78C/FUqBm5R9hV+8YG
x0aBUw6UYiGfet+0eVoojuCUtBLpft7TUsh9+IlTejBe3QxyLVnyfevf9SiR62ACuD1G593SGQeU
RC1ep2ZiV9WsVkyDyYPljGINqA6NzFv0GrYCPY0jk7dypFxlVW3Xa0ueLCx1qyp2rNHTaDkADhwI
CaFFB92lnB+SOY/hf1zYt6D8GKNi37URH7JIOegpWBC9HrsbMacUrztxu8f5syWObuqp5X7POHmV
Sdlh3kQCuEs+jA5yG9ngngulUanDfozjU9Pxa5vbKyzgLcVZ4DWIk8gedHHG5bF4/n36S0+BTMiT
Hs1ake1XuHdM+BrUJWASTk0L6vfdVpVd/1/g70GYBEzfMHZ6Z5FJZ9atmYa3G3G98e8UQ2F62Gx2
XEoUHc/Ef+kSPiSIN78zi5Mz8gZrBik4DsfgSiycy/ylulNbSHKCM4x/x42jSpLaGgxAtZAb0d4E
9nBzvn8FN2YM5LEf4fkJpK26iYSTy3iNkq3/iu/dN1fxFHkMhaD+T7IbiXUb3cOK329n37ZLJGk6
17S3HB08/Yc6G1TEFuCY3/weRj8hOfv/2DAECIsNDnmU3mVvEdXBPhNL37gQVMKQWR7kXbKcgZmX
MoVN+olQ3NMOhXgwoIMDCp85xr/zoF2aZVJMsgo9d4h9WNQc1AUero2QCNOsai/7vgs8bLT88Ib0
fDWF3hg7sYwcG6gy9Xiy4OE4DrhaKiXU7LGM22WNqOaP8aVJbnaDQNLy6p1sbBR5MhaBxiTFYorw
4LjvAhwvWogum9MlBwThXXGxmgAuZCPl5kpWO8ZpVW3s9nVDG+aldSRZyfgA3Uh34enDpmuE5rZX
1ATyRctKLLv6ECU7Hq0KdxrAlwwL0bBsCyv6Dd1oBEScdAZPnKp+kPj7B2zs+00VlYKbQXAWWXyW
t8NLT3QcKsPudPajGvVvNLzSyThrtt0zn18msNOBU2AeUmqkK5JqnQh0e2BVueIaU/6UV6m+fSoE
a3dEkaZLAvnkQl9pSxAVit52dBC/TUina1Sb01+pozvyzsMG6IagXAsVBTkhyjEFeO/C3a7ygFJ+
je/6gHltlzsIAif8F8Ld3N83HJyST/rG4+4/iif3mQUYDSPqjRRvCislqBPaXQSWwzkQU17jQCrv
gtvPRtte7RKfRGxTHnoeblO4TQ5MQ7qRUXBz7ZbCpEhQAEuHydYF8CExp1PuLs7tAdcJSrsy+Tmu
HnRGFV+vgIAdYUxdwMbBdrV6a302UhcwXXE0TnvJLUc6ww6muhc5jKBI/qJUaiE2mbd4jpY6RVNN
EhmCDufqkfxFNYny3qZMe5pocXFqp4XzPwFbJMjLAwjMhyQEq/ZLfp9CLkuUD1ZW2ndqxBqtQTmg
1fbWQV89q4omReVMA6z8GvZ0ADKzGyXiZDtBdAoGzl381RKvW7h5ROFF3ecpnmeuLYEG1WLkVrev
4HQoW/Ny2BSSl8hUUc/bo3t2odR2/bqJnSmMwR1O15n0Z7qic/vEf/PvyuVV14JE+CJxoR48o9tl
VFpER79Y7qurpB4p6AWs9woQYFGUKImczBdUgGgtFHKFNiXs800Xq7NSBZJnPH7aezEPCBZX1RBk
jGTY3TuFzoAOCjVL5gxDgav8VJYAntqVNDlZjGLSEHvyUi3FJKuA6YdvMvliT1gjsGQRj/tYHwJ9
6A9qYAWi2P68QUq3UTkPc4eTm4sN6j2zVyL95C60QO3mSimeZ9zNdjUo0nUSTnMXc0Gf3f9YN8R+
OOkvOxGOsOTJcBmG8vplGRfVqr0fvV9gHpPKOlNRZqVXI+K7uV4BvmKj7OAGl2jR4sfeMVm7TEx7
kM9g30wwQe1PKflb1kyKfwcuCa6lP+DGhvePzmSukTrMY4HUcOS8Nj9SEnf48LnPXZwGvANdUIH7
I/hJErd8ZkrpcI3BbJQmWevaUD1FryrMG2ZWpD1lDwodudSRPR1EDmHd20SEIOMbfYf7Trh3fvPc
LYbnhZ4w63VUEDVHONAqJNTp2tPAkWx3UJQQKt1m5HUzEEtnhaWtpxIlgjGt2PORg/9bB2VTuel+
M+DtlIgHv8F4YP++LWH8nA240iZQJS6wm2i6igX4YDuekDnEFqmclhY+j7KIkcc3kYVVv982ZkGs
omBB63ZC66u4gTrJZlSl9ccbG8kXz9S2WMn8OQACZVA4MM0i3qekZ/W0XFHwZf/S/ZL3KICo+E02
oeX75WozllRhgXr9J8m/tf3I+VlEDKalEpmfvm6g0P6ogr8vuqoYRrjBnUhPZzaFT3dsMP+Ixya0
7ZIUj9GNisSnoLnmbqAcLKldSQZHGbJcjJtK91Yk6/eqH4Hne/nqLvencmkMe2SadjO4sj6D4HzH
YUZNn0qHq7yP7xUY4du3D2+D9bBAJ2VCkOLh3aJCZpv8ZgvK2B+BRxxyAnSVTS+LA4b9glxNxNLk
iJURCOd39MRl6iRk6t+2/tqpkrWNFX620XYOmPR9UEYRH9TMjcMZQ6Ota7zH4H9dupdDHjyxBQNt
dVporkeREJmbO7gwO/G7rIVh8H5EL2Yn/af0NzNE+sbb4AvCGtJ8hoVGeqAq6VUfqxS50IluwzGa
zf6f6sJ4cHDxTHw4/oQpGa25Zm91K7O13jdlrXO7l0LRIw3mZtjYiv0wAgaMWyzl6mufUwyvNV1F
VQ9PdqZfqdrCUzhNHjaalsS3I0A5OghCR2VkCIOqhzKgt2scLa/milOVFy/4Xt8//LtRbt9zp5Oo
xnQeXrRJJR9GaxgGIcQMR/2Y7glEa+KkmyLJb0mahbR8ADZpOjU/8sjH2h0Vfnw34bdyoCyp3UGH
4cUoD+Kw+f0OX2QjoxgFJhMjG4ewMaNcUXGhwWJd33DJuhDoMG9M09cCkdgKvybpcea2Vg3xwOaF
2rD+w7qj1XBdVrWN4ngVEDuTT7woBkGy5qioyUBOoEuHSoxRr/+A2y+dSG9jzlEXId8CzdWfjz9X
gwKJY4hEfrpp6BJ27C2dH2latC22tttjfVQ15u1p4jt+DrE30X7mmtJs1mSR0eQs9TXjYCdSkPam
Tb0dadkumQM4iGks2e80jHEQrEllbdiNL708yvU4AhiEqdEsrdLFEOvpQ/eAo+r+tXIFJtAWdamE
QGvEciMCwqwC6TFc5Q37V+NnsOiiEJFXfJtXCKmcHvuOHaXj+fSOv19svejFF+bNdbdo1tJDPxdy
LMm6z80koiymP/4giloir6SPy+eSAqXOPA2N3IgLAOn7GaswPthifFQrWRUYZeS9JHUtzmKcmZv2
4c7G2M+e6KN8pyN1BgfCTLlZvavlHJi92swXwio7fgn9kCAJVIr7FXRwJXWU9QNhgh0iLDnp5kSE
UpFbz3S0CoI87606/vDBVUAJmdpquZV/3xET9lU1b2rnDiDFFXgJ1x+XjbFhlL5/SLxIv/VzKRK2
nVHAMlqev4ihnVktSqCB8pEVCzdhnTNWzX5f50Y7jm8J5JFLF2uDHqVg41wBaiqzi8HvfoU8v+MI
McufigvO4jc6bmvJwzayMG5n89Trs0D2pLIUbtdNLUbFLfSHg5DyNhZ5UzhPrfJzHdr6lwa8l4EV
+NS5ZOrtYdEgeZGln0BL3mrJS9aSrEEvAA8bz0ZhbO0tuz8PplZaNxQYZkS2mHUrp9w6YyCZ/WEK
Bvi9bLgwAfHIGt8eXJNho24+2opcECWRF+0uCOFdPZS7Zs8ajCutxZc81M4psyevcjjoQiBs3xnp
rUDPEGYlKoD5yf1NnSr5EEpSjLiAJ83K5YFCjkH5Sfe5MR3ICFx1fJyFwVRpF+dha4INmTUFU3Gi
ILaKCuBb8tYZUawt67niINKfrWWQf3CgcanSeamRVq7PFQGuVtvVlVV9Qlsn+FMs2XwTYunEnjyp
XISXnaFUHf+qo6UtCzr+unvJRIkMt89wzxQBA0nf5eK0e2mPapGbUSn5IiuULOLa1mFpqP9lTNKG
XmbtEu3GYH84dnh4VyhLA73ceK63YkXqPeGJ7T7EsHNwmLmg3AtbnY7HuaU59j7pM+IQhaWXSuAj
5j7z50trbCpJsekwz56tJZeS5MH1UltPLF4ATYnVy36HwgXGWBe/BJaJ7+VuUuassIlGZ6rEqPEs
DClquIa/USb/0w63aa5dbL2R85HQ/L7sbJkzVJ2POoMZx7fdfhqRRY3l1rIfauG4snu/Tt+EGSQT
eeQg+2GZXMUStzVnYyJVWiQML5oMQBroPVNANMBeSQYZ5VmsX+E8byjxm9ZCbb6n28Z0Hx+/g0a+
zuAo3ydsYh5rd5vF7lImzhHAjMENedFihrXdzcwewlFZUafCKycDfLJTFtXzNTniJX0WUuGokaCT
6GSat5cArH25fvMnlZMPBiyn/fm0KLiIyXg6aVIjFLl0dQu5hcuwFEpO992cUSA+9TVJ9e0ltY4G
K8sHNoCv56y9lv45y2rV4ZwuCckPmrU3/nSFuNeZxa44oxBaJ1Dm5fWtLsQDv3WMHe+Eidk0neKq
Q70lpgOqyehLVgnZFv/wnVRX1U6UI5Eb+8ep+rXco40s+dmiebfeA4H5EMwVtJN3PXEWK1VOLYNE
CQeE+aPoC5B+hqKKUMQXYhmBLkIU05cXcDXShXVwIH4Gh5PqWhTmfOPS3izGOTBtskHCttBFJfrZ
hKH07Psb0KU7MWeDmeX0dzxyy5kvJ6wTc4kBQ6AAkiQByCQ5b71CF+IxOUOBTjbJvuB2tkE6XG2h
ZleoW34r8m/owJGquSKJAQD27W+9LXejBUjbSCwHjCjQfGVRiYsvC9NvdsnvOUUMi/53l88L4oRm
m9AN/IbNhyZ+P537jCUhxWuGSL3Ld9uyEX2qyoyxGniAhzRSoAwfpEoK6yUbqRx9fWhE1695xmBO
T7N15YmPuXYFImpGtwwf83zK1me++jODxWaceQNyuRZ5Eb/WFRhnjU2qpcsVKai0Yril1yO8Ysfu
/T0KlaFPN2AKbY/W8WRQSqJXUz3Ci3el/kOuQTDUUHKXhwbrJMp4mz4i4RXJGXiz2Xjer9k1xYP3
d8/kQUU8zdRu2Fz2Tj2XPfu9VolyfLYXaA9Pf4l4m6NzjQ0NTdtr/qvwL3LVm6ie7wjrutvrAhWg
MHGMyCu36cIQHEZpvjmM2JMyZa3ruxT4H4TcHXdJ9ZeEy6aRD0l/RgTi+9U8M94e4Jm7VRoI+jf5
Rr18x3JTkO6GqR1sxkmWHh9nEsPZAU6WeeL6N2XHIOHIYali5mwkbbEbCbinzsJquspYVPUKvgeg
dcUsZJBuXfZ1fF2MMyJgRDFWjpd3ZCC5yrY0wj+ss7lKay4JLH+4QlhrzMBFp9W9U4j31N7sEJod
Byl/+NP9twiTMiuyHugYr4Yj0um32jF7c/rMixQ+1otADfQ9g0+z7Ti84YOz5QGXkk4s8TnnOGnj
4Jpdph0FOCxFpyQsafHnRP1r2oq/q89+DChqODPSShDWZTAWZCZ2Bd/R01cXdrJE1E0HMElDYkaC
EwYPgwDKJedxxoDkjZRlXs38ed6hXHdPU+W/WIszT9iSIH6KmIM2pFVTMBgmnF9lT6OYGc3qCnx6
ygGMGN7n8avaRUfn9iMcflYGXRC/CDNVWNmpDNb/ZxfSnsDeAq1Kp+kteo4qyPeZDKryjqRDp6Ao
lhfyLZBSbnOTzr3Mg8CaFqqP5iqI6POuRNQPKhUcip6isX+f3KvM//s0yDifRBHi3RvxRUfiOMIP
TtyKI6B+PPH2OaeeQWZ44ucJaeIApSL2hCFLBbSpGlSyjT9fLxaP+c0MuQai8IUHhzyIsqLsvqlA
jSqkBL1RzSCE2UZ2lEpEl0BfEON/ELxxH2fkAt0IFjbVFv8KR6rnEm/qeRgLliy2UkFtFKtcibZZ
P03KaX8OiXjtyZRVRJfJ9VwMb14S+Pcsqe95PqhJzWszpyUerrSLMkzAfxhTN2XJNe4RcoCqHE79
DPLjWRajrpruF2+8BqOFf4DuxeNY8bQ//s9qLHaY4Gx8TYiKSnBo3j5ZcqW0jYdl6GKrx2EV7y4T
YQjGfjySy/Q0pvYI/6jrc5kPSUTmhnZKO5ebb32CstK2CThRlc62yXzDdqF2csFP2rrNVjXX6qNX
iXMaNE8u/kDO1qpcISB//84IH2W9o2+jmTlcDX/QUnzStDfEKrXglrHnUxnndnubUihmTWgQvhrZ
0fKRIquHwqchlHC4hbeVdZLsbkhzKNUCpzvcHwSDQ0NCq48w6qJInaGe48P3Phw3Is0nyAB5EPBg
3HO5tpOBeAznQ+pBBE3+wRakNxh+nQQgR62Y4KW5J8XiefkJDtpnASwiPjZWp3+LV4gtsvm4styX
ILg5J6W5c7HhAEmDkO8Yv8NLWldNmJkKRSWAyE0yMgKdCsGrgutdsVZqTfWaggDbhfOZVZXAmrqE
3ivEqqgzH109OV/eWCSllrHJnYG7r4WWE+IhbK6PKjNu3uEIDgtV1WSTw7OT5jEIKaZkdGuCPUvB
nsn/zJYJ8Q9tTFy3kNXGcnmNV8qDRDcXvuJFe72Tzgw39HbhNbEe5Yf4fYqijHcvrSkW3YR3LAsz
aymHpDcwy26zOairUHg8Gnz8A2967WtUKkfabmwhEpQOxUw8oDpYybf9bB8piewojFBzRPGSy8b2
FFRAKFVY4THQsN92YQxcaHBDU8KAMETuF+Hf9YW0oR2cXzCzOBSA7txTR9CAYx3VMQjGI2idjcFz
VM4CTeYVtmbFrqnoV56RtugsQUXERE3z1nAbcaad5/wpVHYy8dja8Purst06l3qNz5eUBe7xvoo+
Sfj5vodNmFivAi0vV80R6IgSGS40+qrVCY33GP+nXhgm/plZf9sBL6gw9KfoQBQmGhJdq+CGahm+
n3ISGgH51Ho64gHS/dxfEiHg2KR9Cq6S6h2SYJPEwd8zY0zxVBX8TwYCL6MaxC4kQU77j7M0bmDy
MVCFXVcw/L72ungw5+y2L7Wjce2Nqn2PkOKxFZh4HRQAJufYbHWlj9tpNUJaMqB1ZaK8A+rU48Oj
6rrLXJcTOb9gHZpqir3KOUjSYY4v1OBx6ozNMu4/4+2bEszpasv7luy/9eh/SbywqgWlaJAI88zy
KzIAufQiGOeY7tIT8B9qzkglyqTvZYW66rGpnVuMgAXTkatkZjvEnUEWhbSLOVrPHySFFOOy89pu
XLysZPjzE3MLebInOzi2VVGMwiQdb60kfsKkEZHT94Lm+Z7x2mTCQXa44+VB43ElCDub8/2FxeWc
8BlwmPxLRU0jC1YKzelUNNAd+sA4+BenVmH4C+5UHS/cgYlhozZg4082aN9x7/y++QWQJxOT8vFL
W5XZgLHi7nmiiENfpKwq1Gqx6ljwuU+eWXPP/nYC2/WKjKf3IKuNeqU/8XPZB2JWKzf89zzZcXUQ
WhTG4MH5g6PUP1IdI64MyGltG38P0xdDS5x+pfURMEG+BiZ97SH/O6N//D85l8IIBXvj7f5hvnQD
pIHLwOemL+VE5cB+K8bNR2cIEdTaCGFX3nUXOczfOvecOQLyfOKbIZYQvg2vBOeJUDizvzREJUK9
s66pplr8W56n3x7HXsnuAloiXsuhTR8D1VSXNtNH3m4psp5cEIr7y2x/lGNupIPdOjuHAa6qAqjY
5oFQ3zJgkSm2XNxbIAfGQKoN9QW5Hx8hxNt8/UpPePRAr1CyQOT7f5Bdlv/V9l9Qqtz1vr0laBsc
Nj/b87rxU3xjcY/P8YUp7V7kCiWjFUUmnB5T1gTWQ/XDcg2TMu/gskw2eFam5y0sytV6brwosPz8
V84u6jcGcGM6rKixGYsL7Z4Xu/y1qpihX+xSbr6lZ9yt05ajRo2VMX1JUwH7JJKmwZ3Zn0NfmdFb
P9909sei39zs/TjHeQfsFe6SmFsF9c1n5N0sKxU6E8pFVAGiUJqkicpo2VW2SnV4COfK1BO3PbTl
5ZUnkz3/6A1Dp0kxwskSKFQqBm8zpaYC7HJsEwRLPkjaWdYhAI7zF1sTkXjBaji6uFvEQpysbe5f
YjJ32lsOEb7p3j25SikbLHueQYEkAMO46Pznww+d/mCLNr2NiOZYRA53wmlWjlEmpx9DpE4XBROP
OjOK7EYr2oXFnKk5ZysyQ3PeidoUaLJDmcmgmASJQmOa9xLFQg3ltYQYMIAb9eXYVSv8A/qffzSi
fSLA+1dNRZQgVNdpO+Zse1PiXg4yhYrlgXT9JzLuK7gxjErCE65s352YZ6v+1f0NOyEVs/8/Jfco
jXIi+XH3EX7EqCTbi2JVqAYRzqP4n+40DxoU0AtB1P54hHdn6ynwqSNliEcjrb44szXhhx6Ce9jm
xgt6Bnt2Px48wpU3ZobXkFypr7sRJFwQI9XX+nvPfyf1s+tTA+3QwvkxKyTT3otEQmaMEtUSrNgR
2QX1oSBcFDJZg7e1Fkp2wLtm0madhd8zw0+UWfYtKn3NfR5uSJxDUUaTDJFm39djYXzPhAXTTDXt
S06etDAeoSfxPMeUXKct5p5FdMIoU0Ucnht1+hLMhSzYMg4VvR4G1dCmvIink9zye7lOwP4yz1zh
gfwIDOi9ZjsECtoVGD0Cn+96Hdk2koNIz+UVSghpzYisLW3IdrFf7e/wpryWbfXysAuLQ18PKSMa
tsB55lLOa1EnZT0X6U0bfWW9rGiQ2kEwxKm8dniHvLTOFtjopoKIIoF7KOBzv7d796vkbmgigtGl
W69pIlz9I+KEiIUSXbqvHa9MzQe0yGZv+OANtxL9LOsU9l3S4pm0W1j3gS6dChEEHny0OLDPIq0M
30pwE88IJlGVRv9pe6xM0aMRNfZRUUqkroniu5rn/Tq70qxHMk9xg4YolsUQ5/ZVXNALYrhjrn+6
gjHIZruAZOaqzEFBfz0fkR2dMVO9Ff19NDAJvx6LevaFb6uVIs5yStaL8lBbSBLYYUMcm370NG2h
IJSgL+xgABHIfHy+UlZtqAEzsZDjmVsUDhwObpUcJzBOn0iS1DLrFlEAHKWKd0Zd+e5fu4jBEffR
WN1YNbzs7ofPl1gkPEPcPJ7vGAIUyQURSRhsxhywo7rL88DrIak5aWLmO3oq/WhEScGO1i4/7oJM
Y/n1ta3fJ9beAbs/En7Dw/xkk/YtlHqatpM/bYGmxgwDp4mFky+dtzZhJcyaDxQF+rirTWl9XrZN
fANXgPzdzygbyZEdq4E74jRVPfMtk3NiHLG6OahoKdRz5d0Sc6VhmEwLjzQSsKrqK2A0RjLJGC2q
OP8Mk+vle+1nI14mJWUjYsUs4IkvnzJYZb3XM1v1QbCUybLfol8wD+IGB5wDFjE89ZIeH6ozpblC
GEIikEzwmgMHEU/g2qTh18ogW0f14SO/LDmaWeoOPyNt3xQHB34jX423mfRZH/8hLgFj05CoXZYB
gJXbD1ATliRoa48tvzS9TRuzY+HxbeFBruJaAR1HAPc/vj877gujGaYDFwD3FOD4SOkCAE/OpI49
PDhVZ5OT1Liuc3/OfxT6d2o8gUVxutfFiFvR8kEvUcbtKF1dOtv9Z2PoNtMSJDZ6X6YSy9Da8qHP
cuPBsiyu2OueGo3IeOl985f8jTtEdTErdPYz0WVif2RbzU9VbJmpolSPjoepJv/Y9S6seuf25OnO
ol47W2sn7huZAhBwKW+k1a4oyoiOMa3jppCa7RRbgYeXlJwgE7GsZ1BjaONIShflAW0Ey/JyA/yj
fD2Wy/YdG8UMV0tFtz1aW6VFXMTYxdqOrarQ6dEMlkQnasdyMKFrLu0viUbV4oceTaryLL9TPk4N
rkvzwmG4MseHf9hHKeOEwImFom2F933JvSwqUBW4lYANwlo4lXNYquCHt1iZOHQkkJDioBEs01RV
xzKP7xUrN3MTiMR0EbrOacrENGkfPATSZkTletbm0d6iu7HaEcyn2XOQdKUrVkvWxZUxQrWkOlzr
2MXZif4nd/kYYoEA8l4QX00KFpeKRUl5nQNczq76WQr8ZGnXS0xGDLm5luTWUCTdTzN+TsSqdiDK
eyYM5/jH54Youp6A927L3bzMx0O8oTnFB8KxdTvcdcQI/wCBxD45Xjnhqeit3I4YLvj4mfBiV6sv
bIcLZEnSBIswRE/3bFby0p+wXjWhUBckuURuxxtnouO17I11ZatZQBvRTFed4qLVqKnXWTU1uTyD
/QJ+lqpJebUEFyQAuZgP+lpeTNd2vZU0q5Yrj3XzdM7tNMmsDIUiueSojtss89kTopWMhHdtlPgP
OHv8WI08ysX+qCabWku+cNc24BCU/l0kkjne63rSyvhHSHQmr7AmGwPDT+cxxBtwL1Yf0jlKSVoE
ANMsECn9X3rwz7vNizw5/PiKVjcQ4wc60jdm1CWYQ+9Q82k19p+UoRChFYO+AopN6jN7vAdD9KVd
Wo2JjZU9NvCYXHRgQecjA8jttGawTQXuL9zOLW0zphzxzpVNjGB4uqJM5tGpzinlY4QqGNVUx7/W
sltxjc7aSRB22FIxptt5T2zeqdlCf34S0HSDAouWgZ3IcENWO27kD3yo/qT1KrxSXwR78ox5dpBC
sqTZzReUIAneDA130lbJOTOHNSbbp9q6OC0lUig6icBkW2GruaZFzdDWU2/c/TTG04f7FADh08JX
M3QwA/CnJDLD4NW0UgwAbemIqPix/wzisssfjvECa42n+1IThlcAhlY/fZFzKg5rIZNK0tmoZMYY
pQ7Q4vgcXJGiMFfzNElj7BZCEWyRijcSB2zbORqGn50BWuHB2Aj2yYWiLUsHp/k1KWCmIG9zRY9+
BDBjnxNHtXtlGclfyYymX5NqqB2vOqaoRVQ4eSCx75TMWaUHA/pVGOOrORl7HuyielV4bWRjgbvM
jKTBhFx+JlFe86FkF1Rzm7aysB/LiLL+nW578Pcs+YgrNYAaO/dR4kESd2SHMj8YTbma8AS1/twp
qSe6UeppgVSvSJ1K3PMmM3tdbjHBCEbVaTS4lBRN/jUfXaJS6HGoWZAJWQQhd1DOSsWD2rVXs3bR
zDJcbI7erH/Rly+DCES0DOweFB7c6RbwPpxE29+wLa1pGs7CYUb5XozZjrKtDGqighkSxnivwmCr
UAo+LxIuoTFWy4ANlwwgl3jnP6R8vZBQ5Luv5Ab48wKiNFXYD2KmbrqsRLqcEA7QhsvvM+y6Iiqb
sFkLTiAP1otzl8S9VQZSF0AZ97LnxXwbXuk5VnbcVo4Kjj5qhxuVlIvnxYkUG1eb14LxRw8c+MlP
e5c+5IwIqtPWR6ZwsSABVU7c+piyn2dlNerN9ZSoIYB5RLe/quKU57pVcBm3x2RRro9GSwpQjFhH
cTSaUO0h23pUXCFI6FfbZvITnfxezGEYM2RHOTiIWgl/skZgFOKfsX9cQZ4iYU0WLXV42/qhpQUR
+xk4wknmmZM8rRs3zZaUN+UrDiu39rRHYdG1+VgonDYNoB95Fv7Cx7qlyYtokeWYwDmbYuDqVy6j
bEAxM1QVDkR2JkaV4rIKFKloiUR3i7qG21v4JmXtB9IHvrdw6ndc/YX/UpvTv10+cJsK4fRj6T53
Qt7uU0d6iZpm1ZCHnaP7lWagI+FefEOHjC+9eIYWcE0MkAA6996PnqVsbD+jlbCpYR49sWh4ycQA
W/aCRuCuS7tOLhSDOYS5bhdFryKxq4QKNLWECbPUR+ZMsuHw4io16UF5XxchBmU1FHE8WHbgL9Ff
sLFfYCnHZmEk7q1+FIm9+Se75ZGa1YqtSKQj9W45a5FUBBqi/8gCpwVn1xe1GNOVR7ViRWHpdImI
bODFlzJxMJF+DLuAaGjV16s93RXbr0mRZGnzs8mB8uHibW7sA4fp8SBM/zVA6H53yfGqazPDzFMc
STkmRnO15VDVXpIDZ0ZoQg92pR3GF18D3RFFoL2r8HicXchyH8HrLYhbCFMLhYhg5ebBcJSXaErI
xM7KeQHCxyFenbUw3nDDYtvrnKPhsPuaYornKLSsAYJVrVZSP5BMBYSk4r5qFv8kDk9aPMz2gP8A
fj9HM4p1KMmnd8spKPzcK+K8ukid+6taJ4Z98mJgE/ER8NaK9QVXj0NyLlL4gZQrQrB2w7IGFJnZ
YyVo+e5KqsQ4cxXgzEtpigMYYMDz/yYny+f13xHMy+KvV5Mn8RFzzJWe9zxUDxIZP7oLlHdIwC1j
mBd3kHjviaIe7fOKS0IN4aCTwjUsgTv/UEowwciGtn69HjfqWKcDy4wz2I4Kgf1qYpfwzQt+lKez
r8JKKUJtQJnHJvBJdiV0XhpFL0f3UI3eKsIoNrCNqrI40Ey2szc+l8EEr1OTtQGJMRydoXiM7tQe
+N1FrhrWLFzhE/ZEuJ0QcCBAVB2bokTk7AiD3BOBdIExNpEmza78VSLwraxOiC7v5wx1e6kIkYUH
atC5cIuUS3iZu7Z+fLQgFXEnMW+07Q/TNMfQDHQ+XG6Czm5Jy2fVvnG8k1XHJB4s9VZD7LIyLWrx
gBrYafM7196b3ZU6QsqJrQtc/DzPlLmiEH7Yg6C/USmTQBp5usJNcKLTty0jptk76We684drsmiy
5qHvKpBIcOL9ylq5s58wdCIi2NOxcWWB8j8gDnJjRT8Zp+u7kmFFZxk9QXDiM/XLYmhhDrY/bgA4
4/oiE2hnkdKWabMqyDf3aKvSvcEpuPhXoVInLbPh3OVQyvncO75fGwm6UBCmmdcyx128Mwf4Jx+8
jFZN8iIVCOliigArall1B1JL9xvbx2zFfSmYU0UlSk/j8dwN7nMGeDtSXdeYr37eZIZGFi7Q1Ug5
WRWreHe6DE1UaCdf6XhsxlNhMvJQVz/VmwmyVkQ1zB24+2QKa3ZkUgr7BqNFalgaZgrW97v6twDo
P7VdDt4MU2dKkwy13uOYjgvlXyLEQutx/pSTN7Xj4UeHII1xD/darI5QKcvLmlAQSoD1EhFb0c8j
VC/p4QgQKf0tPDobuiD7Rk8ZJUmuR8mtUBrJi8oj7eQDqrSfDJzcuk9rsf47pX/qshy0NmWi8zqo
HavyF5BmD3Mm7+5LTBpeal7tl7F5lznb/62xkJgQYEBOVNE0qsNgH1AcZRLHaPogJRZL7bGjcUOz
4q/IgZb5FJDYRs4gC4LtBSTFKaxIKA8H3VT9ZqsWoC18hwjR2J56S1Mv2c7tpmU4Kv5uHPKq2gfK
4bTqffrbfjwpWYz6QCfR3BQSBGwE8YFbQlllB/1PDCKg14a+LQBrCLYTtsT9hASZOUIKGc35pkbr
dIg9XgJdebuCI1C8AtdMYf4Xt9cpm8JCdTFPPRa3nHElMYsmlEGZu4qZvQ0I/LA5pXRzGTc3eUz7
adffu6/WhzlDizTpTzuV51tncEHQAZkucGghohn71hj3JiXm6nLFV+TG79GvV/vxncfvtw8uCzhz
EA5uiovwS7GG2B+L0PqYeIlRDsy0D3X7myipfhN0RDzrFqOfh8zCcEzVNPp5ANQ7n7I/BEn3nRog
Ujm4d89bm77tPxtEoBqaHt1r0/OZF9X9rzaQ5s9fniwWQnSA26/zyt5n2v9Z/N1OKAqCmbQ4yT37
Lv7i/y0gonfp3RxWubu7NnS+/tuoEuT2J0qrHFXBz0WEieniBunomiqZyagDNm7it6YThHirIARv
5cDRhoa0EgIjAlJLdyEU0Yc6jZm5rgWnhYKydqBmbiL8QTjIDS0SAv5bzHuPJNyyWY/eJgi6Rm0j
zLKaU5cY4D4kYk6Z51Uzt4GRQr4aFHxWYILQsF6DQor0BZlqmZV/iCc41p8+WVRuj9MBYpcroZOU
xg6IS/wNm4H4qQ0NIjY6okd4L4WCdOvfJj7WCdoi7y7RX/rVFg8SIYZs1dt/iiwlLrJXBqfJaahc
oT20zXshnHwZRP2krRenVePJlWPSf6YfdTFx3HfuuFA9xUOsucO05zag0+bdIq50r5MTyI3D1tY0
AByCHDpZ+kxY0P1dcoCMRURe1lWSqdsO8uq1J/XBKw4t4yWJpZjRKnFNHL1AGVrlNf/IFIUSp2bH
knX7WTxXRZwYN/Oqga/06fRrvFcH4HDWq1Kn9xuoZbf3vE2qsBBG2i/mpFa2QMqocRnk06lxvJ3v
Lt6nKgwrbGr5AKuOq31RedX0JMo6h1vf45Js37l0ahBuncHRT5Lqu+YfRB3/IzeXYBiPiJa1BitS
3pHQtx7PU+8FbQ4P9vu2Q+UkGNaU4q6AOS6pFD+Lo9LU+oD7fTchDMmuTLhAgsmBaevb2kD9tVZW
qf9+kBPq1dXpeMTT6Ae413S6xYxOOmKUg9Qt9mLueH8JBFTUBKFBv1SnWvzwDZroJIm07rhPlS4l
sacQ9xwiGJiNzJk+TkOQoLXsxn5WJ7MBlC5OIoSWR61MIoJk5KwTt3Onbjnt4ssH+5mqZjsHN27f
yQaRtU8Rii2kByFOhZ5F207nFTUd7naYUTHKeW257W3umpVGR+67rE2edspVcvBSztlH34/X1B1P
DQ/88rRJyIg8EUj+shN7KZhmOKHdHL/ylLK9SQREjZiX0ozPpAzswhjoxBFL8friepf8uiu5FjQw
82+6ff8lKFzFfqJnznIi9snhmU6WIC8lSiksX2TxzjNjdwDbOkvTptue3+0Io6ZQsfgFBbyOHGYz
sv3wNyMbNO7Xee0BJ0Ox0r9YMLI8jhlBOlbp+T9fvnMOZQKTfMF1zg/Qh/DVzZFuRmrXzO3H7IfZ
d14oBBCWGI8gUDjyPJRwQqgrBpP1g4rZTYe36hCMLigIpPx9UWyBtLT3G/U9sXLK6g6QIp5XJ7Yx
8hTEzHvbqE2hZAc0qGwQ0bmjnyLvPguIFTZNPklae8Vk4zuEdfP7eO/JeTwAGmrtuK17Sys5wfAY
l2jJVnRULtCtAMnFTK3yQuGAdZaNVN9drh1FxnZQIrfy0c1d+pMgwhqA7kkZrpJMwDUr2RLn2xAy
/v8iAteeMXZJXrgA0JoKNwbCO+kdMV+Yj1iy3/AcBAmM3jqU1nQseAS4Xtk3lKJzvTUKJJqTV74B
bRRlHxXeh+BFiAHDlUYx+9O5/3I0jh/BNVy9d9qTfNCQ5gsHhqRjYCVYDR0GWG6xbuWlp73HRFcR
AIsOoUllvV8gFgxoy51zuAEWBcvkLR5A8GlxvchvFn0W1E4OCtkZdT8KoD6CzlJ5Sg2Ir+BFx89D
hMz+9/D/kdxnl/mkSSu8eyOJXuZjQctqwHnikPH45DKeHZ0shwiSHVNSoS20CPB+nfv+RsthQiLh
+bTLeb1ztfOXHl0dV2d+QcQ2zA3qQRgG850T9dayY1PKJT6SjJSeUM+ScZyAJ0TUR3wHrXEq19A/
aS56nLp/wlzwe4JMY3mpHCjovTdhby94JkjhY4l9MT9AVJgN32k880dlCoJHss9jyQ0KdSz7HxMG
NuWBlnva2nT6hXb5DsXKCL1UnJDpKbVQorG3gkHAGwFoOmzK63YxeZAHUibdgUfmmfAYt2vqPeyh
+Ze62Yztd+RiEWPRKaqRR9xT4lBkx25nbgQensh3XGJjNj/MJT+6nMWVgdS7jFCZeUUpc6LQdGo4
OjnYdoceCOvzHPb1RQgDrUEbOh0nQH/DWH7yVXkVyCHNbwWwyw5htOEw5yt+5MOpP+m0xh/tdblR
vWpp+a7KXna9Nz8dnV8tPzgWQqCQz62TFEJqeuQlrOnxHXVWH5Hn/7vM6R39XyXZXafdM01lZYE4
cNZSNJgrAhBk9PYJHjlRjzOZaF0xdhgOleq6410XZWy+0awFD2upJkHeviqhI/sQEpbZE2mfvPKI
9CVyKaGbUFR0i093bBIk8a970818NlRMnFAlfHaZ37fhsILaKoEYeUMlJfhf3kgcqXphzR0bTBAJ
K/jaY8sxopoYxZGw82KkuSv4N8yxw2Sv0bBoPe1vgIdEiGqyi6C+c46p2yd0cmTKyWhGKgQYcXTp
KFntIC8Fo0QW37pyg/JRUUb24zNKPK19tmSTZJHEDdIZqikiZ2f26B0UL6Gb5NUmgbiTrD1R0Y1n
tBocoDTw6+SBnEOlij0RxlgiFWJg6++hA91zcAbOH0WHGYbnBM6jqWr1UbecS8vWpTPO05CWvZnE
oEh0NToeIfJAIEnFRto0tUutN/wmzj8Qu/Nyg7YTUyHz6QMQlv/YrT/bx8Kdt4w2NrSnY3fgVvGZ
pPN1Id7dRxfHSXu821vRp85kVBZpvY+Dtr6h9slfQxS1gfkE3hkCiSJIG9HJjbmzpg2jU/O+BHly
Zy9FXmDPvz7c862KXwdl+UwSp5o77dm9SKyuYCf3x/oq7M1zeVfPOVIkQMlvH9knOp5QfMfcvJFI
zn6qHpXkvwM4nTmtcOIKgivCWvSxn1E9L/UHAYCDwYljkDVwHiqgBGWdgNqItfLnDvuK5Cp2/z9l
EjyGHDmAjhm/zBoiqplEsdxmZWHqmibPt0K5Eb1uq+VVM/qckYmf0nJPHNEdmmj+s+VZU/gdh+5i
wpJvbgXiW0ZsYYMcoAGd5sx3L+odzU9I7/xmjK5T9kWiRX2nOGISl7+EfbNofM+oUgNKLW1RtYLs
kfnbkDYvnU6mlwj6WaLcJvtckjmKPNdRCpX1BctllbM+/oxmRM4TgU8d5xYpAK9xNSp+1XISznkn
/0jQxGiBwgQhJdiUEzCzaAUNr7lPFzUqaY7sOCsNi6LhrllFfiOouYGDelt8EVPYfz7ksxlVoYf6
1S91zIjKQWqvdwUhMIh8Bd8lhYJSl391+PKHd8XdteyrFlt8eXS104sh7rnVnyrruRahFggYKc3K
SYL25A8lfluiC6pxe7Ebcq09mRcc3VBddmzZ5sUUxIiRJdbcc4pYOJQZZoyq3zLpttSsjNmHSo2g
ZI7iC/zuAl+yKsEncF3m7gX0qOPLwdH2aoGyiXHoGZGojtOHgvDZ/JWJzjbk8HVS0eEVCTS/LeTo
UV2Gt8W2p/66AFCCxXSS1xRsaaQ9DyZ+37xtynYDZkzlWDnn5t8dD7+phq8urEIO8Wjzdw6cxoT+
iY+6KviPo0U+byXaqHxJNMjsNjjIuA+iO4nzXydjFSPB3RVPhzm0CmfMYLFXEjYBWoABoPGxRdha
4LoELBwusqSxZd1A4gH0jxVD4LUbscYTXIAsjpNcwDpgUDYPQOodpVZh8FYWs0i+zIiK73coPWU0
rz4oOLwOGToB0gL/NXKICYx/6FDe5/6Bu4Z+0Qsd/tosdla4RiwEJ8d8aXH5r9TFL74RK4eIDRmU
KEObFefxWQpGaaxlmVs55mH/2oUdt/4VXRd0Hy8oTQ0eI4evTxdGU5KpjgO3nHHDnPnQ3rPxO1nF
Y1VNkZwd6iWm9ra/UUxDPrepUxoOJwZ4M7GAaZ0w3AD6UgWiytSPMsUdnJlP37G0/9AWjcXKfwDq
F51cjRqZ8Xkt9DaTJin5KeIK93YKg7dCl7CX6MyDqXpwYFDOzv5oCsaNmSxDUuaV42KPlGNmqa29
3zxigNL2/gyNnlA2RSc9emodj/WQmNFjSoQED6z3qv0dFbBpmAuFwXlqRBGWvVGQFNt89k34O45G
YfikXvS7BBz8lsz5EOttKbr5WAqyJFwMs4AcCJRv00KMYritnKZKnzSftOcz8RXakp7sEPCPfMAR
+ZFmDu0GnUazwV80st40wPe9NG7ebSvVgrTjdQjaSndB1pqE4dV/r+1QJ7Nqq4DoGlRSdljt8/+m
RpP+XJA5X3/OgvY5m4mBKi+8X4NxRW7cyc3dMZkeyqjVM1fGFx5TFVD5basgS1qAVTfq+MI+155e
Lc7o/LGIt+Mn5bFuhfogUNb4xz8MLIuP2ZJLqsihUi4fFdgi1rvc3nON6686QoHRgAB+YY4xzBYv
ChFVzRem2rlrA2vwwZj8D6traLfivEwPfkhfVC18D7rbYkmkAFYWnA3zbLwYW/XpSby+1pN4T0Hc
ipjntEeXulE4A5MMvxorzZnnLOKd3fJAx8DLrmiiES3XVG5aSapIczHx3lJ4Bo5196VJtDpjZuDR
+58ubwyX7UZecjjUo9sox88zeSKSW6CgNyrt+iVLQBZ+aGyfeN3KA1gjXY7T+VanpWEgzZsi9Efp
8aFbkiNMo3i0qYVw/TNMT2ZW1PDaKgALyT2WSg4NGA0zmxZSaY+DwQsVhhJW93i6PLOI/IKRll3E
g1h/P5PwYcMVYNGxmYjVAkAnKFKmcbqaO1CXaWGZH08+cQDapKmZ2VY3NMwgpTjcm6s8QHS+Rnsc
kBU0nu/d+ISRNykH2zfIm5Uvgpgk10mNyhb/xgL2uENPmv8aDQ7WOvXye17DZz3K8HU1zw1Pq/7R
QQvoyh7LHHF3Kf8t1rwpEhIdX6pdBdj3OWWj7Vrs+t3VIwX7MibSA7UTgJDEIJnPXicyhLLyyo8P
g1+hFO+iB7n6N3nVVgKbs8ZupjqqBTnQV5VbbDGqpHKMAzqdQt8MsydNoFotIaRmaJxLK5Bt4RK5
07WYMePlZNPHeM4WhwJcNoXLoMRXPQTlq6CJtrBaU/CgiMZwmomzujz0ikQOlL1fSIzHyf7os58m
VkeTYsDlWJUYcu9GNYjpd2VvskWukadR99PeMyAJiNCJ90oNLobCHsq1DtIKbyJp7zwTUCWojoeC
7H6u8KVMKYpWZOX+SmS39QlfNu/gpO7IkjnAiRU9pV22tUfArQVvNizBbIq6uMHlyha6kpQ+m/8v
Msbf+OxJkYvZFWtnX9dmq99smLU/kZ7aV7oQKIqxkEwaVHim5xnzVtuwTr6FshYCihh8v0/ALqyJ
BGmKsmaiVNINsbCkGGoOubLPxDFpMJltWowwmPlfVapyHOqc/Os9n418/jhm/pgsn4h0m/BqMsh7
6afg1ZTUAANmMr+ZktQYUCgweVqRTxioEunHAD+1ypFwaiS7Py5JTlySei/Fim8hKAzDUNxNXww6
6IQ2WN5LttICrN2GQGRbrDfKYvEWUL1gQEnCiO7evrodgpHakde+WkuTwSBD2VgHaBQpnfkqihHU
rahPnSQvsLgjX7lk+k7pbpr82EO7ZL5u8HRvy3vZTqmCQiPKG3IHPyhaavYVOM437yziW+/k8M/9
RTNioZMKw6AtFLjex5qLDlGoMy/Bs4XWGtDVAkLtujTMOmBfGQvSWJKtVfKg9sr6/ww8D/2o6qgD
3yfEMYnlqdPa9v25I1JZFgpJmF5750cJfraD0EzNAeF7AiqrV3MCJLE1zAWarTuR29MO85ur1BuX
/EPOZ031WaNl1bpKJbuMeN+EL9RerUoHG6yFW0RjBLgtD7zEY0qpKtQcUL9cGK9IkoqpPP4J9Qpt
zwsfzO4LUn5XGj7874dldhp3g0NvuD1GItVKi1kT1lVb1QUBr0ACB0d1UZ6mNeXnrGNC8fGp+th9
+nMUtD26LDWsKnNI/l5JeP3wkD8cLfPr9DIL0ECsAaYOkC7ZsHqVh2GWyiR6K4gtHZzrH35NpDD0
aJHiGpChuRYxdZefWwfY9bujR1Io3sNFVD2vCV2U23HbbNRoSMQPOHPM1D95Zx2g9sHGS858hpva
uLbyUbe1Fux+DN2YYQCNtj2sl6RSTt57Z9WnJREZq79z/BvWvJCYCam9dXKE57ppwlDkXL8nGPvC
XS+30eC+ef5vQez2G8iuIAMQN7u4njSe/uFslokQEQACmWlOrY+3Yw8VDMMJNsWPvNdW8V/mSKKi
8sGt/n0G/f80kpa7uSBeJuOFxuAs46GN5HmOolas1WbKSQ4OjjqQ5NmRIkvNyQneRdwSXjnIN37n
gA2X8ve38DyNMN3A1uB+J7t+J1XlbZgyTWUdrOZ7SWiX2nuA+lG1qv4tw9bwM4zE2I/L3aAzyey/
/ux0gP/KYuisrQpeA5LBWbxu/2YwkK86B3xmfi33mo93kWhkPyIul5RkeLKNgqp+Ox4W0S8V+Xz+
XC4dyHftrTu2GZhKUA9XnU3Z+jIvLyEAQq8cWxA0h+AMALB5BY9RSL9kZN+sfsy1R8i4fWftRdj+
45Nc1b8igbLZ9iMAIVlhZGYetw+Hq1y1HrPoDjY9FMddcey9dcjCXIpFBUneeX3opEiOD38ta18y
FHbH05mWsPqpSjSkz/j1l0w8fkzfGhOQglIvEhfjBFCtXoO0gHiPkHyoep8fJ++xDBe4AdLPsuQM
ysT9/ukuO98+5ZuO1CeFZe9jOFjDAm8rt41/xoo9o8PJnIkSx8ciiAXow5kgRlzaQTpwUTvJICu4
wh4GGDLMXNtSxzmrDrRH3UYNo1KawYAlT0jSAAuQtmVX7k5l8rxx2w4ky+ekOavdoYqvpVKBz1pk
2B+z8ghaCvOP1OJZYHXNB6cPcB4lmA90fvI0EtF8yDIpfangjfvWtJ/ozq61Vo/3FQGELsT2hCOf
GQFsq3hwOT/9vbCOrk7QhPf1bD22PBCDvtpQeDMoOXQAuhHA/jp/LM+qEIFd7svdF/3ziQ0MBGQs
aejuRvqcX/puUc4Q4eOYkgInS2CQfVS9pK7DNKoBnM5yiTP57wNoVnxcbmlvl1YOcg+4w0wUmX/D
Pi+UcbPUwm3hp/Ov88VaCmZm+na47wtoyTfACG+Txm3+7110zOet1awHLcubMrQosPrbHhhJ8pyv
fhy5JHWXqXYCrypYSjU6aZtc0WbFGUs/uDYboHoUHeIHpzKKmZLiZeYC+49hA/LdG1Kd+Hk+UEPs
7+YF/itY2qpEz3D73YMFtc/qGig0jOwpaWmPbNhMIz+felws5jxnyOBO5auVEUVtfofK7VFtgxqZ
btbgytHNI3+cw2+SLvx/sH5u6jp08QASt8Rr+YoyKPop5aKhvZip/YEhYRPzWehQi9t2JoA9huDO
g6Ol3kzh9l8Sv36SKqyKeKKpKNLtSHYSeF3YyJ6HNzLbXpZKggAu5QPKMERs9kGajAkt/QxLDr/5
7LaE/FXfQBwR7A+Qm9FILbn7AeuXboIk2sb0b22wHaZtu+o36RVjpzmEpWMUGzqk6LYKrNPNR4Yw
EIBAtRMxGuz9Dt0NlsxJ7RjraHiEaAUp918qmQTwF0vXOHw38Q9WRPch6if5XeSJ2N8bUjiB1AL6
RU6ttGdJSIEKAMDJi6ME2eTSZ4A/eJd6wT0GR7YhKIwGoSrnuGdkixsXMLrgI9IadTtzpFsNydyq
5jrge2NSei+aXg5Qrd9dk0Gs1LGz15YuZWStL/q25OWy4zOWla/KtK+ZfbdaTZSZL/NqqQ3kXIdd
2R4zOKVVCX0KQVktiyY+ZMkxs+M1treKi+pS4++fEt+eUNdJ24zGlFdENB88As3wKqYzWccLg+5u
em0gxBS18A3todOvh9ykWxWMdPoGxS+Mt6rvCgyJkzA+enue05YRcp/Xz6PhNZzXiw8GfuWAni+j
8xmvL/thQKMP15Od0v0+Z6LesdxvU05JBwDiwPMlm99+Ngth8Rpw4G2g9d1gxZQOG/Z7b/tiSfB8
CUtBZc7GvpHPkwTx23sg3YEgPUVv65sWUllVrfoQoErT2fTc9oMu68aOy/uEwsMfEhT7Y4PqZID+
OnlFEvheUoOk3A/swNxmSe7RhlfD4XT5CFBmgTXx+jEYMez5aSM8/Oq+YO7lbluRNGVbBTaX5Duo
T6gQSqIitERcxpjr2KAyxkvQOqrjMoCurbJ3cM19zEi54NJ98Mx47R6i9DY9yBdvhhVKb3IJ2sV7
2mTYV0VHdt3HfnVSUJSKiqfICs2YynLYCGJIOpmP1F1ToQaGsNtnVA4h5vTcC7VOjkNVe6yvov7I
YtwBY7mq7vdJypECwXxMtf1KKXMLqTWBue1MrrmqxuPn79Ftj4SGnBwufI3hPhKv76mvuQo3Sg1O
HtsamVUDB2Pp05c1AU/8NQv9oYc1ebwhlI7DQ3rx6W83VBBu9RwEPUobO4vVx3yZqt2fW6C+Xm54
0rgyX/+XUyMnIFBaDr1ugaJBhYsrn3JpDLYmRhx0oA21wEfig+GFx9aVqn8ki2nKwCXO/Ysi6jji
OJ4s7WHQtti6kCxMl7shkQClW3+Qd8xQkaIxiZiVC+WBeV8x7pmhNpwcMXBfRnLIdizk7G2y5xQK
2ezVqwTML6T/QEkznmRyIvJQOUJCAzcEbqhy32cLEFmrfqSnSZTKn624SMlUpG+wcGukotelBPGy
qZdbl0dzIHBLveMIouDBzbKNaxeKEvUasqynTjCUrS0gC7IyPm2LRaH6Vb/p2jGlKsgZV9iACKAG
sqwvNwlxjxCrqQLUAskz9JQYPldQyAd3fZ4R8asbRLZRN7ueYv5T9KUVCzM+qc5uaBHP1E/oeGJx
XwfGoTvMWgMMg80JUjfrQimOQw65Wvkh5KQFR+lGQp7DFjkcitjr9/Jf3DGRvnC+VC8dyCG6Thmg
uJccgb80pdfG3Hy/E6DG6MCqGXakpGzMjWiFzyajubrR0rCNUzn9XVd4MkfSigq/z+N8J0RPmocS
eHW15epEc0cYs8afyalwYoeiYZ215s0UympCQJ9Hbv0n2NonbTJyeHhbZmme71+UJPc0h4WEwV50
raVyRbD+X1TAPnlnQsSsYv2EM3lhJNvhd1DXg5gNSQ7VMHv/oG/Dj2AWVN8YHtUR8vBh+VnVQU2K
hcr3TMnau9Hr67pCnocOYLymR2lnhu33QbwR++Ftska5gkJAeqpoXz5rdgJy3zCgKJtJb2Sg7YD9
eeR0+mHgYPN5oyiKxNsam96L8QZAVA1CDCiLPKVArCTLv7DLXnbFk4zwm3zwzyCNDC4VS3kYh/7H
C6ahCytP0Dj0B3XkCXMl0LfEu2a5fUy6Q4chTWzUByrt7Q7NG5VCcarbNF3RAKAdOzU8OYnGaX4D
EPnjBQSaNMJhU9K2OudR6N4acBgqJCcoAD0C8DjV7ITxcbCpc+9e1l2i3UKyaFWslHJ8RpAoBN56
ay22smbTJGStukZB54Ku+cLCkzkJmWeQxDY7huIV/oGSZbLrukKPMZxbaNVHh31pKJMcMPsVNuo3
iK+oLRVIWtE/5WQE5s3HL/QKuJnaSmohe4a5wj4qNgvb4DFDkXAjRTmuu5Fllrj7HH9lEDbGQ591
GNSf7cQ5Sn/6hPeIY921w/y/K+5ZqPGeYMxGs1iyLpAcM8+RpUFlN2sTvCw++43FH6dESDd/2hm1
k2tgbEP/NUGMfGu0+dY70g1KYpa6xjk36OCDBABn86CfnjIn6WHj8S8yRpkVxFgAhETmhGPNuhrG
mcsdC0h77TrKcnVVv0mcmKsDI/9OprrCCSQUehK8AEyQkXJK6jQLV1GtZO9ZSrTyMjWekkZ8CgZB
g2CMB1CbbLl8oPf+Jkl4pmkL0xyItGJsPWM0AYg3nFiuET/sryo7Z+R4UospmLtaSaMFPRaAm8Rh
CbGM5B9W5yX2WcCW3RrsBTlcLwJlMzUAxME4zFxkD+6PYPiUXU9HSreSkCGRUwyV++4m0IsjZkWS
ZNXw0z4HqJPwQzbuAOM/R6YjUx50RMlwZh7qr19ooS0J4ED3GJiqQXF0JpFl8qzY0HlhTpRqeFEW
2F3xiAJvTzUzN10mHgssfd+FaeXHn6zH/dmE9B905qnLCNdgRySSpY/Vk6HJyKhwAT0vYPFbU1oK
nQHUVumMmhwQJnV+woBpglK73EaLJaPgw/k5aKaC2BNC9KTqYti0F75Cv04PkMAr2owMROHosvC4
25belW/viXs/dUWzYQDReeICOvep+X2OQOmQXGh1I4ve6uNQKzCcQX6tBhEQ5XcN3NquVn3yobDU
QKApB0ikpeneaPJCZqTs5oxMp1XqJoX/4qw5xgfKbJ5H/pvCmyuLCLTXvzjOn/2ro3FAKJe0OlEL
oAxHEN5hf1VVwJX+vynN+eNtgqJr8KVMj1EG45E8ioil+pI4OzBtpB0UFN+IGUuJGK0iyn+BA3J3
TSXSkmlGLwtjIb90tgCbvyC1bXFYRke5gsuO+sYeEbmaR3YI0BA3k/CSU2SxdZNYbQrbws1OptAJ
k1W2ap9VhMUMbJGlltEjCxPZrn6YfNGtjcIx3pk2c6sfmR3LonhRiLBWMo2HsLtv+ZJulRqPcnsO
e3qdT6vcunPrX1skMoN3ENcy1ulW/E4N3jKIeRLKoGqYifjZ9SsKQXWMoGEQBZr6SXCceQdUb9Md
TlDc2N+9OtxH+aAfd4ZtYuFUBqFTI9vfBAb+zr41o8EnktUS20A4zOwH+dqP50dFycMGbXkjMPls
PxR1dD3kZIKLXoz7oppzxaZQTBikGPXK/2q9UkuQu0DTfcG6thqj7PUsGKBwlWt7AIw5aqmzbEzt
KqVJ3jCfLDyY3iKKau4L08ERjTw7QobENyvvQD4qIMja3A3e25UF1bPNAKtL2aUrrHzhztPDMmW6
j/3D7DLPRFdr3xUrIwaLjw9ma+FmZuzplkX5zp0rhHeg4J/2Pg4fCLccDuxFE6dY7jZLk4adj4gk
gZE8i+yE2KP26RaH0+8ER1XzcHmpHoyMF+s1+HGsnsywuQqTqdHcliX2ssa1mDWLyMQlanCp2Os0
qsOOb1ydRJlwd8LtDtXLXakMHtPXRd67IQlis/gWXbSRRw2pbagimFEJKRlAQJYW9aFFZlBqNFBD
3/FQuCtD4gXysjzeOdXgThcSXFpsOO4SikXPgJ/isVyyrOPTHlQAO7Y+u5oyyBRMxmyDJtQRgpMF
19FHEMQ4g6Fl7fZwvqGqT0gVV0BFUhb2836vuvop7gm0fuqfzJd+4ajg8uQDYF6RcrMyfczpSq5c
CEgnT6D/ZWXhX6A0UFrSSL06Ht0qjYqatcVnV6gGhbdEa/9XOLbG2QzHUv/QmiZyCV+kgkF3tPx9
ZzdS6c4XN/UVzkItSt1sbnYUxncVRbksoGiv4N4R3wgen3oYBCeMrsQdpiLo9hZDQFNjQUal5VcJ
hiQ1vnbNNxngxsL0uB8gaSQXZaPov6o19a6WYXmRQzU5n4qgw1Ls6MFgyqBbCdO0QCT9KSzha6Iy
Wc7dMFydlUfZqg5Ms4cg0RWJ++57s6/4shybQhIUNF0lVcZpAPTs7I4UXbsKswzII9NQ9UZ1LWs0
FpWmE5WNhwNOJfhAqfxGtwNBexVH755jCDspYRWGMADKHlHL3naSXf5SqCqD5GyU2A58s0VAgmeO
akQCnUmaqnJkKEVKW2yoFh9Cx/yhwwsXJjXLnUl1fkZigvcSFXZg0+1/Yu8DNvzhHMT7lsDRvF4h
oT0J7tLdHUAwI10Xust0j9xwHtDa0aIZ2PRU819ENpwObVb4gVxH56LfrUNVkjNax88ZDSas4uwm
8JSTXEeHbOWEBeCAnCDHINM0dmhxFs65fzBpwE8/YAY7BhQDkaz9SNY7WFqqO6rsg1GOtlR+xjU0
l5cupiyg13To/3wGpc4YY07+oxdD0pqlm4ARX0blB/O3gPrLmjKwOBDZlaWzV0nQtUmv5WnZgb1l
7HktTwwG0VQJVHPc9XPp+ZRMF/CfG82lU0Y426aKIvMKLT+oTZT0bXWPjh423lDuS4ZFSHlxS8GN
GyP4OxI6HcPQe2jQE++/oHEnPDbkp93TB6s0qIPX7xRnH5ETwhdK2JJMH92xki5N0WpYvBgwQ2sr
xsSUlJYVqW39I/pvJINGUQNTFeJcsES4AnztF2FWZ86XygpgmpcltuvNGuOlZhcKaURiup+EAEEv
j+akDbOgVH+0GlzTUV5A1OnATE8GvU1RvMhBUXfydlxgwLmsRwC3+w0G7/Td1lChAbf0U4VVDrI0
dH8dCo8hLEoMBJuHaEOH+wICsBpyYOiyMIAFMpdCZ4qEo/GkOxo/oOPbPdzCxllUHmuRoQF8Ah/L
otvwsSKGWVHp/ALO7yERQz9U/tD43TrGfc7Kk0NdZM8tQKBk2LyGY0kCewmJwZkZsjmWNNcWUkp8
yk/LEDFFQisCuY+vkTeQoPGfjhC9G0MeWtqBPDE51g3bvABlkm+Nx7IOSWnSeRa/bFFMwHNj1iWn
bQsH32QHeb/wWi8IITu10fOgBOXilNpAGnkAtI5WhWxavY03C+1zW4l1oGjYlZNKYG1C1ItIRoni
rPrShTiDnrg+NGR1oYCTGATEvs1Gz5H0tRPhWEwhimMF/9+Lbsd8jJuab8b9Pxm9GhQ2DnqbkECD
gXHAc+24gh4eJOie03YFavUHv4WJI6b9zzDSMHEAiMYY7qax+4FM2A+Hlnd7sy9S1tthxCY2lUiH
G3QagzzfNdaGfLEmgX38glejOZ+VnEuQeEoUodJvAZZR5Bv7URtuxLmvPK58+VptMglB4dkDsLme
1gygE1u4TYJRcSy8k6qaBrST1zwN+deod5mmR1lmWzwNiMxRXm1CJUK9uVrzOTdnXeOdgTYFx78r
PbR60R3FVhfTVUGDKhxKu9TCuBUix27Brf3+cZ+BSqg66+JEFfw3dVBg3++TRfvlknLOv3Cis/zT
LWFaQB0BWTY2CD++NQf24W6QARvdTkEvqyNE2NBbsJIoa0tKZ9YTrVw4uboblg5Lc4KxYfjC5em/
xT5eof9W/59bwwIJJNCRtuofPq7W5GgRTDaV/RPu8q8O/VaNIOWg41RfHiBlO9K1+647/R8ZZ32x
mkfoOH11VGfHAANTS/3cxbzCSoB3WphTpo76s82xdj+39wYRKBCinQpNNFoNpKrUw988+6wLdON1
havvQbSjY06+kxQN8oaOFSbx2N7ZW/ijin0mXGJXqi4H82j971QYcK0F822/UwHhdDkeCf/aZziO
IjkWg5wqmPyzRNgFWTVRn5fMM545wu2u1FK48b0LpkmUQW1LoOdbwLmVEOlAr9haW7K0MdyUZuzg
Tjs7kGyqQUEqhak8ipZjGVnlbQKF+Zo0oGYteP2PetxI6/8x/q+1+nGOxl+ilu61WJWbYYA7mW2g
fu7ghcaOVyMhNbvXT1fK2ZnmoYQP9XIsalbiLJGRH6joTFFzrCBh5KQiqGbFU0uoCH9aTZKAGqfH
x05nFbjHFlJ7jPQdCmRHG0zCzTn4jKeYtzUBVS7W8Qkk8ZMsxYPsRgG9vVbIZicAEdg1GHYounFG
nlMY/ODFrRHVGQW3qJCBt5Ihea0qAscFC5ybUDBJiLOcXO4OFwGQ2cIirAdr8cBYXgZ0/RH6xGTr
gDyqDWue5e3fLR7n7NUOSWcRx5O4tChwaS2wE+monvjXrdlwCABuFxjLNdXgHFEe19OyvIEm7Aj3
lkenHSMr7N99FC1ZLTAiUTdzwVJVJQ6PDA99b7QDlQKYS7defM3jwU6hguLbn6vGeTZYjzbvshix
SiO3XbeCuh10nT5K4g2ebieJ+8eBOn765IEXdXiHeGLBezRToGqkiYEthxCnJYczx258l6YONHLI
nDbqOpcnhYXXS89pBoBF31uThdBlgsOqTfys5tyZAvC6dG5AmGmdorH1DyESDF7ld/u1/1267bnj
fHbKBBf0xLwJR/14m2l3XUn2l3dJfqJVWIMmDFlwihXyO2yyUzg4me+h3+pbKkp+23iNNFETz4RV
lATIXGugXEdp1YY6DcEKtsQexXE7ckPCsZKBIzzcGrHEI6Oj9JygB8h5a7MCmyH2A5daZU90iVRw
P+0BdSRMqWp6hyOOJO07fqyKAH5YO8QIe9erdqzwKu24ogkrJ1QUFha0cEJTMBMzuZODeTRrgByR
hIawakxAhNFZf6nXOKolvU9+bMqM8xOlB5izHNdG1v19S8hpDYQ3ItWLtJvmMR/qKzNWLhsmJniN
4uwP0tdFQZ9UghAx93zI16QYfgInt/uR5mmvbIamRCNJCPE5ni09cCEmMcs9nzUOEcCq+o2kQmjR
fvOF2myhLmYpn2hXgb1GAHJQPh0gaznkiTSDDcG1U3p9u6YlKUitCLC8xFxJCBYt26LDTUsoqgEi
Dq6XtZjfhcGbFbbd1cORmtPej91k6WDp9w7hfwlML1Tqvhp5R32Wx6bLOE8Nsu/Et6KVzyXUBAMv
2gNxLwkWoBL3o7T+CqWr/SMVeDLD0k3Omvo7yA9TJup8VsSTKKLBBYSnLwSZD9vVRr2ekL54/wsh
sBOSI6omALYYY2tcYIhbYFyWwlO76+T4U8ZuiLShJhgNU+S0IAerdJsFbnm0KW3LbevB31qujhqo
c7yy238qmYKfoKwz4qIJwIgBcSKJikxnAMB19vnREAs21UGxLmG0UYLNO6YeDZwCrSWjV6EB9AOt
BAPtZHr/7TRume1iwp8XHuLnwsiuYbPDddobrfEN3tQYABUaRT35ZQkxP5Sj3b16oQsAQ1c8rw4V
p5gw8zbIU560J/Bi2aLZKGEBSdjHlnQypdjDMkCiLgYvnbTtDAJsHUOlXbCHvaNTPL8eXOVUysCv
2oc/MMWYtvkQc04zhiA8xXQVADsquNWmg6GPw/tOZuzKVTn3jT7lxjdtIHz4iC/J2U7L0/89RmhP
tdVNHwFXIIaVLDcOPSdj8jsTdGg48B3cO16eEGmkuHu9VRxYS4Pk1ejJXuqaWUs0lUYYlX5uuxQ5
Pk2DFRtqfraFZEv7qvvSFFcH18j57H/noSK7Zi6yHbN7niAhgOP6sOR3eP7ECYLmmWtD9RXLCBhl
Z2oZWbZtDFAw6mATFq3NJJzEioH552PT/oUdTalGlI0euoO9I3PuYAuNgknO0KstJH/9YipqLunW
9lmBnS2EcaRfDt4I04OP8zv8p4c51HH5PrmjZ/JvWPamV9yWOVOtCbAXfxqspR0aYfnoh+5ZViws
VplJjzOx32DBF1ZNsRQWFcMT0NjahPZYK5UhPESD4GwchVUWhd6uiGgFQnh3fTz92h2Wvd34VdUh
RRuc+SKosc9wWshRDJt0Al2kkZfmg+ZMBaZIkF4Ni5ZjFqH1mhz3mVpVQKb1B/XjbGZTBiONqP6C
Gy9nE60Ytrf3FvMN6PA6ABgEuxD+6BiQaB22I0FnNQdNkTDb8Oj6CGzU6MXhnfjZbzBZmN3NbFyD
M8GZu/z1o41gyqWdFBRGo19ZNC9J/NZclft7mL+VaZjh6Q9q+HsLAi/2VbQ7HzSt5VuoPbGzaddY
kib9k1EavD9CuBwpt0qFhraq+mzvZaZK3PLMLDTFarvcWyMSCkML+NirlLgNB7t1sKAp04pP31MZ
XdoMhgGXc1pw/LTI8BqYTlc/BmLrPCEdvC1qsB8WCPmnT4fEW9DbpNfpm/oDBwavf/q6lwca13Ax
WD9LLNufBh38zOyhKkC7hTc//ZZrciGQtc/P9c1FNzokbkORW4Co8zXw9qAhPsE2yriY23gkEhne
6AzQ+4czK7I/4MCa66JUiu2BDrT6h6/2sNp8mkGI5d4iHM0468xLLxWhFViFeb6biPPYzlgpbaxm
6m5usSaXxaJzbKgt48RMzill5hHqYIQ53rEdCYdKtXr1cMKX2bzX8h5Jg39/IDCmEC5D+WfX5dFG
sTQSGvTI55f6l+EoV6U6RVModnIOuBZrLSfdbCIb1eOFAMCUnltELmaSvDUkPuwlZ+bvqeRTnc6n
Db65a7+KwhmZdWVxEwoMBBd6Pt1bWIB3SkSmHEUS34wlhiyp8VNGvlOrpGbtnUWkEs5J+H2o6KaE
2yKfP6PbNonNzHgtNWf+5dA+kOGnds7kA3tNOKGNvWItyeo/PmtyzSQdgo08LuSutVU0GEgqD5+4
fhaNLCobl7iH5eCE4rAN1BQQxaXa0OG6J/4PY8Ubm+9+yV8TW3OwtfjoEiMpUOokNnWfSGa4Jl2X
L9vc3UcOZXCdu479Y3BJ1OVB3RO0RJfgVANpmbCsomX5l1CrZ6rSDmTL+Y9g2YsKdwJraS7Air4v
YqHsrbTlh7JeTbpv7+S+o7T6jZBdi2NEPDfEXKSG3Its+NxvADOn9zLJMUwZBvH4CKqFKsAsXiBy
SDCntw9TVBpFD069CIsb+Zj2/4TC8FpBIqgikc94/0PSEAS/wdUHkNgkwO4e5YBCbmE03ckGlcoH
dJ2FaVd98+TZVjKvNaNboc1gfHs5zI/0izXas21hYZ4IkAeoeK2DzXTat9DolEug+rbEs0zKp7Mv
87nRyuVquKs7bWJ2jDQnoRvKW9PqM1VCpBtx5tUpjnREBtT+NCp63Shpg4tNIouWCwxjAyzRLf3A
rxl/UrI+6cHAfK/C9SeBnuEeEN5MEl/20l5Xi0U7G/lVLQiB98amrphiSYUV5h39bvRPMGtFAMl7
+wD9PMwkD/A7gngAaTrG9poAV2qqow2ESvAZVIgmyWntjm8B0cstaQv3MAGr8bQC8BOvyD0Jmt+Z
J7ljAMRK2tXNDn9tC79WZHcE1hYvFyTGO29Sqhj3spaSQzLkdQ1ktUmg1VdHQMkrDvF51Vc96T21
dv1dB9en1S+1NWY4Gzl1Z0DCE4wXucfXEqMlpmmEDkLVLt9b3FuIPmuhcA1dzim9mccw1rD0+4Pu
x5N4z3ESCxZpggMn/vGiIyFGvRuJwnVt8ykqW0YVZKoUJiz3uAQbda1chTSLkL60auhQKGDTIlZu
SWwyJDoVeiwrXiJUeENyrFCTpZBgpQC/Lh/qsKmBm6lT++AYKLjiG8e5yX9uTaM18ht7nEbOMPHg
61Y8nONtRs1T0WrMdYotFfJb/uq7Qvk0BBOK8BUiAyJitCwD3NlNnp0Hc8ck85ETlvfUTfBa74Eh
da8KRSBBMTDsCO9n5KuC9huLL990zIOJTp2ipGX4Mu0RvuXRl4Twoxd7ivHpb5mqM5ufTVqeYPzN
Cz5pD8QHBJ/sR29bTX9QAA1tWtiA/hHLqUyf141UPmRSYrz7/Qc9I1qWGpb+vAlgnseTnqVgr5CF
fH2xQHNNHJgkVgRGkZ0gOcO/a4nv0kriOkO5Xm9evGu3jEIATTMfwRKk5BHdL4is8x1Rtx6+momf
eBddatMWfrrKQwmDynesom8HWFMYBiSjqo2VN/cBL9p+WF5thPEnHif87AfUTfvoLYR4xIUSojpP
70zqjeowKbGIdMsbA8h0QkhiI1mak6ju7rPw3ItHdsen/XyCNPRSdnKRmXdUoYuFA8rYXuUQ8Kke
GKl6ySy/R6JQkG51mKGtyJxH7b+LUSlwT4oUfod17J0SssE1Zhjl/0DZvRsYP/1H8o+8DL0rkWxG
vnttSr02Yb2ee5A0nNJecRz+YVImp+zvkq6QTTn8LY6FxTkWhhaFfqfsfYodbwgemPEzxxSKrzwQ
IePnuJCMaXXncZAXW0povHEmPiYxTU5Jjv5eoxzyujS7N1m6CxSTzrLAgwIWB8C0qUgXm3tsqLng
L7g2lBPIyUp5gZ4bmXxacY/uanUNfLSo1gBzJO0F63bnR/AJQIhLH3dekfDPa9k4Svl44VH/z5WY
37CEUG4z8PysAhYWId4KOnRSvvzCpndtD8tZMFzLyGKsQJSiOod4EsYE0xK7duqURdowY2Iu01rC
296YsWpG9oMaF+cbzOA++OC/WS1ykJk5ujRpioIx9m1kDjoc6WdQCSYlFCa6HIsDjMRtqUQ28FSU
BGbExWx2YiCWnJWfIuGledxz+vbccamIQFJHXnuuGviESN853DyktePCEb/kMPkcIYyX7SrRuwDT
Tr6Rub9MJZ8nOsoZgECY3lsrx6goYSC1yevRG2PfKsKFNANNG12fpuDx4jCEVTVEmrWrqwexEJB1
iPXmEBZtc7iBjuDdX9Lq5iDSes2esMNsctRKLIEKCWaXJCctR0NOX1KRCS6alotLB+zlD/ofSJ2v
T5511J2orP7h1QCFdD55COWj5WZ1Z/Su5M/MLrts+41k3i2QI/H+FgU+4SAq/03IZjeQZ1zg0URT
Qets88hxOmg6OE9bXSRtitBDqdl0YlZYqLaR8MCAoSpKSEqxO9wlsx+qwIVTUeUCkCdtBM68g7Md
ZSBCPwL850lAvMSbCcvAsldfdbwF8fmANu1Dp362o7KwVr4TAH0D/svaR8nWiX4N71gvDjqta0GZ
Jk+YSM65xcRAPeB1HjBZs5q2JAMMGfoBFGlX3AkMCdPWKw5Kx0PzF9DPYk2ZxECFu2EzOkQGt0rC
lYb5xjQIEgO6mP1ShC/fZrWxi6eBoc5HGK8VnrH3LgW3F+VfKmku0FMSBoi/hE8QwyEQLmyYMijI
8LLRj/mbpYm+h45yubJxJw03qVWeW2FNnDkkOmle6u34PImEcLPA/QPIxAbPwMXNShLrUNV23gv/
ECfDNuS1QA4MS4Enqncn49rAjykOb58Bdq5x2iNKNsALimS3zKFJ3YXXMQFwyRpLoB3b40Dy3oYJ
d2gU2dFMiYJ+kpkyVKSdkJYSviJ1BV4zrhGCupSy1klRb/LUCPdsHX+77GmFMIMieL96sEgud3t3
yEYeTdcpF+SdQY6QPqzuqAEiLZVKgdghIk4EsV+AQwjU/qKyk6oFvhC7tda60vIW0knhKki2enCm
o2UHFNe0L78fzNxFLfiOJdsCqa6wzOawjp0cYSdoXuibup84RzILWhM69gQEYnxKlrB6yZ7Mkrs0
rY+4yWzFQCMsmYF6ggMUOogNnhhj2O4yAV3z4oVckI4lgsL5qlBGYZn4BTS7Wd5NVBdFViNB97VC
jgnaxQiq5JsJQjtqDNjjfH/v3hH+XWGXIFpRE8snUFknz5i1MvcxSP6JaJGVwOB/zmA4EBZNkKza
PI1qWJ+XSfBBEQhGy345DHt+EIriq+Q6ZAtWHatnBMyXQqp1Hlmy3vSyrnFBnWsC05Q1JrFrj4Mu
5wq7iLbqfrHklDX1f4vB3H7URKcSxCr6UZLr+2j0FTDlDHqJsLRu0puKkRPX2hsZqwksus3kKErL
aImXMjbkJdqGkXWJGVvJ6E+eftlCr8DxglFnjlbVeVmePjkK3PUHp1fjBoV++btaiQoqNECLFE8x
InVj/Uz94y9ZLfes2eUg+JY5VQQ9xiDibIeob777eirfwNkvFwAChApgarwi+wVhFSityMgjgVh0
Sge99qKbuS9jw90OkSMIYYnB51buabsD1VNwNixwaKGoZcOt+6PJrnuftsXtHW+a/3X0xCUHqJ2z
38XKEqEwhMoXfEiNJPjTbch6AD+uGW8Yq0JxiwQ96Yj8JT4IY2Beg646jzXhsdzcWk4BAMAIt+kO
+iIeKOU5esTzhaQNUB26B6vBr70pqeCmw+6lYSazTk5QVpOpr45J2IiFQ77JzEFAGVPhAAHhIYxC
Kzl1TMjcM5zFEowEZ26GgMj8kDnVyKXcqpcJBptRlYmVHhpa4IsC1XNBUvpK4dx3Eq575ras8Mqr
UEBBITb2NjQu9FFt1/rVT8mMCJd0DSerGDxTwZmovkfluDKiQLsYsOeE+EniBftPYiQFXyeLv+iN
1apnbJ9i1TSF2ZYt4w6nmOuj56t+aHUU9Im6lrmBNJxn2r9BcsPzRte3pfk+nVBTOzT8cnVL2hb6
N0gun3XTkvaQT3VlfVa5JRUKcu4lqooyEuN/1Nr1pXlIvyzOYoFdSHsY58tlRgd8vPxsFgFmFxkE
OHnd+YAqOM9pB1Exx5PoZLYMWyTQ+NXg7/mBNyk6c3o+FCGLUrqyYylew+w1vQhzAkZcxyyEBVAX
vcNBg+XLlWJKRlbNdgj27tYvuGgun9A1kkZfM9LhWF71ecZQv+nCk8/gIpf7QjbiKEEeqSXVE4Ec
E8FweUxf4tqGdeDMlBzz8liAdOJDyHShSsCeFFz/k2Xv4Z1ulJwUQSKOLfvrc0Gv5nKHJnh+gd5M
vpoIyGmgRh5W7wi/+Y9IHVhY1CmSl1D57IYs6iIfWVt7NdMhGWprMCuK9brPS6iayPgU88poRgHj
QwCzTvY26qUol1KBUUm8dPVXVEaRpJnnRar1TD1eFk6d6oE7t+DmhXBQhPKP6CYzwOYPfQs6FYNd
+Pl1QLoA0gJknZZOyy7nfEkv1Xz1HqYau9VTTvXNOCa27PVDgA/VVdV+4Ly8mhrbt7CGLlDafZs7
mzUz2vo3ytNVyDNnkxTwWApuzmDLLJrkMN3u9RjyXfIwfETVybSPXCSbpvo6Ev0zR6B+3NkxGzGJ
visrCaW14PhuWA7nYUUitaz6/ExlmqOpwWfjlUMt+JaKEZ44npXLKLygzw6Ot/AympDVS2vhhmON
LPFbayEY24UXGXejEIB+Ws/SNPI26DJKO/vHmWjTTkH0Q/aTlXY+/djOBa8ciBnh/FAFtGPygCtc
fMoUMQJs6+y/O46Ov+7qc3he4M4mx8iKGAPukFRXjRXOklczHCq20tZcyZKIiPRhGeOuyKSHizfL
lIJpVEc3W/qYv99GeuNZzh+H2lH5o25gEJVA0sYqyzN4pDUkIazqvBNAP+TMk7/0KSTYPnPc9qOS
orETzZpJ0ADSRKWltNLPBYulcv/UZS8RuMT4DJGc3Pi3BD8IGBTfd60JJPQFHtzyx5rm5laSV/Gh
xCQFY98b8KUzaXSdLglBGC1uO087rbAd0FizJmfurnm+ITQOv62+bZlnmmfAtBGrfvQSe7lq21T6
cZo6aHsQC+Au7I5kC5gZXP76Ggb3V+oq075aTjvqbQf9kudR4tzXrgql8sptJFfc2SgeXeMg1uVz
Qeghi5SfsLYrm+dZyheh7OGlnlr+SUdychmkwOSC3SyBE33tJJ4/Ax54syfOkHW83uUXhjAWCXmO
XKHu2k7uGe0naQtubdezJHt0yZE/htC1owd6fg0CjioU6intTw/ktxod6UodQFH71lYKKjq6DbC0
1lfcZZq2cx1LmiaRJyp7lM9chwnaWGHmPGkr8eAtwZA/QLMwtFtZI2Xz65cEoVN2K7HLf9QAFS/w
DZSFRCnDojCtiZkT2iu96F/0CfYKzhBTYI9TDhhj6ItgHHsGLIHcz//yg/947fqNG8OLrPGxTnEB
c3MKVTvLSyq4g8cGyr+ZDbC5B+24vXTCOU5Rw2UH5yi42K65SwdNj7pF89n7znNftC/8oCWkNuFq
2FUPFbCDYNjfPSHeTIvF846KWi5vCnkvyX9ns4+LuAUQfUIHSxXJ1iUfmdjABys/ig0+xjkDbKuF
atB47D+/4zkXuvpCadRSMFstv+Jd4Qon0ZXU3cz0rms5sNvqpntOEijP2IGYoXzWhaAQ1KVPGI56
m18cKXoOs/LHAg97jNiC4jRSimPaYM2hxfekrHKMLYI5lg9iZU+cROTtq+07eGByOx7XFQB2Wwt6
BQsN2U2s/WZUPTBY9yWo/8ChEJ1JGDtFrDnTM2n9j97UBYbzgscmZxbmqQTZILq1D70b4s3nXabd
JLok7ivJjB6MYDyJ/BTQfxm1kvd5xRKAKzD5r040gbTVvG8jRjUxYCUye1HUbkfjf003izSovqiK
4OsTRyPFPaBCU9hwSxJYLm8sW6DdG0zz5YhtnKAtAetHwSCFWYsZT0OrnlzCiXwMdRa7CUnvU5Hp
/D7gDiDutCO5Fgk6GjRtGdEp6JhA2WJXh/uL2pd1neBM1WwB01yzYMDWKf7XK4AxrZtn+bXs48ak
NyvWBrxD9QkkfVYxCRIxdXU8wrgGmCDPu9oYvtnX71bGlZCl6usWU75u63h04vzZEQqmQ0Iz1wTA
2PJtoyF8V//6dLOeQhKKe78yAAknfO0F1Otalgt1Ph7BwAqPYTOrknQlFin+4ufAU3Vyoo5zN8ia
k5R0Wr8CK0uIqQ3NG1ec3iBBLDJhf/MKgu1pJaM9aFwpVVvROceTAiHxyWZwUPJfg23rrt1R8QqO
0EPO2F20R1X36tQGkf1kRjc1oLWczjkvrdvvH4f6dxvK2tFZC55Z4zgjCakLHaC1Obezs8f5E8ev
iCFerukRwEWCwi7XLzOgi9/eCMb05f99o7vUB/mxHUbqzNrdGbtga/C3ujMtiNJobtrvpCDAOhm/
r/4zkT2QYzW0s98NSd+c90fXAPkQ7iLn6t9KLwIGCVKSfa53RLyX15zjnjMt6gsbkMAkGa0sRiwT
Epm8keriIkUlWD4tzK6JjZrKwkeJtWCXXx7Ytu9/Dfpur2zvwm/JoTePljLbgd5jZj88HpzNJ8WZ
eg/xrbj3mfls4YNBN1aAmbqdu3POpvPfo+sdgQJvwFeeY1WTlF9YCaTilkEnQop48mrxfogiqVS5
9KIWuDrXsyFBYl8jCpUD7XrfS7QIA/NvKzFO0cBQoc+hGS7lKmnjIfr7jTJDtv8H7Uz2BkDKS4SC
muuhQPcJRmte6Ua6HTdzo9T3txKVGfpigcvVc/Q8DTo5D6G6PXbp+z8etQ0uU7gFcWD8Kd7Q/8Lc
TEA1f3DOfSXgdYdyqKUb7/pQPu7XnYG2kqHAT6xQfdZFFYWJoKSxGqwbCp4q+NPQfCcVX2wZm100
4L578siH+SKbXIaEIDBt/KibdeS7LDW/FEMH8349z2BsxIhFYZX3QYuyLBZ/Cb0oBWP7q4haVp2S
nd+x+HGqLtU926WIQFaaScc+AyrPCzO03gxCG+0w4VBc3mkDGb3CXxDe+l71Gd4u4R5EiEQCSUUd
tbV6YdAavfVXe/9vNfvLbTe3u72gbGsuxkGxt2M4TZ/+xB7T0rGNMMmoDbDw5WLP6k1QHN1Z7MKh
SKltKE9cEQqSVgMSVA2XpRyBMUJaFTxXLPZWXYZVVOSgnw4Bl2Oqkw90dEJEgztd60AQvSevzHOR
HoFCwqMbVHaSkiPlwruuWS8nYkWzNNoj4KRJ5wdSnw5eaxwemJ+WH0gqJu/Euv47l47zjguLUoZL
BZQqvmSUbfHl68tHSex95JTkVD78QZJLPiqL3+RZTXPWixNrGErmMJQbVBxhDaah+/J0YPPFw1m+
qiaNNIK7BBwEGtPx2inxZkhX5UevxlnEd64RM9Dv0gcXqDHxfChILLgL+2BOTW4Q8+0hZfNwO46W
2fg5xkS4wW/kYrzY813NgjvcKjNF8fRMwFj9xRCRxJpVmyCWIZvIbAafMQ1sqyXYzT6yfKblVaSu
2aTdZQxiEGg9TPBWgKxAWB/ZuRTu0X7Al4JZacHWdPRkYQeP2x4PFJTE/SZgVbVjvRhC9rmmv+iB
3/QlyZipHHPuTEUzFF3prxBRKRDwWzhR6E6pocVth6krlmXFbv271nLs4HPh1WCF3G0wHvYFQPWu
CdHNeTyFuaxa5feigW4FkafsPIr7RDpeoQH0jwpY1BUxEqw0lcofil5QcQJen0aKWHx23R4AY9xz
SZBsg+quorlklHpo587EccltQMf+Vq39MFk7vplqEQ6y8Hjr/WcPjet/xWtrwto5PjILEuDB37JX
ZQC6VhQzfL0WZPII1J71AJ0uWwOzFepjk/Zxay61CGWTWUY42N42qKPQ2wAMglLSnoGExaO7oVSz
2VAr0ogGy/wVBvd3ToBHsL29W0WmPuVpqQsWy3LazHHiVOrkjepUFr9JK7OncGeN5LxyAgbzq+iK
sLv9ukPA0c5cr4g9USlFZRAYLRhYiPvUZd3hFm+Ks2uXoGgGb4b9Ksvvx75E0mX5FdLYaS0PeRRq
3WBeClxHJaNsDwX4+kctm8/RTf8vdRx+x68CLCSUM4ukTnPqBbs9oLXoaxIomVotAvIU8B2pZSxE
tKGCWGRZUS9lGjn+Hjc97X0l8S8RUIljtNzZxL5f+/2jIx4Kzz0BVJzUgZ3bRyIM8rYQmO6PJzMg
UeDN0QudS9rg5ykUL0GfICWSbZLb/CUjGZBQSAngTGJfFvNzLsOOTHQsjTOZ2Gge1rgIWdleU+6M
2ykbhZdv12D33BfQdzGUAVQr2/5a3uZVkc16Eadq7y09qpskZHdlJR95G4eEcDkaAIpdto+Z5TXj
i4kLKYIjmdH2mdKl2W825WjTskJFaievWIVqCSQX8k7VX3HmLhtKaTX0Avv3iJIFwdXwtHbRoB3H
BM6UilXLhGtKfizZP157Vp/ZLZugaKYT+Eu1pjYtWqmmp/yZY00hdITUfXAS2Mj1Cl9ZuvIfD/qj
mq+e96oQ4KB6X4qnK31iVxhedTvqRxBlzNk/NV48ePEn9lzfoad+q9qVN+KJTH8bJ3HvtBL3NMqO
LulSrZSSl0eL09MHsRwxBE7ehyM/GJ50cavJb3ew1XGWRjXHYEwIVXDbiIyNMA2kGA0NrI70VHuY
mp00IyijtlXbSC782Gpge/7q5Rzs1348vsEH0NC0T4yZTsgn8YUgVOIXQykJPp3NBRSvFalEaUUO
58UYRSgL43mikmXKnHmpqGu7LBcyzRL01tv0dj7tHW/VZrLamcAwVXr+f/XUywPR64KBN6M2TDVT
po0muSf9wxtgspHtx2K+kXgj390qmHYCl36JQfPZxIYAWk2/82g/Yh0q2GEyUZrWWgw8vH1V5Syt
GRMZv0/Sn/2e0i5DtCk6UGw/N1RAz6tEmYmXHpgrEx1SyxvghBVc2ThiQW7ARXZC15dUbw7Z9I7o
JZAbkSAkFO3/vXHXJ3HhAh4v61LBnStf23V+fgS3OIgnUxLZhz+tii8mL7iJutvEHgjMbteT18JP
f8nbPujR1MzVF1YzHKY6mxMC7g/HE0KOR5KLsPa1/Om7e0syg8j4m85NRDKfxo2OPGlVHdBNzAqO
7CedJz0YYlHf4aNxjilTuvholWODMnYDcQ2N+y0zFFimY74Ru4/y0CCf7SNftPBoagg7KeyGOvph
L4n7hHsY3ROdS8RATctog0eziltuhd/O4XKXZceZ7BBa/vN3Lf4gUTeA2xWJwRCdFG02GYxvmTef
+ba/UYFFhF/uYV1iHy1MufEbg+zm8y1cJ7vK+tXEhrd3LBo0jwT70+lhvEdMyZzQbvulM7psSenC
TabpdPLOjp8EL9X0FgzwcKJe0UnSKxnJHRM3oj78YM1TtraijgtT9eWECScVDIEd535Ce2+eEUvx
SbnuK1oBqQJjyVm6zpBh9CvjQFKZEpUBN+LLo9ntr9+uFLm4SYC7nNuliqv7C27KQXbiFaRE70is
+DGKKvkS2VrH03rfna+Xry2ROxwSQowIhS84fFA+s4w4Xs6rjY3fWlPchcmPlqlscVGXYfuxz3E0
CkSI0KOet+QszBL4V/7Bj7kn85GYIc8rp+WjNM0Bgj92TC+Qj+7oa+CYXrcGEiX1rPabeB11iqkq
0g/jirw7jolaSbO/q5WRuRAt2QaUHgUUjoO+ZN3hPvMVTuwKhMAIMZvDcg86WUkBCZiqK6yLsfBr
Vc2jkPn32I/HkJJ6ZMEieSyhA1QmaiyZBIjoygR7jXmKeHtFlhhwildrmgIpUTQD88VQnIWTidVs
Z7Tj4amW8wRBkRuV2GOHdlzKv+AjnFk5JCJwrb+WBfDj/0cOhCa48RnSratDwVFO78mshhpxDk1A
tJNgYKqSieTje7pRiLbZnMwLPNCps75Zv4cCRZhAFu2JF0ZlMBfn/uNn6swIXZ+l4b+8TfmYRmbO
sbazj38nHp4FyThsWKa4KbD10GapM/axubqCZlceIYgee00NkAIc04RihrcEaJF40Tf+YkHI9kaT
J4Qwm7xGWRj8Ge9ESyKiDzHS3QqVCzcg2RRD0irR1aVfpRGJxelerWQx+/q4ukj/uc6nT4o7anDd
Z3PfhnVeAbBCF2QJxLUWV3/1tCl705qAuVt22TnxoI//DE8xMwDH1LMfShTXqqAc9lCNA71mLnEz
+olnbwAhj9U0p+AS33v+V7HkZSYUppSTq7fWpfIT9ax/M3WZf8YnOIHDTed3K9nqPkS5PL3IeXxK
9P+nnL5xQ3HK0SIPB8CYQ0z+NkptbYMVSqxzURq3lsGHJ3x+Vm3V82yrZg/UJSWjV4anNqhPGLER
CqomczbpzYxU8BLV+5aFAYg16Fnw7zGA6pVqU84z+B0k3bWzJjGdjmeihw9VRqlz81hlsGAZYJ/C
hUq606pbTmO53e0AsxdKCR2iB/uwoA1xGMHBjqWE2pprLptLvq6hjwPmtjgUAykggaXs6Pt6JT2o
W4lIr8JmmdhE4sW7FUIqLfwXm0v4ZTNhioCPPc0yzaucVJa49D80zQlQaNRxjYmgqlseGs4QeU7P
HrYAbz5pvNKSBM0p6DqEdalrbjBLxwdFsvWjNdq1xLGQR036Md8jbytsZQ0nJS5t80xG5C2HvIo5
JGnhWH6NSyUlvk2vTedkJbsTghAMvwmf6Kou+7dJTRHEw+D9IinXJn1m342SlNRTgr3BkBabiE74
J8daXRaoedTlLsyTAWB7fizuS81Aj2FmRhKN7274rRiQUYF+6ivIuckQKLWBZVmVTecQ1IZeCtqS
2Kein4KbUXt4Vk6qgpLGKYcVMpIcuoDfhWx9k4W9notiNJtNeQzqmCS1wCnjNcGwUkLONhD/BDJU
Fa/V4mdF9f7sz1KserjxIjbwGXeSn5ilPL9R+Ya0kRsBqTVFTVUH82OlWYjureoCTjjH1zGQMPfB
MEZtZdUTjtw5Qvd15vNDUnQCC0XPICnomgk7/S37mMgAdrbPZcmqi8ib9pccTBYvir7FNzPOJ4eG
8jmWJF+RzRL1E2QR1/JFumeUPOap9p3EkbO+ZWRXd4bxc/G/rwRJbPQLI8TVzYfXOrWUhgQCLvbm
MF7j7e8Gj1kOVtnrCRihydzkGMZwU7vAxL6tlOxAiKz6oUY0u7jB3Pg6jf3MugGd32Oj8xUTIRVO
baLAYiASgpLp0QynfriEPawixui+GORNCc13ujGZlTaInrZhQwJ2qn/cAz63n35qdujTnNzLbDDe
rvK0IJoLPgI1ZnxYsG04nawiAJZUeJWX7bxqStdG7oC7mTR+nIPF6nBKRqCJCbPoeYTdvNgLb21r
PlfM0Ha5FqdIShngQYxZo4BNI9m/Q4ZNP79s0vmKzWy627d1VXKdslR4fL/MzlQv6dkZ+pqvDZ/k
4POmRw3tWWEmxDuLMTYh9Kj1uML8Wprx99wvnkOnE0AZNZEm2HJesyKyQscwVSlpLJzivD5tNzvi
XNPa1HqOEE9xEJA6DWk8113iysiRWxFwYFPeZo91WTMWBqm8H+w90r/5jiMxpm5XFPRxzcoN09Dx
sxxX5MwzlPt6mmP7ohCRiX2DYqmzeSjXjjUgZj43NicqFB8j+FxngJNw4Sd+aOAPOGw/Fk7zX/KJ
uaUFyST6x+459btKio0127xPFWiArKbt0cn105f23qdTt8mXwqPfEUtbXjQWK2Sa+ENqRjDYxibk
b4DEtuEnm5G+Md1CcHoiWdAXZHetdEfWqyxo6HzaZXmepVihpLWdYM1GD2tKBlZPbkSAJezeAO5C
s1gahHu8gy3zq2LSyZSaS5oUZifkQ3ODTF4vXPMyIuXpSwo3HIWh68iwZrLglDgn+mr+md7Cq35i
35FrvTVuhXAnWJTTgsNaTMHlygte6hYH2yb3+zHk2kXTqY+T5DABWiMt8HdSGdBu3JJKMIkw3eO0
O+h/y4OPS5asPHHpJTYw8xw55W9+KR7i4G85JC7kBbJfPX+nPJ+jvJEQf0zESiUfV2RVeXbUkCMh
bUv9ZggfK5w+A/DyX/i1jmmjvL4IiHufElonIx2tbgo8agNcSie3s3+cu1QV5bV8Zgm/4uOOoRda
lFotIjiBnx5EIgzygzSdESVdrIa8JQwHZi8FDhyXJ7lo6MviYj1f3Qz9nl1zvEkj4wnbeJvCEcEh
c8vecl668/O+W+FJdTma6y09CncVIZyHZC54PHuIHOupgoMUg0bkffJ/6KnIaMoQRg0rWVgu1Avy
gLtoUgc2Gcn3U0Jylz4RySaFxkHaDRtqonj+sDfi6sigopY0wX8JhcLOtaUTdZgP7kABE7+mZl83
JfDbPtXawXd4WelJg6byXzUey69knd5G+O8Tfn6NIaMXm61Hkx6OOv6bdSGwmrU0F9Ur7r0td721
H8sFjlGHxgmqSFoIIhvSDGng/dNAdPOulxnH88lSK5XzJk4txtwi36p9ytzqq3yBGPRCormanwfE
4qCqSHYMOasMyyvoLMdqOqdduGlqPRtvTkQ2+LLEB3DyTvWIFFunxBJhCk7k4oJD5uiE2LroGnhK
Hffeq4VqchDust44fhefceJ9tqrO9bamR2FbL4xp36bx7eSOtjBWFwkRCq73o2j0vrXSgRzrY5Dq
DfBGb+34ooKlubDBMLgBxE793Ib8fNvv6QcxW0pBPndj6PYmCQQAFiKsCj9Lspmm5QiP+msDSZyZ
Pwti4OkY/KfUdJ1VJBRbMNb3hx+KMROeMYoAH/cQWqtwtgMsOufpn2DhjdBjwnqhun/VGDIZAMra
XWru2jLDlGrSZu/3KX6gmWO6R1dcUmtWiHVM7Hg6x5x/YQqWBiOAc+Huh3Q73/Oe4BDt+tZKs70P
CxVJ7SptlqXjiSJJmzu0GrGsXj5VbXPMxZKQq8zcoMK/iiRQxX+0a0VwGAsNonVwsPWHqUsmrV6A
S7AnxmIOU9mgQ1ZBYG+wvhzuzbhYSSfLI0h7QvBTFSrdhnRiX09sUWXXIIrr/DiEd+rwowdd+Oee
oxtun4VzhLsKGyaLavVqWtSLYhBVbJzmY6MvThcEoW3JhjBjJ3g2lvC9tEjOEQakBW8Jl3I3YCBN
OpLsnHJBNOWn5kAd0mU+xwsZqh4rzc6g/ca5KcC4UMe7c/YNHkvLUmrt5PkPllL9zPk1mChmmiGr
7MWlD96EmmAltmGgAcs8dHjn4b45r4MBoRAwnB/a2yNs1g+CnmdfgWrS3afMR3bK1hn45seSzZCt
rufaEhXCXfTQsUMdTGqtdFijIf89OsyiSTx+7kXG7/FLLZvQtqdUwkbSjhAr0UwtkbppAF5HFd10
QMSeGVkAtN0RTUirvRPBIh6B9Io/eqZSe+yTrLAnwOVTPaT1YfFYgBxWLdJqVDZi+GFGrCZF8LDb
U4wk3rVgtRKRrBYp1HRLRWUT2pe+KDoUJwNJEIMcZy37P/dojygU/Vop7zTWmIvgCLxtZTb562ue
59q2h0nBCOZLIg8tE2Us8hA1bjuPpdnuChZm32eRB5oCFDyzbHtFpJJNQlCpREOgaS7XWosFmV5i
xzsbEFKpnm+02OHqxNXgOZLzaQug1oOoM7omrO1yfI/kvxAngeIxTYLhLcZJ18u1b8a37FXbHvCT
jdxBCo+WXDW1i59Rj8xp6B4QNAg6RxQCNPa3s3b96ZgarDyTp9w6Kh2survIwYMh1/teeMSpcyto
rJb+R2RWFgNVzwHWyoihTRqiEBkDKNMvfk2bgev8UZHyj2L+sQGJKDm6p81ASC+e8fkudXMWkcIW
A4cLWk3A1zjbkNasFCqPiit9EE1Q+pZD1msY62bEon+wzJyXYSWx1UZ0YZeUL0dYoLtRJeQR/H57
LlyHqm72W1HN31kZDp+XyKbyiJ1e49WmT4jVbvaaVs+YSgWTK1CYIhDEa/NUo2TZdDoZInnTsw5U
/cjTvJhjzfEE0PYbrPPvDPPr45m5FO8+GLNLyXRCjtJbFo5M1epD3p8z56R9Oq3W13wL24vHPFkl
QkBJMqtg8ErGa/CgYFQ7ZfRy8QfVFGnAgveWYm4FsHhHUFW+Xy7/wqfUipsH/3j9ADN+9iF1hG/F
ybkObwLM291p1R88TqqPCGA08f/gd/OuQcKtNoeVqKjR2WdPpWxa/nnG5AcPQhX1tCmoaU06wq8c
QGU5TpfMD17bOsRXPcq3jhffsHJPMoRiRlJx4nbrPALOLtNSP8PhVFxKp1Zjfp6O2cfFLBfroMlh
c61DMY7gLLGWBgEjqZqfpuCNoZPkFEuJi6Abi0umIyPH92LPeHDIUrGzIaFDi1cMzjQoAlBB9zBE
B+e/s8BXAFKCFJiJFBSSJoYGQ0YhoZEw7xMMjSm/tlK8alqGWjQHKm1Z86DSJbPu4qiH9nmgUmIV
rjiLTOD8zSGw9kj4xuqQPMuhG7NR+oLpfH5i5vH3Dn1bWj9am1dP20yRESpzoR32dD5U8mQ9eHzd
NGni1dQ1Bc8ccU8pA4v/b9C8c88swz/es5H+lDqQOPYeWz+kA+CQhK5plBuRt/gSO6montFkA55b
d55dgzV0F8lDw8FINo+v++MJoecPx54FB17a/2vMvyW6ozTy241f0vZYc6ujc1+yMGzWgV2aPa5a
HrYhWLqERCZ/79cvcK9vgum1Zyv0cJ+FrJef9D3QkMPqTk5NUFO4aQDH/BDGYAqzSmDdLWBeoWk/
A4YM5suseWWSFGKMtOMH+QenI6+0Wj5YN40hkcanBhhxE5K5lc+aoQkGGVsUCS8R9CncnOxwQ6Ye
cBkQeSDNRtZtiw4DgHwPDwiA+VgCt8TowO8BcP70UICYnJjtdWxlWTHuLCCXtmV2Y0Ke+jBv8u8w
d9UY9E3B/rRZDpQXef8twjqFAFZ4Uf4aLSqo1fkVdwzewY14/A53zvyv6JOY+raI2PRwBhD4/ezd
ENyROHHG7fuUI9VeY6NuhDFwtLyXwdYHQSuPwQHJoNhbQPbWOiP+tmyz9T6SkxNEVk6GMAo2URiH
YRCyPBEg8lFhuUL0zWRaSKn0MoVeC+Kcwg4IMyE3buLhT7/9AJTRvgfsL7coPHoMcpZWJhdyvRUg
gx23sUAVrqht3yePEd0U3GHwDEGsS3AQWk9oGCxZAU0t+keMx0yX1DDZOEDc94SOjWbvji+Fi+cQ
8ojc1WKAH62kdoV/miiCi1uLU5L6d9fzXyZIh07lLEwIDFhCvpY166NN94PEPfyW9YjNOdKlWTmR
/5BcXxRNtHpB2PG7XWWEodufEMNVK7j9TXqPx68iz45Usm59As2F5nkeTLRBMlnvsnWkkvZVJymY
Vq8v0AMn4aM8/YxCO7+c2HhDMn3H+KC1hYHvI8+gj4NIryLViFL966FAfdkaCCq+HAto3UHFBDTp
+pD79r6zOKcdiUJb9AOkD2W5xmEcXB0u0uP2jF5gz0WJbhpefiUSgT54rduM0MCXufzSLKHAgj14
ljLkdEnJgF+z7u/exB0RKF3O49qQbxvqQ1iYnLGaj6OaKzqh11ktHIKtgWFcKv2dVNYcO29wz9TF
EDyULAWlf6Jk37hJItQWTA8TI6ks2X9SjjrOEid8AMeobJYqRUu0JI6BmbSn+eKS9cciNzT0hY2A
b71T8AqMC3MdAJGsu4dZ+r+2edDWJT9ssX9dOszieRlCkJMoxg2v/uWl8n8LZEkq4FFvCRkwrV3+
oIPwAKg85JeKs/jsNRPy7t0pjkKBophpWV+aUZRO2zHyqNN/5AKLyjVpwv4gNtZP5a2BG5a17Jxm
Qj/Bc0wKMaLc/dnb+bLQ1KjWy+la0Wf9wCxQRAthWlfKcwOf/I1veISyzbqXNgin+KgSXUgmuqKE
B3USAWGvrnCvknF/ta/8p5aKJuZYoQRjwjegSSgxQ/8qbVMWKV9R5T+b4bDZVEM7qndMCzJLaiO7
7/7UXdyErUd7KKo+7WDLXfHpzQ9l5tag8Kg8dYrqZMIY9DWpXt+3iV+WcHG7kfYpJsLBKDJU47+Y
QqMUJJz7NjKDGsbgnDvqA3o8snUUgpMIwvLrYXPJZ+5QEpRCjdOvDY9plyN80iI8+GOWwjvMQW2f
BIV4sS3iVviva3uKjLzTtv/Re16IU9WjBwvRtO6XGBoyIhZc4u7qrTJO9g2LkHByWryn9Jq3VL66
OugQbkpuFWNmpqI3Ya5NYr2Bs6aB6rE80Oexv4P5wMmLxCZbiD+8eHQ2X8wWTY2VP/70FkyePyb/
JONZZILzfpPUUxvAEJYtyHwRwMb1ibJhc2+c8GL74WU296RhxQrbXXTOQDj9NsenGBSxlL4DGrB+
M0ChVKk7lqU/RHS6EBmCKTnvGXDQacqXvlfj2/z+dE/NmOrktzDAgghc7Rsm5Q4cFRhTV7OaJ1Bk
/ERGIRVAmNaMYt0lKVr9yQj/ocZiUFptBrFqDVaYnBQvt7+vFAiHvHwnrDHY6c4/+sugnW1CeMEo
5zX89GI24Ooiq4CLbWHq+9RMWIOGahqTkozBK2g8xjTsX7YbhCag7Sxd1vPuZo5vgolc7cskMkgN
+0rXGP9vDReAwKRMFsAYlfj6FVSoNNxH7vXPgpocJo+Xf6EBOfT+RZvKZSGsNJmii+ccX/6wSMxe
+Xd926RSg6f4M7AmyPjtL0TBU9MD5YK2O2O43jQw3iCw64dTJb3/E3cbn3LjU0k979sUWV9oPQcj
yVGO6tOPcd3S4jJacMvX85szbHR4B3TzqhuCdtbreI+2CCrQpURMWGu8DCcxxVc78p1Knx0iNO5W
ijcZizMkmMKOizUiPbIiX1HETfHD4//8oqSzd2Af7cLNs/H16N/4t2QoMS7p95FinvS3eISdaKb4
AwQ61AXFZtpH6dGex+KXeH8iVNk+SJlCZ7ZowsrUhheBANt1rKPg5N4StFLCqkqz5LKcCBmFTPPP
/zIIt2rWz/iuNo26S2nhk3W2+i0muNIJLm0t2HipcabuARDCRc7DOiGkRhAJi40ux9wm18bKDbJd
Jzjrd/h+beOilbmDZYUbt8cDtJB6w98XWztyBMoUUztApUc99LrZaDlHeGxKpNIUUGW2JGaaJ/Fg
xW8sM8doR6DdlJzkZSaNS5eOqy1Oq0IWoPh1VUYd99Bt3E+aNB7sE8Xr1+jtKsvMXWdJIneChTz8
v9wyB4P3BMGgZDTU7SYK+iDIjg+a2EBHIApSrJMVrGP7TcLwj+6m69I5RMbnsQopUq62vJJSiTt3
IZLRzR65sdhE+iTwzX9ukuScB+OOt5JfYdbDpudTyy9fsOiwL4WBWvFZeFRlKkEeh/HoUkiVJqCT
dYFwCq/LJttlbvcG4ZUMwKUeizQC0YR7bPO+QClSMvPxiwoWGrvGNNU3hJzLjSLkSyf38CUQeToc
09FyRUMiqGDLnCZ/AcKn5FL4F6pb0wZZseSRhXA68Kk8Oj2NxMn4ug1VBrNMInHqOJW7P7HTu+JT
bCZjz065AD+8ymQl3PBxK9xCpBXcdwRId7R+TdRlyySPJAH3IuGvB1FyxczAm/C+5Sod8yWj962r
oQKiN0Q6mZjbMk9GJ/xwjtLOBU44dJ3ToJn5x0A7x+nFdY6gKmqwopHtlrM3leo7bnLd3mdkWPoU
FG0PMWiJ9DQYGJMJLxAF4lOItz/KmQwdDLX8A3yPUAN4mNv1eahc0OK3cgB9Uw6+CVF1A6kMCNnJ
udL/gcdighIVxpZY8277RC9BngdGtKA5N4BPezPNYSM+cY/TKEDSVZAql1A+g0FbnLKYBOde1QNV
tpp/5e7vZDcDatYSx6uQv2xXX0jYGmqaf4CoW8gDcZuucQ4LXPsKREpeHr0sr3mMRrTWhrmiSr6G
zEjTx8O97hVHLDGnN/fdoMPWzDK8ekxInGol38CrGWc7uToHlUAWWzN/Q9cMwFtGivJiMinOFepm
jQ1fO613RzKXH6egwyzkWGbaiMCfCL0tWK+1LscMqj6P0rzVy7XmRJjMuxSFaRyVRUX89g1xJAY4
2kZanYtwhmQU+f+DSfB8Oap3ds3IHRJRbzlJAIhg+F+jBlyuVJk0HvkwmF/PhXI4YI2gsh9oeldK
slh1yT1UTPEmXehdcSyinq8vf/SqjbNr/yIlIVZXDSp/cryXxic1wIyz0l0ZyPQAEJ8vNxoAQ395
Ykq8SgJ09A4su7IOU7GSItohk5eF9kyJn8iNwqSWJUw9UhXTiEtz7njPlsPOOo4+piI67iJncFIC
y3SBg9R2zbCLjEftlZ7cwSWN4VkaXF08j0Mp475nH7DjjgslFUtvwvKR0ENXAgGaYs70JKucL2zv
AJ3+vIVuwuRTcXWk1vl5ONlUUyytrOLhdagPqniqMWqFHZqd4Pf0C04i2ZVpcGDyaTi22CbTSBtl
j05JrhKGK+boG3+BS19xNYUvzEKGm4IMpnUANsbV9kYqUIB3elO9VBlmguauCRJ1j2w1EgDjholk
PN8UnTPojV48ERSXwr+6Gu1tpp0MycHnC7WodYtU36a53jjF8vyFq5f/vvdGGEaMR4w3e8ZNRez7
SBKbf2IRcxNUdRkj+H4DTd67ruLwN3alne5q4B+KsfQHwx1nNF5gOz6UkqcR8gnMQ30TgMBgMUFJ
e1dbwm5JyhPJnb4KphdI+07nuAAWRRGTj7sinOdWC3T3Rrm30614g23+jiUvvSG7YX+4UdOHIo0k
MUb5L7rylaubVsOMLh3eS5zH3rV2hcOUJUKMDsAbBGz+Vhy+i7hUGinfXu9+dQV7p6xZoxlljo00
bZVMfDmFp81vJZqjwH5YrfuS4GNyZ4gUMES+MX9OwI5QspHaNfvxwhdFvZrgZdsxAEJRh5gO7kVT
qxkp3kDARMlXGlzzsxBqxgRVmPYOLGe9cvKjRmBuOyQkQ9t9Hvh5kNBR0de0vvk1kT9nF16PMTgG
0cQuoPyE00NQXlLM+2cABWOLDU+oEqnwbgvtXrqW64AyZv3EonH0wZx3V4Tu46OSf5mz2PRzFXOS
+nqf/P95qxuAnDCEZOmIfQilpxmjX2rDDJVkhyEb/sithXnFXFn2Gj9AtoYogW5KMj64Rj0q907e
R8moY5swg4b/9bECOFgJZCEOGaBkkQJcN07FAh9UR9F314QesE01aFvgcWgvHLl2crb9v6cBRrIh
5lhTwVnSRVIFDsFtcgfNXNrQyvJ17F3Apigs1T6WVTLn0FvXIOqVgbReidtd3ceJIjcwm7tIuyqQ
HKsegyvTka4j0c+9lIJknrJx2qCrqNmkia7Oob3PhwCaWKfl+MwP9sOWul9Lc5cqMYHXr4KXH6j/
NUbhKZr/bkC8Kf5ILnN1mOHXMk4fJd+RxJnVbaj+w61roxYDdlgYxvX0dTW8DDsbJbV2AMhn4qdh
Fa4UBtRM+XRbg0CyFoKbhJ/+c1p6b/JXFskGVUOoAWahSq1bHgzfLTzJQ/zynSON3bkBkp85fisF
3WPUSoY0qrfL1L/5x8ToxZutlpqOevRD106QL42bI/vAh8DH5PCTuZIVB2biNrHWAgUS0iJZFyo9
cdaqLDdrQ3PrzjZx3X6Z20+qVQ2bDGdcHl0WQzLohx2gpKCy84lYs5usYxG+vmdvKVdYc3UTVp6f
3pAZLxA3q6aA8LUrrE33n7S3UAKIn5UgxqPcDZ6Fo2qY7Gc2dIjpd2LY8J5FcIvXZ64vLOEKXmSt
OSQVidXbVh/VLnO6bk7L4j/p3oGLc36H3sEptYZReKxDt/sOCFS6ffKQAxYeB4onzCPSkfQ2BOaa
3lJpf74yvoFSxhfRfrCYkglxQruMRGrcJWX1A1ePVrsJjDxIvXpnIq7QH9IjXqUgWZATaVLwHRTw
xtYaWuX2pMHWpeE+7M/1/9An/yfEav2fH+g33yP4urjzk/4nT8RAi5g7qocd6np0qqCLpZyU7Qrt
4HVj+uAakldTqn+/bzlAIB2+u5haglvxGqjCfGv9WRtqbZeiiwYyeoo8NKAC/DubVW/9PJJC4tcr
5wo6/yv3D8eGXFTRF2lGJucB93K7Xc6z0BJcxN56T+I4Y2D5m+QXZn/kh2FqTWBhpGWDKIXhRyQr
vGnVApwujqdFtmEkzkL5kDEp6E+Myqa6x+GrtSrmJ5HJNxElOYoeWZSY3jsIR5lY96/GGy0DkmLL
FN2I7kdGfISE42HcjqjJ9Dw4P6J6q9yIFHY8Kh3NChUYzfVfWWZ8c+Qepopfts3/sCe07hfp5IrB
m/EFUJTE71YvKbwUnuJaL11Tk3esM5feJoYmz1uEWm0/+kHmL2Z2zoaxy6o6weF/c+c4wCszvqQX
PNUNTC8AlysP2pZ732I+pYql32AFP9ffpdeNwjwlJozej+7t86NxjF/YiWoc9/eHl1V2vb2peUWp
bKFC2FgZ3M0Otj2tgohzcwuyvTR2YiqF7UDAxwtMpao6dFpE+2AIMdy7oqqwfks3Sk+uL/63t29l
qKeLIZnOVnAFz8nc+t+vOXibmIrGD9ZywXzy1jwUIiNRvFRn4onIHBP/vFUO4Nv25yIdm57FABO5
H8kHKjXHKeEcXpuhI0mHFT//niq6ov7TVdhKXP/2LB/3NjoAo8UE8120yEgSSolwBml1uLS0UACq
a+JB0FvELyjoH44nSqw4/jwEz9d7DY1Mgb2atpnFHwe1PBfKrlta8HGga6AQPBouuoIn4YyLKtRJ
zQlxdT0RMeR7boqL6HmZOgBHvFbq1aw5Sv56pAwO1cqUl6ZAekB9hON+xU9XOLUZYxdo0f5YQeSt
hawVG4aGJtLSs+QbuGQq0zAQ2xpoGQKCCxNqusgLlMznLeo0M1kVNp43hdGw441mZSoxfZRI3ELi
vlsPsLT6SDOMDpHM5gQOFekncAtNPevw3onKJGCZZTG+OI+tLBWywrRExxj/EIZuyQwUwRJ8GP0B
e3a0Psefkoicc9M0dzJzofCloDpgfUz5+jHj1cCYOBmIPRTaBGh8fUKslmb/YZ1zJp3ZXBC1R5s7
l0jGN1v26j0mA+zcx9pUfYLPKorawG0XqAsIwOiB6zjTmEIipIrosh6oNbkDXwaBSvIIF0QlntqH
nOciHRudqhqGVOwaN9c+7Y/YgOr22l+/pNBrF3SJA/w1juowxrVaw79hiyBHXsqydKD4IqhAakoY
GXgw0+mu+nv0SUd5cKfQpJV1B5QeSUxdWMB4me0YxKGnoEIm9P8iNnUKYS6rWHLvjzKTKJOhQbbp
r6ilvITcq8IdGf9jwfSGbWq0xfmXHHS2S24IaU+zvgp+04A604s5CKQFw+p1HFD42icLYjGg0RTy
+ZPpP0QxldG5MMRtGHRpsPwymH6oKV3Ny8zJc1BpSk8kbu5Jjs7zSVpjKrm7psCcFi9jIB0E1XKU
E1Kkxh+TFKA51J52l6tyXQY+4fISo7HRgGaNtGhJJ+g0tj7zlFew7bnqdEzamnoj/3LvMvfUzfpt
Io1/uvdCzCG3U2sMI4AZ5+AV+D4zoC/Hmb8NZj2UX/KpU3ck659nPT82fAqj1PPql0qg8zX1HXUC
4tR9lyb0TYuQwdFWPWrKCmMTgrTY9ZElwI1NNZ76oz+tjlely3/Pvp/eZivoCSfb43mCmMww0Y+L
P1HN/S+XxLOsxLAASvG7A6tXeQs6lWFVXWyM7VOh1W2+ZTldKWPjsEJYHSrY347orxYXEJLFQ8rG
gYCAiNP6zOCx9RQRM4Ar8hbPSozu24PKE24ByUKdh4tFfYBwkOMG4bX5QkjKFuVZ+4XY4J92aUw1
fFX1JIqzOq/yZBclYKNqgUsqVFmJ+UGDyZe0Zo3uD/H7Wa3tU5yIkuH3cj6YzrL8BqY60yN0KGI3
oUD144FHMXTHnhL7wX1ZFo0126QBhNcLu9nW6oZ+/YZvlDWioF6i+GFZUU4VxK/iGfzrHCnBHzbr
ZcIi0WmPO3qD64bm+lLHx1z9a8xv0PAcXmkpV7g9KTnb4167IkE/hiSzq0Ss+ZmY7nY+a9EObIB2
5Frv4r0graI2m8sGN1vBIxbi8bzqq1Pj+2+V0JWsP2g9td+RL1AN8izF+T7rBesQFHz3YWtK9xT0
K4pHRsEu+ayMtfG0fHApKO4nGVl7x5H/GwLcxs5HDsH9aGpU8DHLirvqu7hr4rjwCU2zg3afbopB
DrbUC4j+UlWvV55924vExcNyBCseSdBqe2OBkwPjEr1Zhe8Eb9bjhXF73ysYQol8DYUNhAoact5n
nMhTwd3nIktZ9dJMUz4O7lWCQHeCB6Q6uK+/en7xp3c35h6YxdszxYh3ZvCImGaAMntwUgwjLIbO
Vd4vOz3Y1rtJ3a19ylnnTs0IeThkInEF/Dsd/R/83AsG83eAFD/cfgLmI86IOpL/nlFNfingR+DH
O3QPeuLll7s9zxvnLA/RVF366ZJeZiB8lezs5OW0KPL5ewQmbPq7uqSOsUMV+wYsjGMoVh6EeNiP
4g5sP40h0B+clSv94tsBPlJ78Ph31N2TvXWVnQocpp8JLLkMEh2n80fiypJI1oF/LA5MUsQO5Emo
L1D+Lw1Zu2UOWIcZhhhU0QlAU4u2m9QE2CMpzI02Bq+LQauiIadKHWVDY5LKU9KMZlm6RLd5es6Q
H/3ErZe/fk5lvKgjpMUN+5zpZ6qDkeGgS/V5FFuzV3LtfF+4t7KFlZ9bF7iRy1nrKiCniVF6kDrp
fN0JcOiUU23Ra/FTpCuzROJZVeDmpttYWMR6d1WTQ6MqXxSaUMw6wNpC/gsRJs1C36r5kUAGl69f
hHugYTTMSF561vlIvlkfu4zpWzjYZMqjH2B0I5ez3cLY/CXDuKd2Qb2W8iyYBDYhtvRe9DupgOWf
dzKQcJrHdw/wN/f9LJPaOiR3wokCWuOjI6/6bJPiy+zFK0MEhGgOqAEIejv4FRSYqN/epPP9p5+g
jGWSCYXScMABjSdMOXR7GYWYe2xSFpG8s5CeYZKEV4h3SA2vfufDR+6T8vtJ+7RVXRW5aI9JhFef
9rI0CZwxuVRqrA6nmjOR4b7+n2IgPQn2eKgZ+a+C3062pOvp+v7gZB6eVeh2rdXSIeocsvke1fzJ
Nw25URN3a/pg+l62FGxXhWFPkWH2kXJrGwnH31IfS9O2JijxVDkzlHALjd0tLQydy73yS/ma2nrT
mbd/tre0O4zjMWqGXpiCNPDwa3dlGFS8+szV9tdD4pPZHRhJTz4XdGn8AJcMhzR8+fol8HBo7pny
M7CDuaU2RpcrDof2AsznD0JWc93gm1iVtTjaUEpbzyeYMGIkOYymGyZBoRNcRjGth/+ce6tmI78e
0NcNZVWKvQedBtN6l/IanSOeQsWtl1fDo58RTe+vcJwYf5fSrvBUiksxgYYRWHlFrRmWGB4veXXz
qWhq6RcY42EBdPiOa2WcZgCWLEOB07VjJaN0EVcYvymnfsGC9nx/2AGSK3TGVu5uTPoZ1li8RIQW
5rSvhIEd7fY/ExyrbmcjJMTupfkTf5KMZCZhIEqTQHv58Cw2JUr7x2JomU5kwrJlAHhs06L0z0EP
O8OTxQq8YE+5A/+uUD3k3X3yPYp7dDb1tONXbiKyndmyoruMzZXvpwh7EP6K+ancKPIKO8TnBJlO
N9y6EInYExVb5p5kRQHEtI8TpAOTGyxmAGZg/ECeeg4I5sTAMJakMafyY55Z3hctJJcUi5ha9Qk5
kOOZs+cacMGW4M4HNMyu2WMsxszM7vzo2k9bGT1lrD5hjz4fT1ASXKkK0Zu2rYICDbm3YCX1mvEj
kWd6RvWX4Qp51pVhfzAqT1GpxUihmNZFWtxZCJlTwZNA20NBlwRIO8CoAH1OUtclexU4BD9dBLTT
oJChty5OkfRZzmCjbf64wBSczth2L998I0Z6YJoVqYApEXAZ9ynBSvWIRLDH8qaQlzAycWcjbp9H
uEVqsDbmbefLdMVHvpjoJKcaA3X/nGUJLmXXM8bpay+CIbJ4XeSHH03dyWtE+KXmHUeg3EEQA41b
xa65LCta8kq9rlxgrypOrtf+otSst07v476Ov7DTu5YegZUUY2a2HyATnxYWpnLtdnknp70ukIqW
Ke+/ODegGZSfL5kp8v9dsfHQBlBcYSHHs5pw8IOPptsVsFa0iCahylyI+G5v/XQlMktQ/8iEnIEu
4M7deA1thbY+oRINYvW0hdbcD8AC05Ggcym6yZtkBbZIROWV8rNWUUDeljw4tqRe5vri8G/6mXh4
OIRLlxPP3P9MNUjQUakqhhjUTQJRXWFjCzyW7OHFULZQQSU4vKU5Kj0Pwd9JaWsWgu1k7UMXB8S/
gwX3VUyDk+ubC988mG3/vmg8WN7iZxOu7eGX7b5lTt31BjhPqlGnZCymiGGdAaMJWQmjN7wG0LaJ
eta9OutFwoy3Amx5+rNvzDts+hLrix5uubyYZ6z7NXGCaRtFI2k9qwp5fDCnJYSfVBe8mTOLZw/Q
yAZ2o1VuaGsZOtFeSvewZouMGrQCHqvU50b10NsGyt1paPYf0FHfpHM1lvQatqnbl1gukWUiNEeG
qr8SmEZfZSaqADC5D7gn3PVUUS/XKKkVuvPwWvU35NhHZXQE6WJHwulqB+Wj+C25cVZWxY8JemxC
2yGaHWwNbTcdyM1CCgNxHEM5pxBbMU+Mtpvc6BKetWnWnrKjmDnIoagCQjK4FHUTxVY4QlKYScSH
8+P5bGr7SsNuMckRT9C1egLF7QVqobTovH+fdj2xHc+R1bb1/p/ePDUR9s1e3/1USDAq9qn2dhnT
pSZK8pnUYEgatZndjkIJCOozVY4D/C/U0TDeLe6m9CC6OgNQX8pogk9wduaYS2pXX1ER8m1o1Fw7
yaOaGw9LZ8K+vqdwYc1vaLIx/z5nK3mP1zNiGMNx8jzHUsPWEPm57cWC5mIJ9GCCenIR+XfD2LJb
8ntb2Qr4QQrmrfyVXuqO8HSmYhsdna9+i6mrZj42cmNfwvKNFyFn+7ZUCDVyPzyUgxq3vl4WPt7D
ta0lXUs0u6Bhx7hOdWXuWbcqfYDKa87o388l6gtV/TkRfSq5JxkJjz++cT4GpuAm4ZJFDAXSrTC4
MvQoM8FCn3ajZItG3LxuiCl2nCNqhRuAJrlgfEM0/AAWJa9rEQACiBru5BxUQ+iJYWqRPGG3pmGR
ZOqPMhPl+6mM/afIcaJIUigrg0MD4CEZoMij7wir+68CHF1oG8WQSuX3OAMVC+m+VC0AV5nh5ORb
UB5WOmvZvQZVOBrSmM42MibOOcJrK7qnKvSaqDrKk29xOzU/UMUDpFntj4t8MzKteBG5KYiPLOB+
nZ1eirzwNM3Xioi16HhRyFEFoF7WPErPx/+4Yb9QQxVoM2dzNAPIHIgIFpS3sIJ3z0qR6hp4LxQ2
6qa6iaWuFKlyQEHmvpBA9yx0f2i+cgyWKZXQpeTIrK9Fxp6c/w4jgjYt8KPNQRVGpzVrLbRV8b2d
n677zroqe2tViZWI1sUQVneVhN2oovhzCA1qachuufrRfd2LQveCZhgT1oesvRmKKruBEXyBzNi5
9/ZSPxqRhoF4WuWW5RJASwg86lOar1U3pXopgFqmAf9/SRW2aNqS9tokywbqeMbBj41r+9+5xVn7
T3LVJNJ36ZLEcPYvLYLkdQpdphPifEwPJ0OEcHBsQE2ESM+F3TDnv2dkQlxuCWD0seG332NpAsvI
4KLHydFxRCODY74Mq2wgl8teT6U/EfIj7UO25sg+nZXVFdVQRCROb7oSHmDDUZyhbuTrt8JDFkhw
s1UUnXM2beBF++/9UocfLQ93f9rRTFZAjv4UVMAwExXwGh1R+DNnc8bOt5JX8hWRI2zYIvYYfvch
XHUVmTlcUFqK7TVYWYsoArdSr10Wg+qGK7D6KL3vkdpjEqbLXn6TPOg3RQqBA+Fdi4KunJk0ujQ0
GqX48s4cxwKutGSyKHNt9yWG0CJW32E6CKBeEzS9/OhbzmpGd0MD2f5ksssQK7ykzQFAoYoDX8lX
zMUM+Frnq22VsU6/S6Eq8Kp1fHtkfhg9N/kXa+vZvxaRpHc0nAujOz7T6VGQyOWGNfXZ1IjEDmrX
OAHF1D5Kjo+3Bc05A9EXNtaNEip0vrIl4hLMFloazVPgq/F3BTi5+P/SQyoxLlgeon5IkVGml5MM
VAAt1INkHrtWju9KU+C7XVtNP3rBgjdWsA6Rh7pS+GFtWI98Jk9DBYlvgYdaEB1xMN5bIdrTCmDY
DmSWlDJDY7kAgjN9p7ihQZfCayst/fg6clqoo74IJEibkhWhvixrjDM713GXVYhccCs66wwxpHyJ
aJvMG5hFj8/em6bVzGkG2bU4B4yxBdCpOM49O5HXFzg5otyfMu4k0E/dZI0XRLwD6qkp8Yn4WBmP
PXKcY66Xst9aQ8iFgXxa6z2348oA2GJR+Cf0INnB8VixrK55d01UZf9b7KHX5q5MBNPvRmGAUE7o
G9Z16nNbtPQdXngutmQgoVCikWXq2TvLCBaHClmjplMCuuEeC7znZBSElqIkf0op6//+NH4iSdG1
8gePahNJ3FSzelG3VFPAtX1AOcHBWFCvd/3+f0cJr20RBPtbJRSScr8RZcOBE2Aq1eWUB1Jf6V6G
F8hJYg03VrojbF3gUx3fK6QwgZr6jQxSp9fc7ymUFs6/YRDSvYZv7Duc4Xo+0x3QJmH5E9l78y4E
hcB3XL1GR4fempIoR6tCxasDJZDXS9SoYnv1yEejuvCzL4crLlwM2EJDXCma3nDQXWR1g0U8UeKJ
j8n0GSdFE0uXSqmP18ag41LnwrmnTjJHoVy/FzePyAWL4ApO0Rv3Em6QGY0NMpODrlgrsmb6v4u1
DudPsF1er8QT3uaPgibnEmr/YfcRft/RohFdj4pkMTmoypPfa/Jzm5LpoGUXonkoP6IIFcXEiYIH
mho3KDDf2PD4BfFs2O5PkntoFcO9JKrQgkoUnQaUQDOuVmFnxy0l/n1IAEu9f1YqzgeWpUPSHYmO
Sx0bx55RXCPIGvppsJmXOfLeqoE1N7IWNv8KsPYHRA/BMnyzXV/dXW4m47ju7fZjyqvJLSB2/Up+
7X+yHhj97nZvhMewTMn/E/+0iLZrAgm1LJB3NrVRKJmxUBitWbtE10PD761rfXond+j8xVcx0QwS
ds3VC+HeEee/Er4eYPumURn138o++NqDzsKTaVuby5A97wEBd5N7PI+3uZRyJBBXKQxAGpBubMMX
sPkBorwym50g1WyFYQgnpcyNF/BBv8ciws1aUifmbLhlt5psR+z4XuvHTFxaxAXGRbnHr/QSQnYy
bWtetFbNsTIl4mhFhJIxr6Z7OsbdRHVst25JhW8daI4GK4gOvK6FwY2yl4mX3/ez2AXl4n3o988w
kFqjhgHLwZzfpH8MMlmLcG3ZLApibxk91FyvQBMgofpBIY6d/+2rWSwtJ+0LaOkUdysnOczbKrO2
hxEbuSdV7i1QuwhIUMt4q2plTb+KFpRyNC4Q4XD0O/hcvyj8kmohaRUQD5yAPC7fKBcEuJIUwcY+
Z8nQxOM2i6RE2GVjHHEIkh/ZKB9JqSjfsMsfSsd9AanDVsZByJMSr1eUUq8XVE+sBmNjUxhFDgES
WljixHfD4ygAmvjyaXCqm3u2GyrjqQ3baDiL/iPRpSa9o03PtmFmTJPS4+Xtz/miBUzk36Vr2AgI
Lk2EhPqnuinC6Djb/aww4DZm297Bz7AIdBrZ87aiBJPIMIFvj7T2/k7vwvdDez8fRKpyn22/F4SP
d2kHxTuhrOK3Rr1gGM5Pe2lY08S3Lq8t1+RJNzxLW+B28TRQa9PcJV8rzijSFh54XQqdBw5MVUU6
b33ITQVmBZivANY3XIseJ4xKQyd8XXJZnVhcmY1MB7T86m9MNG9OdnPPK4bSDnWNrYFqPNWoe5Y2
GuxaU9Ldp/qu3OkWGokRA8F0zBM+dsHYuWxEmKn7zZkE59Ni9LGHjdygr+ky9590cvP6IJ5XIXJR
70dc996FedYlwgZA59y2+mDiA6VVICdv1xs7jSsV7mCGUUgcd4GuqlG8FTDDGlErnAm27KOd9/+L
besEEtGjAkKVQuS+AWySXQ53gaU2wf81FlCSry8KqH73HJUKyHlZVMi/ymBikqc+Ys+lWPtQye6E
IY783xSinADG4PIQjD15HHxOYaTzI5aFraSzg4LBAs+z55j0Je4CifbcFQk/nMibbdT4e0ig924p
3pvOnih6QuqHQrPp8N8jstXvyRGXj64XwdTw9qaQiz0DdDNDchkRE/pAmGRL8lXh/LyFvxHC6Z+V
HQ00/GyN8D0IjZz0kTKivaMrsH5NiRuAz1DMDcnwuGZ4MAZiKNhYEJknWzFdCHJHXf7jWsIxpTwA
4Nm4X1HTEO5PTkFItBv97zMLQ2+VeyxldjkXBB/QrCkkmc/LVaONoXl1r5Xz//2m3y51k2gWrTZZ
Kw/KFj34QkwLGyfQj1f25o3G+hjrYDJHIcuOfQrCSBLF8e66tBSGw7/kQn2xJ2DcP4Nm0D/nYG58
iqfpDimpRzHpsC2aUx+XsLmqoYGQksMj5ZdXDxJz4jE7nuyJ/JQh3e7UXEL3V/41Wr153Uwctm6G
4aRn1qEu0uuUa8yAMt9ad34okGKU1rB2UTsaTf0xTdoPltP9ST+pt7bSdHVcpNmmi+aKjGe8yCtY
q4EeSHHgS6FqCNXQ/4Tlb8jsvzuFgNPZ/jPNKT5RY2100Dv51K9QejC0ozrZ2+iXoppU+h0omfxA
Jr7xgXNLNIxp4CBbTZ6TgNmMs/FuSzxabXi0cFVLghxKxLgF344nf8V+liHJK06ShrG8PC+h+NIw
AQfbb9zpeqdZWKg4+AAx46rxo9fGR9VzuHNygjHxz3BfbOMpcXjei+xiDrRwQNWzlRKZZOXskwLb
FcYHR3y3FwHBrHAFLYEoRb+2kBWHqRM/aZou9U4msx8lk8IYrHoW7GVkt18VbknA15OHpKDTfd90
QyL0F4ObI3h0BZqlqGKUGl+qKuYFmwlzHUz4A0KNvlplVh+/5v4E5OuumtKpqjpJxIPW6zzfZtvJ
gGAV/6rcZdiIuviBT0Kyxy9OhpSJCL/WwdvnnRulEwHmkYjrwzBQBCEriVmP4ljibNp9i1VbDN87
rpT1sHgaG45ly+iQg2PKAnMCJWdrwXJIiLHkx+mmgZszEStjDVJD3iGYxWT8BGROApiiZg86i5qw
XMgqCszDPrSlXg26AIsJmSCfLIMHHFynTyX/qMgzT5PNReJGKDS/BQsg60KzR2SArGTJQCZAY57+
E4+irN+k/WFfQDXHd6h8Zn5T2PCS+j0pizAsypkgwW52BAaXryCiW/D86t4dm9l814yhrAwzmS5R
lgoQegI9A4YcGJVEzgooFRViCIoVaZgz9cTKGMkcY2dvsUcjR00R4/ON1usvDU088YKAIa4AwrfI
ykzvMYYjcYB46FuwboWrMWC5qzshPvziHNPq5LRaqVI3q2P2Ird7TFSIb861WhDwnvtaLHT8nofU
HUg+9a1artvkf/0idzTK2BS0xmoAuOfJ+t4drnMNvX+zaxGWpZ0M9PUYaDFPg/P4tVg6SVVPa5Hs
5b1Zy6buEIZ7tgclCKCEZ6pWrfRvjj2h1YSTdl4EDIKfMw1OsJQGy4Hp8MemvwBZg9UGnF3fhM+y
UlVFOKzH1C6zYhTZl8W9zaMv0Pe/IyPmYNpc1NSwL1foi49f/aqvT5tKa0kIP41zb8yry/vxu4yh
SPvvhZZSrQcQvl9lhAvtM5HXxWe10NK1IwAsRUSWicIWIl5PKE+CMeGpLU9KrTxpPmhGILzsyCoQ
QrBt2BRyUNvqJ4zFMRmw0Nz9rBXk+GP8ns5Z8nOlFqD37l3g8DX/abHXm87L74A9CryITZOP952y
IDvxkq88zpf24fdZKaUhraijEb70oNzlPkk7p+XQVpp6XGg0izRazQ0okPrT3u3Xufq36VMLw1nz
E0L4rc+fYqSC4o6Ki/oAlemOM3hwGJWiKBCA+msjJqLqWutUNbnMIpKIGizXwK0lc8Qeof3RublR
Mq07klv93FuE+uXSfb6UhwvlEIFLNSafjQOXTzDgv+ErEVKMEj560UQC3dSjDrhWYDn3cq2Akx76
+PqVNp2Exu+OmLlDz9YzFBrAPPlCnBmp2qN7qV2In/CBBkWCHZ5UFIHnhSHlR8wXkeQmjedRRMxH
35iBZRaaQhu7+k58S+vXtlIptN/vC847cE3/SNRZbFU3SEtslknXfStCwsWM19ZmKjsNERDHeeCF
4W7wFnI7qARVMQ9mETy6RWDZLq0NKCRukDZKQWRPooaatIUytpFHzu8tu5WRn0vYmPPane0+l3Gt
ItoQEFxbo80IUi/nOdID+3TtIhUihGUQnnSiscOCGGuwN/3Vz/zyG0WMXZgiquF7G6iQEkjYX64Y
/HJUCnC1wYmxP91zwxVQ7yDgTk11wawRHfA6ADV0WlAo/ClC95ML5avJ4Lfb7ojrVLuUVXkwEraT
gA7Hl3nfxySlWv1Lbv4svm6WjcXFAeP6zoENStBSVG2k9ZG2ws3wq/iDF42MNGaLwOIoB1UIlIDu
9x+LiaTnb6yxNT0jKstUtNcFbvvtTEY/uDHiEVTeGdzP3EGmOrqBUJBKxBOWb6qW6Fg7UjEh+Fve
RYpfLoUAQXUhoVG+n8sHpl409iih2xozarWkOC+92l3oGm+knUAebgUV1HYSa/jVVnCT4tMR7Vv0
Hz4pJ05prtqyaw3ZGQtG0EM1q6JtO+GxY113oGDluZPylJPLm5OSfGXlfiv74EP7Og2EoOIA/veo
YF/BKuxdOxsYig0jyAmIsG3uFodI/jUZvJUj4/ec4UkyjDvUdU4kto9r0ao9F07fhcxKmXmRY8QC
GZLJ9fuXLF3hKRLufFCEOGxQKkt2iW3/mJj4kcyypcFm7h3fnYyJeMtoDaNuPb4Itr16sZdJxkwb
7wik1j87sPni06JyN8MKhW2QgK3Kiz3yGeEJhGoGkIpoqXugSoUrWWHu3evqtmrXUWFqSxlO2cOu
oPnjJKySTbW1jadP//iT6Tc0m0tN0+syt/PPZoyr2+dmzKMDY+L/wWDHRrddDNgk8ihZmnccRf7o
WhqndZyQE6TOoGY8SeALCx8J6aApfHqrVKASTSrxS7YsMnuRgP4YBkLYAZRt5UsY/Ivr6c3anVQ4
iJ3d8N3ds+r1ShvwEWLuFRmkuz7cTOan7uGcWjKrKr+3c5FhBSsx8TRdG/OhkfbMffb3QRZhOldV
h86/4TJFHakyks496vMYQQEvua2WVLyTsyxD8fMwAFIPGg8qxLSRpGoA8SpTSRWUXxsQLuqOmKzF
S4Olan959TFqYuhjAujwv6ejTeSs74EBqt2bb458DV8MyFcXK/Jz42BLlrq041Gf2eYOqmY+oXEs
KKwaEgEpH5sY38pDbtayEe0ItNYqJOUeKYFWgz3FcUKaCV2ZXHlAzGJL+TWLz29RGkivT7LBRD21
5NOQYUuer2NPbiCuEI+ii/3EEQEAkUZAOINroYfST0AvpqvvooWatHkULhGdjTscWYZY6n7ni9v5
AbWebrHEyo4YuMYOHHqTluTtQhJExPcn2eD4tjhtQc1p56k0IVzYj+FIW9bTyVgprZ39PXiVvdbE
sgvaMQrayQfh0lDbh9YhuwvDWtTaVC16u/Ll47ldn9TQWRzNf9f3NBuE9cXzN7r6mTTaTY2zrv6m
tbW0zh6BabH24YK0oktaCT0dP95fYHEkMtO6NXFRwaHg+lylMK0zHvQVHhZzh8KHhw0qaIwL1rc7
0hM4DTxptZ3Th5zqJci+pQr+ke7iuY9f1yiQJxs2j5z8ozC3Y3L97Wc1LJcmcnDEJv/ZO5Hix0Pg
CoHyBG78Gm8o5LLOvkF26VyH5ouCUgW/3OYGad4MYeY0mN4mTicIwFigBWnOblgD9IH6Q/Q5EpJ5
5XUWu2sbFlWxH4foR41KUpp5o19XDJM8kU1Dx7d8kW3x4Zn8RkqTV47S1LZWfEx6E7PK13BxOjgp
5JnIAQzwAvaeC+aObIdA6yQgiTouKKlFWWT9A7At4EzrCrwBxIGU738xhBEjyjvvAERzWe2mho7m
xfhaAEWf4+d8o3ogJHGuOV2Q+c2oTsSgv0QzkWlYpxRzJItrp7eEydOraUwVwTsoAEUh7KcwmHI4
dOb1BUsl77EozVqEvct1ixB/MbrWPl2S4xtWZFmuHy4FghMwlZwxq/ftNFPVbbeUal/Ff1Wieheb
HzTQZ3vtpGjG3tr7AcQ9jz/W6vPrBnIzQ+g8Hr1tue24Be77/FdVpfWkIYbcV4HqZL0bDpKuPbvz
2JJ9jvJMLK+ES4CxB5Jh7W140ydmOytMYMX5EXQQ8yMppUeqMXbRe6/U8zEVls0fzyekZFhQj55r
unNpvGNHazbQmyNuBAQ2upRjlqEWYWb3n/b7ULk62JYLx8TXo40/w1FAU9H4sahdGckvVcN+fZYi
7+wjAZV0QKmnGAUr4xUUJyC35jCa4VbCytKkdqZ+1P0P5S7/BNdo4+3qX2NLTMePGXyD/w4AZlT/
RGtO8LizMaoYe3YajTVW/Q617zD17GFdIHD8prl4uf4D6sHdLzZtcMJPf6cUUSkLRJc252Qplglu
En7fJ3aRrF6vnNVGz23TypbXWUBHipLCozoIPkK89azFSTF75XCIf875evZe5ZoOrp3LsiZsRKAj
gxPGTZVumdnKyTK3IUo36ZwdC0WWwBghnmf+huRw3lJogJbGchL60Lkj/XAdL6/ktU1oQY1jLLzH
OJWplKab47COrPHAznMOPAgfw/gKyqaLv9CBKTL3DLtasWODu5ydgvAF+mLIXn20Ozq6ueVrqJVW
MsJU1+tOAU0xelCZF7L/D7JSl4CUcW2eqLi5Mh0zjKKitdGYwPsuD2QvlTkafWHe2vZUP+sswPLF
W9pCG50chLiz6e62S0ARP06rynu3y+trlgiKGfyOE4cCGvE3ekY+UmEEHarPb/5M770Jkc6YYxQ0
8OSBefny+3+OanJQD33ugFCknrxnekZBIONiDKQqIGShmmqJcSgWg24pgNwei/ATnW12SPD3Yulb
fIKs6k8DGp78XNsetwu/Mnmkwz1ddJT2sTJqHIfQYZAjiLKUk1e0QZ143/ffll67eK1Ruq6M9Qox
9tabPPhTd0fHcGAHtZ3VUDyQ9O4eZjMzMShRg2hXkqfOwX1FPS7rLMYgcDvUqcO81WvzojDI5urm
1PVkKJvJ3Y43EHX49h5gav1d04++Iq40NUr67spDkAdbTMRRy4fmVaHdFaYQSPpIYRrW/qKWhOxM
g581yXWjlI4s6RlsRDRz/G/zLiO4K8HUMQN+1S3JxFVcwi6V65ocpdMN3xeksiKyhAVCq/iQaadw
IdBEUghHqp9IAjW57xhQPIzPjjl84g0Su/sCvoN8KX8yI6tlniz7CWP1Y96eC3q4BAM7abQwlUVB
Vp5ZtvVbfvVKc6OJKKOu+WYlbYc4w3onXYVvAadvZP3v8PILp2x+6UrVElkvCStyRpV4y61c9On6
Y5Z65BInViidJqFwTx5ns/8UNHJjkP9k5Z4fzyDPdgAJ+OvmcAJc7aOEQYM1i79UwHcXSPJJwvSM
4XZM0A+LNZ6H5auI+6Z2MwXuTBdy9doYO9P9TnLtU7Cy9xfG0Dy4YEOK+HVas7w3VRsYqGm/AxrG
Bao8HqveJ8gSeeRjgMqEan9K/Qzc5Mui9p2AvF93Vg/NvqZJ6dnMB4uUIWXKLbXqpQutbfZtk+aG
CncaJjOqDh2OhcQbKiJheJh+CVK9EQA3l9YSxuPwOHJo+85P5bkeuEZPoqVddJ8g4o89bKDphANo
+su31X62Nl81mm6lhe53pra94pbDadNDng5plU7ZFJtHfmAV4EkOjj4G6Jj3nzI13Lpfy/Jk/3NE
rTewQ1ZhF4mXBL7bCQkv+3q6bjBC0vwwcdlqpfUojxyvuK/2Zr1CfQBPuChQAAg/WuPLJ1d8j31g
QpS92B9PKKvWB25Z88a7+vuMhDRU2HJsIPoTQ0mN0YWqZM+N0bPxjcpPFABfwRGIVmtkcC/mMp6t
OckbSHOcVmbWL/xL2Fr+32i5QrpGD8q5ZxJAZUTS3C0yptmHqi8k5w5dSDHQCDNmKy/uP9Ca9ZY7
LZ+VafTb9ZPoQ2Wd3dkY1N3R1OMWnHxGsyt+M8xpebPx5Kf8jY/G5vE7kdc5KoABxXjsS8BcevSB
BCunAyY6P6bdzspj8BZOGF0JLaPxVmX7OAnq94cWqtjXM7Zy0lrJDeJrqXUrqW0XfU0Tg58W7+Uf
XM+c36p707/qI9HnL0nF+xZVQHiKmWvzvx2BVX1gvwY4jdMyl84hNmTQEVNhlXvZhfzWaYcVI3iN
Uh6/v8HdC4ht06gl8ifO1X5Vv9yAPa32lhKU2+TlYhgzPMG7Un6WPwfpC5uNjioLTllFzkn/BoJ+
X7+moZBbgko58wLSTV+vZEqk+0ky6QgH1TWM3ADBZuJTvQmhEPv0bCsB5Fe8c0SKUtfS7KEYW+DZ
lv3TMI0asFvAcHXiiosXXfMO9vR/nBG5Z/fc+Gn9DLwG+ANC122JOX53OtLkRyYLxmqQSEpThZh4
QU88VFC1QNW7kL8ISk1ET7Wr0sRciDbpGrVI9MnERDW/v5o8lJR5OkhCFJfyUgktg2lj+Zg9uL6f
diaj08wq+/+Cpx7SHifR97hSX9CQwnOukuSVdI8zsl0ZCYM2kNB6qVyCUbaL6wnkCGailOeT6/0r
x3q4bb8Lch9PLiJoBHwDrpJJkVRO9qAHMQieNvI9mYL7Zxs5EUMG/cb7QXOIR/Z57XqWSrUms4i8
R1rdDOr9Bgs7H35964zN6MeA9XrwFs3tfEFF5hAhIl1LuPPZIkdP6WFuIkW3TQ7Db54GUJae2nUY
lFf0Syikan6JLc2PDsHvZgh3+vtpvJ4m3dHZzNQarqZH6YSHgCyO4UE8bXsKLJyYPK05SRXhjG4n
cxcdcaUWMdsgT+NgyUW4h5ZBjShs4hBToLV3OAoPkBDq73CdiMnDKSQBU4AhJxY+NHK0Oi8gjCLz
8pl3tgP3xj9gL3vg0+GAWqdNIiVattq9vOQ1yxbjBZ78JXPC3L9YNwW4jpaQC1Y+8l9HE5/JJFEu
V+6qMdViFXdpVIvH9xWA6Y+Qg8kRdqB50v4H9gNEZluddgkm6n7tLA/eFivjjJG59owha3TfQdC8
P+DSu6elhvd8ZCkesVzf6xMWc0u7EMLrIewTUYhU53KZVJNrRn8yHQ2FGjHdv3v3Hwm3w6ThNUJ+
mLX8+6SIqcgBibsTOT7X6rybSAQpLQ61NPF6JzfDNHFsYZIowiPtgCDswAnXQtVHxt0OS0w0nEOj
V9e6iTdQZzBi47lX2jd88b1+NDFcGZtyWWq+lMAfpsK8oN7sQEiGIPdrrnnadUP8pSllyataKniu
BcbwWuvI8UZDR0BPSN9ivgi29MXlXarXNjNJdORNg0RkrFmlHKrm3ZmJvuPXZDb51HxWDaFA5v9w
OSg5nbKdzO9+0fG5569ZGL3t8brM45qMFKx0wtdAtcp8+TeEkw5/sqsbtMDU4ZHrlCCCVSfLtd7w
/J5Uy6f98wPUs0kLNAL43FFdH3RgjHW1VgnhEX/yTlOSha5WfEmM99i3vLOt+06GV9bBMcLi6eUZ
ama89NpQ8lZxAcF+qgta7ICUQ0xU1aPOfYmBzgbObxl1xNzq3RQleB70D/DiBnuuaJYZFObrooX0
51XszKqMlcW+NRMebo0NYZ7HhDGK5cfcqNLUnF/NhmKZ7+pB5HXo4tH6rpC5RcOe/4ZY6ypxmYO3
BKGLVZ3rA4KXXKACNwbwXlJ5dYLZvLnTrl9Qu5sXI9aIRcXH+jneufNvIUmO0XAshmPBndTP4vX1
Fg+DXsa8XWV0gaNH1BuT8rKqsRymviT66Nsdu5ENRA4HV/3KD3doebN7VkJ/70efGHEBFSicGJlZ
jAgR7iW3no414V7ww6BnwQ3HqOf8ZAAl3jlyNAlRekHMsylX+TbLR/AJxY05AOFBgwLNZYKq77Cz
rKAHuZO6hnMGpoDmFSEXsS/f6GYXpqVmzg7hbv/+zrcRV+LXB+bzCqLVeocUqiSUPkmKi4YQ7i41
FUyNvtDPtAhk6Xh5JAsP4xSeAjpNBbYbmSPebcoaDDdD8KW2Q20YOJsBJGS468bixxxmnuxuzh9n
qXySrQ2mxW/O9jNd9FTrxQxCGSexlGqULd2Fr9yHFsacGbNOpmnVmMuqbdrHBRYK7Eey9AUPPR/c
iMzQoefZl+ncg/3K5Cts0HnhXvfWjm9CQdgDhJ/rZudAQvr12SHH94lY1udzCdKODB8g/EKJLiG3
c21OnUhhsTRYt3EZI8PXY/va6R1kfqnK+jojebphWx2d6aZ8lh85cRCj0NwvZiNisFPVM2Z9myUb
Ix5+2zqUeEcfMJh1Veo4+8n7ZxG4r7ycFv+bqcMx5kX6ZIUxD2K4jT3Vc7vPsELVS63nwwMOQdvZ
ue1+xRUGtSc379MhaMx3OZifo45cFk6CGG7sx39uP1EQi8oUMo6if0Hp6aJVFvwIK+GTRkf/iYWM
t5554qcjtp8WIFMMme2vnCCecARSLSUXgHjkCzJKDXQCSKuUyzkcFdsjwu3aIBOcga2nI9YHLLcG
5orzk2MwroqgHt5c3e+HYd8PA08u0jZQicy1cqlruBiuQ8QhSsLFdeVSiBW/qOH07BXsJzXcFbWG
ViuZ8LD+iaxYrwxCUYhfOSZ29M9kPX+BhzoOJqrirc4/4LcqrIZk/uwWyGPRsKJBxH8ajtzV/x+b
fbSPuy8OToraWv9d5knTbfAPFKXvRqrSZSTEGB3IY62aAta67ilx3JLhVHzTIOnjI4f4cueb0Wae
kCNYF1XKnpSPM8lwQ4f4MoQIjdNOIbCm2gbByTsGZOY74mvrz5gszBuwlO1dCo0t3VzP1u9s702E
WUCCfZmQ0+v1VXnlE0j/zHb4r3I0HQdiNc5YSVvxxdQuiT6Tz2kSk9iyNKhIR4J9VHrH1WKwE3SH
F0iZTHJit7zKA72TnKNx4p/IhBlN+j31DXmC+t+eQIexYX5FIuQCPOfWy2Hkkui8eJ4x4j8x1MB6
BfGyaZZDiZUFDMeRI8gcdlgnP4UUWYfsPjhQV8EW0zXnGGj+lvz3oP5u/IidnIeTREh5gHvkIYMD
CNNFCUS0q+Q9evu2sS42lJ9+X3mXMWcVQOpWB0uMSpc1MI+ovPW+tSVebEW2sabX3E/7tVQbODXt
BODU1tNI4rjyJCREHb+ZH3f9Igs5B/eAOjZAf8kzVi+wJNs/zCbwQtMMP2lKbXJG76ieiTqVAZlE
NdcizOrXNm+eVfQ2zdRpHYOGvWyXHcrLb9NpW7ivPQ2u9x/0aiTCSM+gxKFT3ZXn+fOLHDvBkzYg
sunpTBtvSb1a0vDEeAyXWAoDGRxjmTLjeqDm3x5HGuF7y6a1g9sB9KgKw1aJvttxF+n0PJP8q6Ht
90n+t1phyv3/C74l5a6BuKKBuB2hfV/Xv2fGclK9bsrDHn9aIkGUZsNj13fuylAtWpZW8OSQsPFI
dCtoi61vgBkOaEKqoPWhWNwuPCkz+wIJWN8FqYEleLGIlMnawhLsOUor6jcMS/jl0lrkvux9FAhZ
uTww7ygtSXBcHpVHG7HMHsKy9/hYyF96r5kclHwPNm2yrCQ+Txz2puB5pDv2fMQFZz5D1Zpiejie
DLzLEEIDK4BdYkSCfGdbp0Ci8DApI+owdR8iRM66kMab9/kpoO1YeV7q5L+1no9z8Py93j7LgSwE
UEyNwAmd5lQy32ettQKp32s4mDfavqXpTI24Df8rDs1y/eY9BSXUNNpPCnSGs/mb1VlNV/jZiLOm
4HTD8ii+F4zpA/iXCuWzQCj40crTk1UrvznzESkOZypfZJRAc5VxKPFamnvWDWPOi3eUV/ZEvpMa
HcLwIbRkCSeL1wnDnMSpk2vtzuV2oHk80MWMC/oSOp9FsaC51AbaeZFkj6VcwjYGXn64BEgsFtVf
O1qtgUw25v+CzHkGrcJz3822eELeqkfaxUe3yYeUrikzglc6l55EX7oe+qNXFOGbaGDJUOdD12N+
lUsG54PxuvB5rxhBUmBU8Wxj+zu1dPvNEqaszYA9FDnibOALs6rS3ffLMUuetY8XI8+b0Ajfn5A0
0gDpSgnlkwqsLnVprlj3w4HjAJdRcClUptkBSJbVcPN5h/AOlPG1X3s83fFK92RmiRDfX1n0MlLa
I2YQ9p1l+jHsG6c5jvVOTfsi4oLvqJ315GNi8lzNnKntupNeg7txNf7Fku4xvbvRJdOWBg94mpXQ
WfGtSvcwDH59AdkYc5/hm6bJPUU0c7WGXIbiZHQd0kMuzQ9Mh6hPH9BxEWVHRA2eLx3j2/frMEcC
+AVlHCx536VOIYXp6HUnKCb5X+MBbtkEIxJcODCBggltpCeqTGoC22s2vXeICScfft+AGVTzyjIs
92MvfaQ3rXmbryerGJ1haTKGXFvmkcIfxZRhEXcL4iQ+rpK36L4HfnLvMDK/yH5umMueGV5cBNl6
7SRZD5u1PvP3Ivf8/SaRHLiV7sba2+chpuTJbEEWQO2fCDJnM/QJCB2UBC30h996bYDlqn4owoO+
XcIZTF3bvmDnibxocAn9bk+sw6/wR1U7P8D9Soh9YqAERhNVnu+VLqkCkPQMSmgdUqT6E4Ct5NaO
sbvoMOAwDKDC6g0nxA++KM0S3mjzT0kie54FWFsRnPBW5lLllahjCr4+QOXFe3JnkKnM3PXzORDA
vFMQz6Sp1AQD36ACmG6ZwLgN7UEO3hCS52hXR2iz385aJLzVK9FH44SErNSn4pynzATPAMRU9dPV
RLi6AfZ6PSXyvA3bH5d93frCWdAU2lgBoksOLVabxCsICCCvM9eIY6lhG9twjrqI2wP2FyONkkOi
oCUq7G6cNu0AjBcbGvp8j94w8tLbHhEbbudjweIiHKsmh/JR2vkfBYVk06r9yvLUYpXUxmsbUrQw
z3NobCFoZIxOF6Wf8l1mwCsvnJn8mbQT2RQ19vyzh3LYI6e2mFIclj0v7FPjUur8vwRPg3LRiIq1
4yp8wc90Xk5p+9fIi7p13wbFDy25inMW6RZgpko6ovDiwn06lRGORhhoWQOMyEQqEF9I6GHXEMNm
umJwOxYMvTsM9ppfKsP6vccPIcVLyBIT4cNHKmUOfvLJzZJKq9NvOaq+/T4wl8mX+xOprPi+jMU+
As/g+Ubz7Sp19/jJvY9XP6VKG3WYiDFDjegmtzl/4nK857FC0XW+Wa5d+yNkVVHUC3cvuWLGIt7Y
4CPDpu3nZVJazTyJS0sW3jyPAPD2hTEosCN2bOXaneG9avmkRhzOBhlMdngOuO/Fih9eyXRuyjqr
C7qXgEYYNl3uu/zMYhg3b+OL5baMyr8pZds+rTCi9zA6Ydhj3Js5LzC01wydqHHLamVVK/CzvgKJ
c/xhJ5xcDwvT6IY4HZPdY5nuNe/0ZA+AZmIdIIJYgG4dOzI0FhQv17NA/l7hzRqNFarvdnaH7ocM
/7wMdHSj7Fuguv1UvAcmsk678UzF9q6OYunFEC5oPuzI73CwEK/VKp9M3VxyIkUXWGC2XkzFnXQZ
93TIEdPIAmiO/rjYj4nf7PIWAzCqlfT/+g9FP0r3EfeXVkEBTMesOraJ8KFkvS0SdL4gAGEDK7bn
MtEABvR8ucFsnSlWjDNaCUo3RMS+KBdbiTQK6ZLfG9PRtjIq7Lw4q9UrFUaj3LnDX8TSbQgu+6EA
K+HdFfKSFYEYHXNshhIk2Y1HSkz/a4rHIRlYfWp7Lj67COqL5AX1N/lkaTAG0PlVfGoeQJ1YFKE0
56E7srHd1Sj8ztY4JDVI4JPERXPceE+vxZ5R1zrtGAOW45gAmYlSs0gCF4JDicwP3p8mjyW6Lca0
KhYJ5U/qNM6suAaWe+i6d6iyC3/OChWqUl0NnaLzW+TFewNrry3WyJFbM8T5ENldCkuySRHy/spq
3vXasBXGaIP3fi/7btcALo6FlSkovsnce7pWp4nNCChnxOgFr/oZwBIrKFRwfgH9HgoY+Ah7u8Yl
L3wmAoMjlPcYDfNfpXTs2MC2dIaYd9FlGCitEz41muolv32Jk4asc/6Zr4TMy3o1FYwFIzo/sV3I
Mxxzknsps2hmswE0q936KO+ACdtQVsd4SWHLEr5sk+TpwT1ZTS9GYKlNfAEASQpKk41E53rnH+S8
p1XoBaBiYfse09aoSnV1ssH3r8R0OFU3a6sjrX6scQvlAR4t4kJwk16NEgnTdSnh1UPptraN9SYl
vLKck1UObixuQ8YWYui8RyPRItJ8S7FV+otEck8MRIV11wgez5mG//c6903l+r2RzxPM1t4/gNHN
TMHR5Ca1Afs8KbF0ZaMTgCsjgTcLyCNJCnMVbdFSiY2dNRSpqiGFOMbJHzI6ApISTEOi1OtZ/FP/
wBTiSYpbFIIFRMthmqcoLbUE5vGGqfjJN0EKh9V09vcYFM1/0p/HL79XG1DAtK9yPO/1X0h43ZBZ
BtpIuQgogjj+Li2PrJMh+16Vl+ezIVsrhCGaERvJBAojMiMrw/frz+1YstBvsJcbq4uzm8gSV8uH
IEWH0jPfv0hR4miCcRBfHCYzVikIpvymgdC+levvkymCPno9C4rQyVFEgCOIt8ud1QZW9Gipaw+G
MdkqDGyHzUqQG+gTkbrLtoRArciEpbD5yXFYR75nYdSj+QWLxOtum59p67BKi31F0F6Xilbe8d6S
Jzl0X7UlIU3Lsary3OcQ85jpJ1Gc93Aw9PP3/sMr2FsvMFNl9YZZFrl6+z2C0+H4I9GEm+X1kkQW
L06MZiEDd75u/jX7awwguEgQDNHbNq7asNIqjFiRCSJSl+aU5Ux6cpN4hCPwTJfb5DWJyEOtzUy7
eg5CADveQeDNTJ7szMPbHGBuStA24CgGJpGh+BzO6nu+FwEqZfpjD1S90JJEAQhomMrzSdWLXPeB
yHQFhYMEQQZPx2nR/layNbFKw6wY+7O+/Ey07X4F2Is3NRMpvP29RHfxCYBS3GdqoCiYuaS8urIU
IOIegROr8cZ7aqC96uLZ/JbzhrH0sWp11auLF55lzGFytaePXxGz7wNFncbGZ880jGTfn/u1NH6o
vPvq9J0iHgW7onnXqfZKJBZGuHMC8h7q0D+BvEfpJ2r+ST4n0LHwQAK9es/7VRxNLxM/GdynV+vl
alrXamzij4wFxuqPG328tmP0LZdTLosIOum4s7W4JhpTbsb9uhcuPq9HJgFpmDEVcPZiBHvj/hEd
xvn4+XKwkBMJO4IBmgMeDrgbql8SRDnmasLqmIwKrpJkbh6xwzJVZoQJBDnNCaUUtUjaxxU/u+9t
AySGDLNfULoGNDvWtslIE6Yzrmuu0z8B5Or5oRd9qtHIQP63zhmOUfblhpjsuMfPkiG1O89yBDnh
ALHGIVBwv7/JsKOv/1NrZLf3ioR0GpSqHiF/tAEn9mKMPPL47rG9s/40DzF/+mdZAY06MJ7shAlE
J33ju+GuNuchbFywJ6GfPyLUjoQLdOo8LQcVyCPsV8ZIjKZwrOKyeVZ+ORcoAPc+kYRFIqyDlb7L
dLnZUgcqmSnUDqlYl52qSe9YaH19Ia6bo5BX2skKVKxPYRvrTUjfTLRXh2G2CtgYuyGRA070k9qu
5qM+mz1e48KYCld1J7XyOKHe3xC0EgzUqFd7VuT0pr+nkUaaFzng8QNsmI/gSzaEu7ov9KB9phYG
YZwqO92if5Kci1e7dIV2vTLp/XJzMFImKZGWEicFx9pxQpxBtOua7hR3Z2S0jT4eFsxVJWuEQAK/
Fy2eB/7tYP4TkW+J06ArENBW/KFeaDEmwL+vfIalUx9SaNCz0nNwx03a4l59MP9ATxFl4eR88oBM
cD4MpQJxPlUDqYs95HvjDIVDgAG2e6RKen/mZtYKX7zcWoPxJuJ4oLwmVCFNsWQIxO4b88dLTZvj
jgtf1WjvBJtT0z8YFYWoxXYeAmdthBLl7/7Ewa4pP1A7E8uZeK10Aappg4a48rdPqiilK+jqKoGr
oP2k9RC/EeSTIPhOgo4/YfBAVLIDCFEzQz1jjHIu7iEPQeaMhdH5siiw4oc65pEpwXwNaMAalEWz
OGZk6tu3Xb7lTzfQMmrocljUJr8h3iK0H/NJqzoJjxHB6jhxKJfKO8OzXRenvXtCMd7Znff8fcYR
n7EHIJebsD7ON9fw08jjvmo8oEKRJ78TwuXVrROvu/WJ8a/FkXc3hu52xn8YxHnm6VY/6S5gDHci
Ie0RJiXxElPbo3pfr4TtHET5XXWTgSB3bW5+gBHIrHOXWr+6nYZzrff3FdG66bSt86UBiPwgetBi
7ZJ4NhrZh9NeiGyjjrQacfwrqy8BUmowBlgx2p7T884hS4YvaOkiNd5r+MOhwNGwDG+xnIuUeG1i
GFMo99UOhtXl6OUm6nlvKvz0J8REj59xOZ7X0xg7H1nYHCESMOtGc+qysz98B9LbTg5ptq5qu3ak
BYVAbr9iejC/TolV5+QKC2TFrvu8mSbswTLIPa9rlWfNcXnorQZZQGN+jew/N0979vBFUj6SBhE6
HCExlwlsowBZvBFq+La/Sg/aDYSwxzjceLcADIVSaL4w3v3PPbvB1LYSPdsv7IvcLhfRwmuEAAIK
kNRuZPKs0z7qZ8fEJpOmIgNrO1QwYGD4/mUBkevF7SoO8DU0c/RD8L2+ntveES+8hNomn89d7IUk
6OqH+DKqzR17L+g4q18dRkTFSGbje+TUJwyO1h/qnxLsSnsXxzKF3IfD8fEdg6SVwragjDwQHkaU
XlSnvH3L8BcUg5Gea7V04tpiQQt9tlp2iUAvIAH1H8kw3FGFJTKRJLmlnL9+heYGNScv/WrT+AM+
+sUFOanQUtsdylQptb87eIvksBuk8xhv+2vPKO4VCLHCjqK9H6HYDJk09XstiscDJ4DMqxRHYkCg
y+SCe1Hiphw9ZBZIAjqvERy/Aczyu/8vLMfNyMU6ZnQsXvkEQGg6wnzP/O9PHn/dq42EcNthpziQ
582a5duTB2s5AeRGBg+BYfAkJEKDHU2lWjSNB8YaIlqTN9Zx7ie0IWzCwCJTdpNRuGIr8dJbFQBa
F3N0xSuIj/vk4sZPHSZa3hOZKwKpQk7qhC14WkEbivdyGIFYZWtnIC5L+JtdEit1B7GLDlz036ee
DkS9ADQAIa8SJs3aBUI731cyLJj1/xdP+/97LQs2OclM79oRw0RnLB3jLnfnt8l+/JQMHms3HCoX
qheZZLSfnF/JsVD2Vdyg3sbkKszn2yWyBUlasNanJ6uawVYbexN5GTrqxhILgiZbkciSSyX6MSC6
8nxt/ZsT8sslWG47t6vhzY/mTDQJcXqo3OCSTmz92yJ1PPcz7EXz8y1KIw7Uvx5yOgQs92BT33ZM
Y8mOaXvv1Yov/0xHyF/H1wF+gGHmxvu7+B1zA22gzzQxRZ5PXRYWOC2+5bt3ncMsfaYa6Kj/RIvP
Nii12evsqdYOgOKSaFx6B1DhAflHkWvVCocbCgqxA9CpqsRvL9frClZftAp2mK6gbDpm/WCAAycR
op5mBlD/j3eH9MOk6XvZ859hKWzhuGFHPTXF593cz7Tu1HIY3ueVhqeUNDdN3baUy5/TDglMf9pL
nIw1JIvv713rKKXpEWVsYqrChh8jYmkWJ+WINDa/4yKoP2aAlhzy2dRc1qH7BFlBw3yFLX4zxUpS
EsPlf7CMB0ytUhas8Q27k4oPIfrFFUdK9mETm/eEXRto+XFysNO8WSl7v9VMHcBAc1PG1FeWMVCr
5BQW7hcVmAJR0T7ewhfz6rD7YfQtEXWonG0vFpoL4zNhhmHFHfIwxqM1WJV7BBe8i8IeYD9oz8Mf
uoU+ZuhVaQyRjZt2UFNaWXpI21tLNIbwzh/3zfowNac5EuUVibPwZyh6OUqmXUqez187HiwByzAq
uJT5tgWc9YQezJz5u9wSKJVFFFbHLyFw2n5I2grp35Bwula/oaoeqNbPzELGgbs3aQU4Nf5RFD68
TiftDOCxbmGhAbVh4KnUqi4d3GDlcjtJ+sW9hfFwDluBKxcI+levzcuyWC5K9hdIUDbVvIVk7Hyg
BFRkOdamsEXU7JUefK6rMmqQR2/QChO/EniDbb9aznrXVpM2/Vngw06DNUP+azJEQXjV6Nfkn+S9
EhjnIwlq+AlYAdQc6bO3r1BnMEnDcaqOGKVJZKez+uFw8Fws7j0whznUbt4o/wS4SDmxFnZf1ghH
ZNT9pBXIqVPql2W3mmg2odaL753xb8ro4QH5JuBGZfuX1ryR46/tsqEZL8dY/b6xIJL9TVBHoKm9
jFxmxUHCDHUUQj2mLbRBmjwT4A0dj+avLq0fKVTrjTwX6JwfcnQT5nAN5dGa+Y1F91QAVHdXRXOa
TqyR3f5UOqLfTEGSnNsV8XaFV2unNrcoH+yTu3a0lTZ0zPTVWwhMdduQuiTgV90fxJnC9zwdQNCn
CNGxVG3k+pdcRM1xCZonu+AwTAcBKYW7hHW0X40SLgu69sauIXz7pyGKhTMc8sHhrl9XJS6D3gcM
5d4YU2jWpB2ev09YwxdEMO2HbttExt4NLHuU1uYO8eFCxxqGFG6VQ9uZ5D8KLJnYXHg31ZMTtDzg
XtpBTm5/R9fKuvgv0dl2JPHL9fOyE1qd7B5k7ftqjirqKgCsMfJQ+cy9X5ZkPRJInMszIPEITHOr
TMybHVUiwOQRuVgfvCyz5u84iq0oWU4NMogmukQK1/K9vj96T1QZ+Sf77HbdpHV+5zLpkESAj/oS
9XBDlbPQgiGv1Qq1IkJVMxi+N4UZvSAGaLEf1oVHMeqNS3tJKLGNRMjtcv0/EKBB9hJdY3EKC/8C
0w7A005Daz0hIZQLkEITwl2wv2mQPz9lBoSPvLRtxkkxjQYpV9ln6GtNcG5uctyF+qaeiKxjDLV0
O6RjQvq4DjB3Fj8MK6Wz8dGHYiGHnI1Wbh92ocJmjJE5B1yEv0RNzR8zobdetHA5ofNmNSzVdrnV
u3pthCorOwO+HXDoJbgZpZ4oVF5WAJonUziRZkKq9aQonfXpZQQVbWsPhOzAS5QKmzwvGhWCIKoO
l7uomhXBl2WAnbuxa4wdrRw9GDqmEXqL0EdFWkZ45Ii0UJ2vpELIkQLFZ+roBiQ4YfchT+h/X0qV
FvPePkedmw3vque2hYXkltVrKApGZfyp2Iwhfy3kbk0a1Y+5LKKT7n+81fSM0cVkvmNSReppML0H
EiF+2RXCh8p2GhQUnWRouRoniaEH9BeF+HkwerF+HnKEvcgfQ+EhVZdwq4If3RRGc3l9kp7gfaNT
TDUhPyiatJ1Vua22acy7h0eFXAlv8iKQBUkLOqYULnXGINNY3Sw0MOBMTYxYcGlRfoBQDIbEOmpJ
aJT3BJeM30TzkNNCmPKnIu5OlWX9oo+aNO9jhzLdT3ZztP/NvgZL8/QFs1GoZnri27675D0cdn8L
fD+Y2Y7tEA43dvdVzi8KIblO/BGIUnm/ifJYruWta2orpX1NFJdw44ovlWW7p0LImj/x850Nkl0B
F6MtMy3z4jnuaiAdk+WefbmYIH3/ZRUVW+hjtvlLJPRT9S0LUGtV2H+3v8qpURWVRc7iZvcdeZ5j
7T1Wj9TZaL5l3GbH/RfpMowqbBwvcyZ7h4rji8xT45f2qMPAtaGw6NV0v4z5mt+x3XWYc2YZNaoj
ObcUbzAQckFS/rpInd691XkLAnlnDpcmw1HGw+Fz9fKQ1znnymQ6LpckpSXe87kzIaA+NiSF5oUj
NROEB5/EoKgGqSVUqubFm6QLHMKOXmPyOOtYNTByHXV/obYj2hVyHTxk3veMyr76IOo8d4ZGohnj
gDMVq9jXS9F9sLgbHkdRUqVS1bnyFzGWsw5Wej/bzElnx1Pb2r9cTbtrpcWH7QvpdQTek8GdG2Yy
d/mKeb0CgwG7ryvcU800fZQqa3CJ2vDczoKNcLdqlmkrPwnnooeOhMxnW48d4I/5nMwbQNEtEHGi
3hllv6nLn2kmAevaKu9bfFT3gMW5ZkqQgklXfINyp6ARt85A/EwGQ9HeXo4OhvZ1PlBMQPxmhyE/
yMCbEOMC+h5A/kPuh6+aJAqMoeTOWEa9IoQU0kQJtcZNOXQ/vo0aHrrctl5pLGbYe9OzeREhQ96+
Iqfpl8FjsHqMQA3xu6ffmSjMCsJS3SV4iKnoQWuLby7myfTq4g/ByLb21QBfb8PPIM5TGH+4qUg6
2AIg3Z/MhjLMPqpulhbwpzJCzCHoLmfSZrD1Ye+PZLuBvjNygwmDv7D/7KXsvJ+an88xKMFmmr+I
xb70pYc3z+N/JtL2KfChdcrNocvHbF1UCvRqB7eto+eOBpEpUGh8WHUEqUOKLvgmj+Ox+JIP/8qG
OeHfSq4WpoyAvAl59CD0m8B8Cz75s1qKvqOIEAxcoXFTgOVV1s5zvUvYkRMgx6A39laEwnBTH1/o
Dxvq8e30qXCOZXPiBEmLHvZBLzvss0PW/1rYogSqvOSKx/lfpAyZFOqVqk7ZPu166FtUaVXwne6B
SDgtvce0zEWErVSjlKFDSN+nKMzZZ+ZyecLiKFMMPfDlDVdUB8ftQDq0+O5pniogaYVeZOhUvJHQ
2YXPzziaxsPO1mBcO1G6CJ67V8XINuMbrF8oXS7NkYhQixfjBzUQYpTX800/WpqaNGn54JOS+9fe
15rLTwjHgPwzXVE42m3HWIDe/3uGLeowZVv2dpajMGR7ubZHmOorvPzrXtD8sS1F7n09orxtx6dB
/60zeuhzb0smwSMiaTDRwvbWxFMAc0rwAkAEPN77lNWNshEGtgrVDngzBHKYkOgWUQ6dZBfh83HX
imL2ohp6RKUhNsTs/aevg3/qfatk3YZgVE/BL/UjEcWMU0NcsNEZLIul3awU8us/zBcLOYtFHED6
RG/xKzTtoTFhRH3e0WGyFvkXhmIldt+ZpIZDOg5kPhJdL3ned3HwXqriAQBRcIGsyQDjqloXFABX
wK/2QF4g1nRQZuAGJEh+umPh3o3Y0O7YzC7ggj4zJkklY4gR8nCKAqxj/fJ2y2U3Ph3aRELzFfLo
xgGq12Gz57WMpzu5S1KauOv3jQ90bN1YAJ9gCuRqpnAU0/NkVmhqvv/RF2+ujJWIgpXtVwFLEQqd
4pUR2YC79twSKY793e8FXzD5WMWw05oWP6Dl4MVbLqB0qdS7mNqAqWLEIkTRmd2hbD3LZW/HAN9O
h6bzfMo2Ys72M6A4uERDsw2jc0NTKT/ZtiiG4E7nrMlImAAmV6h69SSvPORCA7ngO6z0vGrqiNW8
1BrdPJ+Yzt84AiDE71DZjOhowd5WWTZ9FJh1FtxxcmkafOFzvT4mobCJwN+uAf8wROr9L1GbOJgK
wbbIPo8Mh2erYjwWuhGhhFGdEr9fs5NCIFRcykzgebavkDZ8W1bwBW1rhOWBtFSp4MONUZEgin40
HWV1uprPu+DBto7eqK+7LFJM/gtDqmwJOWMwYkSx1XWcMXuOWN+6MrV3hJGrVftwBBq3dYFGAoTi
b8Rcw8pnna7EWIbr07aeVGU82Rx/3WlbilticHoXWY2oMdcOatzocoJlxUtRWhGRIlbRGL5MA6BU
f71lWeWpblC6AQ5nWfl9Z8unSv3sXDdUuHQw4pCdAP86TIJP4PM/oZ76wOIdHUtnzjCbDKEmmq5E
sRAYFZ3fL7ctCzbksGzbS7pl05gV85wPa6rF/cug3bpvnfMBmQq9lSHbNCuINHYn1Uu2jQMKr1Yp
5pvtW3dCOUu+hK90q35voYiyKoVgmE74aARVY/1JIeh90XuH+zlc/DIEY/DI5wLdb1P/Tk4tUb17
0utZkp47Tkl0sJrGY50QquCcSiHnuJcQ4C32c8TX+L+kAMtdoylnoJKt85smCpabVN5q77ND+lF/
ONaEdA+mK0RnTDzRG8E9x7pG+YnRYubkd/MQzUhbCDU40iGxmQMEYInLRxngHBEsRHNkkSzwJ8dN
u929yLjD/uMD0hVv0JNGpYfJ+m588ucIwcqtCZOyYJ/kC5bmQOgHRQWDx2IR1ndHOwswxTqWeLXz
v/gFLOMIPr3xe3Ms+2REQwaXp65e0nQpwt8yJFopYlRwShp6T/c4dDunf8EUnk425axhZ7f+CNTQ
Yq59mI2MfVYFVZ57I4V3Pz/MhNL0xURzMDiHMuIkBFROXP50kkVlzSh9cwnDGhzn3aVuYla2ppOd
D1NXI0ocILj5yUq7u1M9w4a5xLIlPJIYUdfzTRsGVvLZIdgMNhefXZzZBrsqY37ln6rvNu0e0zDq
aB6A9jRdliOwKgMdmvR0/4oJHZzi+liEzqG4kcV9C/4rswCdWFrdh4WCKypcpIjklAuRP5omAgbG
lgc26tV9tWVDG9EaH7Fr+SoyLV/PnkBUZJkSzqo2ryjV788IlZIVN3SRZoxt0sa/IaIZG6r9tvEx
Q0kM6cx7uq5CkO2NuzjkL+AO9+w2W9TCOq7YsBVFrqsCPguUUSC1rG1ExddW1a4QYQaVK1vcbYUP
OdUCThCMZ7mLyM1jlaXZOqI5rK5cabj8FKkE/cSTmF4lUIUhYBnhXoqZz8/R/Sxn/Ss+7XnzWqaO
6dJgXwqj2+SSO9U0oxFXaXf/aGXinEarRiT0+il5ydmfSxOPO+IyAuPNSH09hBsEekyASIZ9vNbv
blyMQbbcvymRkn2felFNjrJpp+PymNDUpGnroDEFXbGfICe/pxRqWWcpqJboODi11unA7N0RheRq
oAdspidxKGmZw86PPkheDYkbv26W4v8RDu/+zgr7Dhp96lhe5KgsTM2SiK10P5ib3Tuo0SJ7otOZ
KPbzCLOKP39K+hQWGTI7gMkbNVTmTZAb1qRbTA03SuJi1cUYOhEK+rMnxtjqtzGfKGW/faQSVE27
Yfj6BZUXebtD/bv20bbrU7bWsxsTEBmdl7rcHImGg4aeCYBXoT2UnQrJTgHKC8my9Dni2lCOAs6p
wV1J67/bmLJSpkVdagmhsYB5pgh+QrDKDfZYxzLetB/AZ1q6pjOc5nWoksvVT/SZ5wZkRXu/QDcY
5BanHd2JU2RBrEVsnndnC/dsLdIUDDvs0dRfA3rDd9ZYtzCk2LAACObLBTPR5UI+FbKoKxuphP+i
bSJ1M47R5GybhfhiXMRUcdxUMwTIreaKxqJNO6P8H5Vac6cPiXrE7Pl6AG/ruwBAnrANoL/aQBI+
dcA/ZiTuxlC2j2/d+PsJgxlEcx0AOxDy8bDHRS5PLND802kWJXD0uamNRSNdtGSlHiv9IUTyjDTx
wfbTtefyXgrtDg7rK7G0xVuA4A7SRsLacCEev1nSCWrAqk35ZKvxAU/UWzhAKvnQ7yGUOnnq0jlw
f3WxNg/U+KrucQvZMhF/aL7FXe+9+tBfvtTgap9mWBnE2dI6LFsK9EiY2OgBhhfXuA+u6P28p23Z
JUMggrMFa5URujPBwJ+imM6jM1RSGOKNwyd9Bvyv6Sk7Doh+ri5D11Fuyrb6D5cZqJCKiC4jqAT2
b9z7wfM+xLtpF0ZX8mYzUMQ2catq7raRtX3Ans8rUE0vD7YSBjtFIuMZRaHpe/4E5xva8VJUrbju
ftHOtZTcwpNfc827wmPiuRItff8rfEvOEOwvkXA9jf6Rq6A9Hu2zvfLG6GFl/Q/FrwtUJ7sayRie
hGUhy3RCwa/lWZ5kf584Oaae+HIj8pXdqYsNRQlbeOv3VCVbDTtDncTzLW8a+HSNcr+dMX65w+lI
WlTtXOc1Ov8QfWtFi+7vzmNGTjh+TpnmiNPPDKtGlXId7TKlXBsjdpOlDBcHpyo3u+2O4GYS79T6
5b9UjXtHxi/DxwIMdgNXZizLVGgsM0nCzg9fdUAJHsIfDUMDmTC2U/pS3getus5p9J/w34O9Ncpg
iwDZEMa0UjkkUTOR0mQ/jRuXGBlRFBRIk6jM82hjurtLvFMsUpFu0yAnnvQPgkdJdhEu3Puf1Yrf
6Vadd1riEt8pi4crUKr6bAbxxjJi1D4ra07py3dTrivq/73dJBZtXB9W3NveM2sUrXEl6BwDz1pI
5zYNZYCWZc8G1nwMz4lXb3NddL43EUbbBu0f36AUyfZqkrIEheKbjxgdcWfX3QJhX1OYOKC7dyML
l4q4YXdQX6DjIe85XUN86AUPJVNGu8rKUffgjkt35IytoN38yUPDQJq/VDH1lTwolK58WNBq3Hka
q4xfNGxKCqMW2X7BKBZHjt2+nEsZyvkoLTa9tZWamVHKbUsQH9BQAk/EhEai8OAXqtbaaWTR6tmz
FoZ7GhV2w0qdyD7mhuw6Lh2DRnnNbqwPz7tue/JBCO1J3G27I25FygwK44wSxvfrv5mXOAg5SsIC
xfAaKOMBhFxOSi/xd+Rf21Uvz6ap+ElX0njlX0tCJMyVF9wmcBPX8hNpKlarSoPd2o+4XB0tzGkt
y+g3EQx+J0ICygwm052YwFJk9SZZvksOqjvz1W7cYXCjBb28DZTgbqg1Wd16jK8XOt1I31lRagxn
t1D6Fkq9lCkaO41ES4fbBxqu8VTFtaGKowz53/haBCHPoruTqrbFUEawmLXDmG0DYPYC131ij3VC
H9Yi5NDOAuJDHvk8cMh9qb8b24nHrXgAS4nW7lP16Jx1dAmjivABd7lWDQ1ZmfUlM78pmWYh5hl9
4BHFzYLIQ+8Q3IOU9K6cZpFvVV7poPxerXyqorUGZEur8tcAnGyM3Of06R8atO9A3eGg5j1I2lX3
1CXzs2d74071N4h7su/IqrxkRvmy9BUXAdyF7b7qKMFyoynhqa7wmik0CbIGGAyjIGEfb9LTaV7L
QEPn7mY2MsLUAsvgk0+o9epvFcRIrZyo6TDFLSfIUJr2HwALvpaUkQ8gxPTQuiYUorY8/oboWzJr
dOrG8I3fSywxMstvkWqLM/8wQPsVbYMSENWE12oTBFKK5KiO7q6GPUpD3yPBaxdBTsUiF6c0h9ns
ENS83LEXKkh+1Ljurqf+nlpzIHGQCep9pD9BzCy/vidZWXD35XgAYveKO1xgUJip639yZ/06MnNu
dXYe5Gni1U/Z9i0PBG/MWjOaZaOoKICZBMKusrZiAJkQt063L/v8G+fx90KOd3hGCIywJwNXcBrR
LiIArbqYp3W6n3pMoqsINqXWU5/uwBoxQOkmKnqyMWNEwCLqxetOqWB17L13Cqp4tqy9FcTvR0xw
0Z10eS9wkh98ScqZf2pGkfScr6E2tpemXMoSub/IOL0GvcRj08/bDfthreb3g7fwin4Jnvf9zNZN
4thyqjMzqr+c8kqaEj/Erv9mmwY8h1b37Smk0BOYrF3WbOXUt9oNt0ijJsEQpfXvLH5Y+EqMm4ov
vvqnz70YBPDAI5Xf7dqNsJy1qDuve6+yIy2qJKJDlR+QRm8aXpXYj4hxgGk4e3Lkn0nMjqXfS3ro
7p0LiAuycSFzSCRX4zZGR1J4Tuo2A93smZxaudWtUP5D2e3hWi2U5BktfyUXgXxifgxpdDjL7bZU
qP/QnOF3Seo1CxFJX+iTvYV5HUvTE8edHBquz40dagSZgNVpAJ6at+1z2YnrfojW2NKI2amqeKQ/
PEMg7K084rD4pW00OFh2YbDdH9XJXrpHBjRP36LCHNbYOtbgy/WLrayOX9Er0hKmv4PMO9Im+dnH
PXONuSSUfqKzH/YlvQ55Tpy/IXMHTGS/M6kwEs3D5Dw8ZkpBSVIzmn74Xj0omPZpKBGGjdBRMNG+
0gMkE5BZlzt6jKBpP9LOM6ZvrbOQ+bfLoYfigq00029nlSEFe/XVMUlBVae2gbkAPKdMlv1s5FFh
s0X9zq+BKSs+/TW0PK1dFHm35hQMau8fSYBFeHwhMj2c+nB6Xu1uOzmKoLae8kGdZXJwlV6QjuJU
Kq8Fy3iz1YCymBRMM5/yYK9zGn+FQjMHBnLf9f79nXeImPeZc9SHRaa6pK4p6x58SRAKCzeSD84U
EEFUtzN8jdXofclESvv/Z/jHWEVLHvuT33BPwZfgWTJ8ecGYC7U0pYiEEZ//n8/PaPnFHR1578+d
AkbcNci0SZIlfqSdtxhUebCB/vb8OSblbseNGKh8GrNWSR5N9cXsJZ9s7Ws2jINgXB64RkozfDV9
g05HQpcRaihnxEmdHeCadDxL5DPLBUc28VodzBDP4l/+gPAoqPxRKZ5+Dm+yEbK/UbDqnxoFHycd
mUwHs/NyrpQ5yO5E/YXNCokLdCJWxghLzb1ZcACglJ96QI/KKr5W/zzqgXqd7DK7VGiEQuxM48BR
BFgMv3xrY52InL2sLxIZGCFbRkf0u9bI1vvlVmScyU8SlVycbPudhYIdTZSnTOS7IifzJIJyhMQc
x6IP/zB6BGiqOOKQSTRJkYEGdMbUSorsq6b6KtO+C4bG+LWIsRaKWnUynPIOOwFr51AGWINrasjw
qXuF20Qa52snBBTKx69CnFvy93b2N2aobe/ZgZdZxo5ppdDGCyAlLgsb0JrBl4whsaZMndCWTQEv
nDnz2cWnvuMTnMbWhFd8rOjIr62Rg3EMtdryWb44nW6tnhpIoNBO/Bawdqas4aPQFIrt0AYm6B+1
ssgw00ISWbvhTvqhvxS0Qh3eX1tBFmFe90QLx8lfcE/FjKBR4rt2UbE2BTp/whsVK7S8D7k6DBIf
TijGnswRUOTXUka4i2W2lpKo75YUEe+jZGX7D0Qks82YXeCNH8q9f/Agm6RG/KvqRtPZCRawsQn5
wqJGnUbdCCWQXWhnQ7egS8XepEU2F0uzXuSfrCL1oPMlRnKSt+yksbwaVdU26G/CAIdImianjlNH
fSEQ6LWUjkiUH6/MDk6U0RiB7K03hpZhgYxt4T9zuq1egjYyz1kL4rfWyQboldKn8LQZT126RJLV
/jezxPVRfYbj1mBspmSxbA3gdh4h0cRndSIgvE6NVTJftyg8Ss5P5MlwnOD1PRODkXJDCik/bCPY
HCd73RWZTSKj/Hs3GvTF9pH07QaAOCwKlrIHKYpLrS3UcEM6dcRGK7gT935sHmLH6TDv9vb6VhkU
FwQh9Lu1XT96k4iSJlmD+1XS/6vsq8PrgKDOwhLIrOpaoV3FLfi2lBD7H2SErZdOPES7N5ZlYjfb
Evk5KUKWnOycdaNrpixnhLyfKfDtWbhXr6tM+gVi/BpYM148uqk4sDqm+yZAUw+bjBRDbFGQTyX0
1N7NWf029x7VrGylIzLHJJJZMamy3yuwqYplU3gURiv4lbwjch096sdsHjs+t6mak7kwOs2Xyc+p
WUdjUBnsWMvKtIqll0ST0j0RNZZzWRaQAx9/Ssk4I4HL0SZQ3P607F6dqWXIyALYgmljmRNWib7b
xXIhmNyCybX4k5qzN/KSrWl8dATfB3KEvgBPhru9wOvw9bbr6c2dH/Z19hgtnT46fXC5UxyL9f71
HV4LLJX8+gv8FKE3HmkG2+h+8PRzz8h4WWFW3k2JZ/BaE0nNKDxP6zZWDzr8dNfTakAaXBH7TwK0
p3ho0T5xAn4sCaHG4DWZpP96GuOsMWC1MfW0SyeTB9ckg5/4iH7g6aSouui5IqfQZWHluEdx0Y6N
e1DjX05I713sFloqY7KeAOO2rewriALE7X93S9ZPPHB0WrD2u1a5fa/4IJ9nIVIWp1DHULNz9Xpo
X3a1KYk30pvRMfrG5LsfcjJgsEp1p9WECD/f0O68Hbk6E+G2uafAPY0i1TEP/nt2vSjRj2D2x1Xw
2mfhLVJ0CDmeqpR0ef+STpdo3lLnIY9OiNgxa6jkhacmsDqAN1VKPO+jIUrPJaFvsUsujhPz0vSo
6HgGUA/Czf9soAl/EIY82JLY9GZb1RijStkgAXdP0IxyKbNRaMKlj6lx5JO+jy5wqd7aOVbqhFWh
6QlAhMw/ooNgDvebw1rFvlYopCS8WfqhOGqPRsZ6C8vGQJWa7uxPCjnBGlKYPMSPBEx2C3vrIrrY
M57qwbIbBPwTLYkajNo6fqqsB7hzjQhXMtiWSNir9hwQr7QAKsPDLlRlfPOCyluW7WFn97v5FkcL
cFX3nVpLdwSi1CkS2GdaX+Zk3ncYM8dJJlPFRWZ9bNF3tnPfW6LtAuMzAl6x9Sgrd81HzqZ+fIHq
YG7JE/viLjRRPY0wVxyCQGtlANRPXO3Oty1sP7925sIp4Ks2yx4z7YFRk0f6Q/PF5j92yUJpN/nW
bdyAY4u3mqcyoXEBZbnPsVqmXBEEdP/2TbQuNeLy5mNMCPNPVbp29lwKrqXv1BElJBgDiXEFGhck
sPwC4nLV4F4PeCX7vj1TomS5lq7x9rK39zQYXd2dy9rVYLG5Hp342llBMIqtnVogQU4gXeo/uG0K
6jK2G5LNBao7bkTrdhJSM9QSQbUyqoZnuqlU8mCFLeD0+tFo0rzNHe5qmf2eqIter/o6KowHArFY
qhIBEJTNQ7WAUBL/yf7HzBxYnirnaEYjDVRlnWvCfB9uM5FaAju/RzsZ6nTy7kcF8tWTAD1bJOHg
XMZ+WYaXkVsjHsh4JnE6gkJo2PAqR69epnFWHK668pvUeLAK6K+CI69YLNvkKpSCffUc3VQ7WZKk
vjYmzzb8ku2Zt1nhTnleZPSl+a3PZ6EM+tmm1PxtreSXKRRJ6iHQWzDnFVpEaOMl53Nq6wh58tK6
+37DBV0FVfvIx8pwTTMCjzBJoEJmbMFGs9ijZGrANiS6U5GXQd28HwPkYzrrgn/L4wTOCjAQfXqB
Zr02YiJxyeY8JdvawdhIvLuP2KRi2MV9+XXRV0UU1P4L0Z/yNo68b7GZJjSMUeKL1D5uAEv4pmzZ
cV6H3Tgf3PVkciVYJw7APbp0/uHyRK5/FVx/LG4D4g9XHhkt+CMdgv0RghWRinC7EPVhsYJbbH1W
VX1fPj7KwVdlHEldBP+eP+4RAn5VVWeM9i0KlSu6GASrzJLIBMlbRv1R8C0xrAh3lmYW3AvqMm+X
f2PuLfbtkg0yh7vYCcAN2yq7vd+OqUjNSf+Nnj0WfQTRCO+szQgvmqKdEk6e/1hLZXZQWXAfWF3T
7kK3d+oy0mf+RjUDrYf7jPhRafK6zeTzHe0TMwOQaDHsseOc35tQ4xExtjk+KRSY9N3OZxyclx4s
+Nld82zuk2f9PNSl4E8ZxmoH1r3unyj/t47EIl4357Tx7x0X9kR2PQTVybLcTrWQD5MmTV12EE8A
WOERolKJZP5fwFBJCsi5vgOzjtuxzoDuX19OEyhdSkaRWyCkZo8Br5hcF7HZhCBiVumRpO6U6M5m
g7bWSwjW4ivp2zRCHqc9e6tA/t0TLKb4R/1YPkSb4aP6hgIjyTVcU9N6vjGBlp6otlqIPMC9O0+x
83jlCs8zteDCtVvK/+utAyU9LpcerZA3OHKOnlEwTjqbB6N7eNdC7RfpEJAO/EUN2EW2FnmAAcw1
RtkIPtTbuhgZ6+Cl3d6XOaFJ7GP6m3GgVtM8Akr4Tbtj6rrJxP+QPcI8e5lo2kccJvNMxVR/aacW
x1OOhsM/EADQ+Q0O8/hrZ4i4weyjXGUXmByKVoAW5AExXKb11X3CFYl5UbIHuvT7eymR/V+CuoLG
1SFW8EFa4ITZrzzoMZ2WC9KedlC4/GA6D+TwSFPshCPY9KcNaZ7dUlUQIMUJR6SlYUantZIjosHD
VGyqgSYseIpH4U79xFGBB6TjNUNmdc9TQapNTtMiyxsl7XV0X77B6LWLu2PdsLB0fcwxfCoaKB5A
VCydqNp5KlARNKg2CDjrBmodtkI8PNZt71UCJSuJ0MEvjgHGa5R+yecm/eBmgzdGsFAO9wJ9NqjL
gYyaoXgb5KJ/wwxcUzRS8pK6yuof3fho1/C/H4QT1nBXtWXAYgprMc/HFtRHYujVOHVBhBUBpnOS
nhw5gM+ly964E8IDsTw//aHakt9z1GRndYInYalVAxIg6g1i8fzjJoWUDQw69C2FGhHp/7Tphoxl
YUbdM33bn9JcORPCOwB+I+WK66vHMsc17BHvXe4fuZwXBNFObORYj1xaYLiGyCmodm14Q5ywENC0
IUxoHbb7+JV8LwEBmLHMR7qQBpZ8qjOZA6SPGro954AKvZklcAO0p/CNiNQh3ylrffqhOOKNQw0I
jSOi3bf9Le60m+OGnr4F+TE5y3ERb5bfZ455dQrNJPq7huQkMxtqYbum1Z23FJtp2uhWo5yNpPc1
ACIRuR5IbXHofUtRFAZaayT7arT7pEtSV0j8vZcgxFTdibESvobqp6XBStM+v8DSuSTtAHZ772MF
J17LOpRC2B9dJxJ3ASwP9veZx6EH0ioM3yLlMWZBGLJyErTvV8Cp3RlprkVXJRQKmDeKqp37DVez
JLIbsLkXKsP0Nuzq5wqcSGqUw1AVdslZp/E6Futoj9/VYhJMeT9lwIXoLdJcM/RsAHX9djjPfNA8
whsCTw0Xyfsc+R4HDZOsWdMKwHiyuwQOw5ov2QLwColQg6tkjL/+5+1u5ysowAy/0PZbPYg2z3Rk
Aph+VSSEiJrS1COaqYykNLlRyVqtjHwBm3C+t7bfQFua2krVzYUOI+S+H9BvAG/jK5A1xjIWKIsE
VcKGyfTDzqnXIO2jDbteyK/3JNgWN+5wHVq3KVl/rJPJ76da1iOWpkzWRem2P9LxXBpQu7xP4Kxh
DFPOx2+szjH7ZyudAfYsQ8I18jrB7C4sIAR8RZjoyaaQDCUMapv2h5xZv2ty7pkaooFOSpjk6PMQ
EQxPfzyXnH5KDSnyFBASN7ZRyvwmVWkbuhZnQyj51qRsj//283AoR50v1HCG3mNs3wU6+JKAgl8q
Ya5xpwZ4GeIv0Zc9E2tqCDd7QI1FFy+HkEnevAnsAJxJ/xMN2h7qQciT+oY3RoAExWySbdiw9cSe
MA6pruICpzieHjjcSlsdDUAix8re+8YRU7OCOHjK8sFWbHlX4Q6yLCJnT+QQwqdojwc5aS/6ZhXs
CxKwWl69w7UGzBMhhPrBAiHSKXQAQHlP6Yj/GkQOReuzcCMOpHMVCXcGnWV/KPuWtasJKQGB3M41
+3CcUncm7EZ0WaFUS03maVwoitbK+q2zhJ9oS4n3pJ0at9nGjYA2XjKCQrFmgMQ66e/hVl0YyUVY
wSO20MybQwc4Ul0hHOIR3Ue/87CwxdYrPStto2zkVUvP6E1RcDP1FwqLln0rzm/jThch9F0Scefj
naFBrc2Lk2lgHy0uz2yW+YftNt0tx96xx65qKVubC8GtFnnoL5rH+PQccL7jyumBEYNxWMeohNYc
bhyhBEFUtvZBdnOBKwaEN18/taLWl8dBIxBcXg+djN1tCUw3dyk2J90Vz8itiPBUT6+34vmgwdRE
8QVN6NloaBBd9ia9QgyPzf0y9o94O5fDIw30oc06T23QXvwavhqjEqkun49jLCgbPXO/fk+JAskM
3qHFCQkFvhrqup5621BRJ4+dhUOOWpXhiYm/sJ6DKh8QaVEQ1mvKwZoKbOjA9nT3Dh9uLGz9Y3C7
vZWFh0caPCKy4l/hxwhcjp4BvD6jxjpRSXa3/BVqJNqXQU0wZhxaAVjtKRYTnJs2ly1zIXDC2ZCU
lUWbGbDEZHpzXjrjcJQ1AC4gJDkZHXD7WUwEqOJdgkcYBFqmSL7YYy4P5838EKJMZcy143IcXsUp
zZIKqfeT7YNyHE469Bwi45XslKkvNbH9Q/tRxURAbbLD+p3KiZXY7Ma/2tcLKESBUyP7Vvn95kV1
Kjte8X9tqMT6cepEFocnGmChqUtFD/k/fZAbd64i7i4SGlfz2w61zxIJhC4Bw5U24mmktMK2j1mB
tmsBXpp4OFrK39vjr6Fhbt71AO+VCoKTy40cTEPZR9lralLcpz2W2IajeZGneuUSnNtwtCieAdTT
jdeue4xYf2N7bzM6zZmU/fi1qKVHdrgVK/DVPd2Qseg7CKsITXESgmeic0HeT7figbFBpIV9VDX3
WwvSUpJjln5+dwhjPiIlQdyKj30jsN2kKW0Q2ZStegHwg8/2U3tNV3MB1l314qxRAsghMQRCcbsU
Gd6A0QtyOnpkbGZNnXd5k4DqTnZvtiio8zJ6FWQtAF9CNqIPm79TAAiL/UGX4+gNU5jVKuq7Jrbl
9nbSeSTc3zxuo3POeLwbt2hysvhjTNEAUuh6Yf59HQuctQZxGuZFoMlOwnDHV6qbp3Iw+4A7tkuE
6CZ2riLpDSUEb5JWq8kkSYxbPwdw5wq6TPiARMdRgijr1c8v7x8Q0vdMsrn+rpqJ2MMYIuXoJCXx
krFyJH8Z3aNUMPvEoYcPHM2BTiaptP8LstWtAb9/oNXcd3Dd7q3M7+WctPsYgTzWlNxPBj4aEoPO
0MVnEwnSD2ixLH4MkPNyuvq/K/SS5s4dquoQhHd7i/e2KxbNL9PGOfexfHLkMkXwn4I4ONS8LsRa
nFoc/igWwtCOf9D2M4TlSBzX/QAl9hVXL0LGMiAi5dpsTGGTusI5S5uFIJm/7I1cJ9frk9+H/2uU
Q1SAABnQ2OaRzHAIUd6grb4AP++eH00YaziGjpadkMUFQue2p20OM/3/tr3oySPylrhlhEDaz737
lRFoz1sRCkmLb91uClD5Qot5f54Fkdz+L/aerjpQJ1oXmDwZy3kTiJadc98vwdrWl7/19FehcfN6
ECN3ASWtXu5xn5gDaKDrj6xIeJFSgvpJbFKlNH5/NFzVB2FC810d8+cVzMcfoJn2wCSqLsl+sMzt
4esC0LK9yCg0fLzn7OoKivlXv/RycdgGRKbe16bjDzCv0wGVJRwpout3QaH5yfuIUHzYNuXMm+86
2xydLsWt3rOSxKYW99UTe7xn02ALyajASZuWd9PG1Kumivj5lQKa04d90YLa9eMpmbHekitLcHtk
EIVhOkz89KN6ga/KR32dtG8/VVVHU/vIylULiAxvwrgfzCh+8L0Ax6Q7JlSjy9nuPnuBDtoDYd65
FfmiDIK5HK7kfvcpJWclQ87/sU4WLCMuj+XiR74kaCuGU1/gCkUS0toucGw9PGemiK+BQU8TgxSr
uRXcEGQe/pmy52oF8LBadk75i3TuoOPK192VfSztUAgCLFrg9A/j8RjMiW7phNLs4yZsBcXhXiCl
Udq2YlDe57fI9MO3+8049SbXd+G4UmSfjCMBD8axrQRIvt25zUOJfpfYCdoTOyHzi5DBpfK/2RSU
KbVfdEnwRC4y4cqnCD0Wn8ayezKqJg/OU8tB54rT7DS3jBANydENwIMqXuJI+NgHOBqSUaossFX8
N/+zYKx4SL1bn2Q0ZJREjXQYGz7Q4dVtTUDINg8BaqP3ZjkQPjDCmhkqmGK0YAzQK36HTVACnGMf
ygwOZ6tIzRbz2p0D02i96471bJfFjHoPylaR/V3gsWzvXf67Qt2Q5WfQSisAfXD/D+mwTc5EwOLT
oZxrI+prA5sCObpZzC6K7hcCWyd856pgtluph2hrWQh83Ot8rhcnBHX9WSeYFeW7hEk1JdIHu+OT
zHBNfeed3SXUJHVp1Rb0Jj9bDQIFdwZcMxhGl86vOMbbpEcVDvGFD7+bymXo6GZxPOrz9JAGi7zY
KaJBVY25g7oPUxaAgip0a8gMiKyKNvVZ0dfDXFgEVpMC3Qebc/lsRfwqfKCwthIJRHc9Xoz9n+/6
1gJ3+ln3ceGvHids1oTeQxpnqprqU8bQOSBXHht2CdPUVLL4o/pJ2/wOdScGE8eWfzZELtRcD8xH
YCaIci3HfiNomhpffP1O+ptdxMgiYBQ7My8dRlgBFzKwFIevOwqKUG/gXueVuRPcAlZMFQjO22jI
jYn0ggKOJhBcQJ2yUcEtdMXj5RxIqhqXl/GJH0B+3ni3utmAZfpWma6PG3PAd8ZciyfCzqwgCwK7
A5dTG9hZved01MSqdG/xhYkXet1kg8VjPnXAvjZG+DrgW/eVyDHZifwSbwwkbTHHGmpNsa9UKBgK
VGugzCAhsGWIRCJBuGq7pdB5tB6Z6heS+DeYl95B7iXLmp9hOTlpF+iw8p/teUHaKBcV/q+rBKvX
F9b052afPEdUTcgkbXWnMY287pr4EFg15LW1TMkI30wpVstc1rMmZ8t4BPYhKzVktj1Q1HdYsaYI
laHBv9DkMSIlCndi3cteHJZmbPz7diMIVAlHORngzX+DeFzyznwwBfJDaPIxmlVi4T/+33QL5t71
7iwqaRXX3/r87tDG8rKDv7Ur0rCOhq4s25WFTe85+2vyBr0Q3i6LpL8gIKuLRCbKy37THvTa4TIw
iQv5hFWd/LS/QCCu8pOaYATdreF/rVup1LVaSFlvFPSLCXdmbM+MlAST2Z8ybXfJUxb9KiMeaC7x
+79zkj2rAAfaF4hVAzEGO5LMP+8gIna4YzoPYjDxt1M/nfTosqyvNPEjJE9pTm72Mj91SI6b605+
keQKyTgl1qd7veMVaho5MF37nsrx+guWLqFJ7Z+NsgLKyozy3v7sa1/tYlsMnC4U8nVr4+VjRK4+
2MsAlPJDcKPtr4L6jemNTcldLrK4pv7VECZ2vfZTcH1KHsSjOgiIRJPIDwsD1KyDauigy8ZdFlCc
Ec5Xz4j4BHXa6wXfuem4l0+Pn/+hrOeXubJMJuSZEKYMpPEYC2d6H3yZKbx0ADWx9ksUmi3yfhJW
8p16NT9yXKmRJ3jKBrocasVQdjr2GXs2IXkEuTk3KYgsQ/uQx0mYplW6RkzRteMTq9p1EQh+Q8ty
fIOENZTYfzsQPLsgf73MhEHPgJZ6Ld9oB9AnVXOwzG2ssRoBGOFZnDRbOJnPlj5wgCgBfZZCR1Cy
ZAVgBzhsVQgkh+tLWMnQdPIWLQN0B6EukrqjA1MDuWDkQJJVoiRnKyaE6qzEB4PrzT5dxjE1DY1X
BYCTOMFHUyDuxBRC6F7HX+skbUIuY6rvrLSxK2043vRh4k8YQMUlXBWuvV+TA7hc3YMQWqIVBtT1
rfACzjjyfb2GYq6KCMIwVOZ79XWqWmY1ETfgSGQ2+3kB3rxLf/FJFxpkkQi20urmFDfkAZwhU6EE
nRvP/BqFrBV9XmCK5YLMXQTY2Knf0IcixGwnrnYrZ4K5nwmOlIEHOSSbxdv/rRHytUhUOFvqKiIF
5/c9i4e12N6mvI8MzGCu+A5T4DBXkxr5iCUD8jM+8iiL9cPodxNxp9dTf05cugIRVWm/OPklfyFm
j98G7BJ/kAYmVRjp4j71CJ5zptm5xi4369mbauAoRKpkOACP1cHgXEUNOxB5OetoNI8vuBHQZLwE
7YEjpf7KPfHHKNW/TK+alBDp6+O33Dw5yzQpglczoIvBD0i8qcqtVaeCAJi76SnW6HWIqLGVJJq6
CvWyPXA3SSauJIZ2+BPvp1C/zdSMhMB9YIhB7XzTFMcgdxR25UCTZUeX2UB3Ig18EzJWHpzzpEG9
G9ywbk++Gu2/755W+lJYg/TqrKsZEzy6yLF9gK9MVNIh/lWJLb/cWlODeK1f79zSBaYNzRKBxzgV
BwbWKNUm9q9zxMGwtBamJFEPSYiv/vf8PnZLZJacZVboHPSlFzO0Xj+hgMswvWvsgEG+ITqwVFgx
CCzFWiR0RTXHZKPEv4FzgWjZNql0EP90TKV9LGRJueWRJNqsXnSf/tZGvpK4lER//VIcGMG61Mk7
CwJ73Mg8KjnKRKead/pFXTqC9hcLsPfu0HJQfvfKolNrAOiEFBKeS9fChvr+gQOOQMIWz4gIMQkR
w1gioa+SPXyTbzRmqCGTl0mvp8m4LY29qHTsN3VbcuW9xuSHLFRxdIjtg1q4J7+L8RqyEcpC8NS/
lgGr3CQejjfriznQdNhQmoOYKf7Uw5mB/xmSlMMr7hx+9XoMGCfcdNpaaggKzLiik25m8AMcQ/89
cTSe5cDeV4NnzzF5rX0hU0V6r7Odv8PmMhWKrbzRzTMg2DWJ2tbSMQmjNuapYW+UKnpmnlWEt0n5
qKV4tQt/ouieObI+58KwlWxn/lS6APdBGOre/z+FBsa4joITWINQg9ZMREEYYeM6r6pGuFQS+7c6
YzznDzZY7vIJRYFB4phi+xcwahYBkXOGZTuFGnOiwk/Ebi3vNHrehiF+doWZEfRVuVHl58qD0Lkf
YaPfyZl/mQ+HjrmhP/UJkXogKSeMrpOCe0fsC6rqliOzzacaCGEV0fASFhPGV0zcV8crr7YhwX63
T/7+KgwHXH3tvuiVNMnNwhX5iXUUnvNjmgNyeVpdEXEgPF1BEKB+MLk69Hurl3Z956wa9g0h9iVy
sqxAsJKknS5xxqnORYF+q66Ln6F1gf0RDRUWSwkFyz0hlW17gGlFA8Q58X6D0/zbzAVpq/cGvnBE
n1sBW9tDfHGE9+CvLdsGf93xPuLDg2Gsg8F90eklc/75Pah8Kh9BIaTgQp/yD5dtCHXbvhR1ZMfm
ZJR2OQORSTml/2I3dGqMhCSwuIvGHpoRQQ8Qy7zCtJrVFbvR9Ikp7wuU7tyxen1ZOT1z+lJkpJop
pV8SzIzcHhE6BAgdPmlDoa+Stsm+cguOXFkYozs2wavPLzm2x4hLW0YiL7Lz4DK2JimuDX64rkpL
/9I3Nu4/L395ZHMO2R2sRm2vHT+Iwbnlq1NEn1QEqNBcZIwujAdysfTvmH03HU2SCk5K7O2FgzUH
RsGGdkkris4Hvgx4eSI8PMgZmAOABAy8I78SMMpGMFiSiJHzqb1k6LwoYi6GfWC8pedxWac38XG9
qkGqTqs2v2HcEy+ZjOrU7rrtSclZxdOfZLC/ijt5LlXS9SD7BIEHttzeSsXcvv8zYWULTVLg9enO
gauJF87IYyTZJifYx7OrA77INTdvTXZfiWzFNU3b5g+Ish4gzyv5xeHlBQQMyyK5i/rw2+ni+uGK
fzpqo/d7K5ULpCm9NnREJb5DV3P1kxMQPjqJnGobRYfDgmFd8NerUF1+afngCaoytaEgVrL68OCN
XuZpRDHbtixogMZ64Qx0m0LDVzgrK2pytyBvukjM17EmhGp0hGvbYC6nmjitjkvSHYmTa9WDac5B
QcN3y0M5flxmSgjw18+QvoPTeZPH37AtYz/UV374Rq7yNBRyuK1kaUGNNpJ71d2xHvTOx89B+laQ
9uaTOvgULvAOSpuoV/g0slhz1ggJXxPkUMo8tE+prIKlVOmNuUACNbWs7/kD2AJtTipN/2UIVtBx
Q/LQzqhTqDvrZG4mnKDk8t7KlzcD744vb/4HCHcHcITkT8w+4MdD/XHY1/uh3YVfy2jBH6AddDsP
OlQidB4SY3gWEU+kXvfFJ6zleK8KJ3+VRvF49uxfLR3vP9nCwFMpFqdi9qXXlVdt/ykNXDZ6qBB0
kO1+XOmZQYsDEfjIjutoM61+fPc+faXY3V4gHimGSZwCqsB5caShoVlfmud625xouQX0S4+mr5ly
ZXpgKw+Vnmwg6vC22SwJem19isQrZvVDJQLfTLklrVQK765UFEZpL+EW/GM4SHAHH/tSGvOBI6ps
Ujo/fLBr5ijndKfgbPmgkDOTLKWlt29BLD2z8l8u3JkQ/I8cDQRDAf+FAhwsu4GiBRcoXiJ93AcM
BqZj4IaaQOkkfKpyiNZder0XhTFTi4Emi5lHXheFoeje+sauTD+P4CI9wIoMLeLqCd7nsFo6rPr/
VTy37+W/AF6dusPadJr4LA2gitVSrfywue7zZsGIjyyKIiqHyIOyrMJRZi6dswyQQ+Z1W9p9RFyZ
m7nCqt1B/myvLoFb1J143ClYGUZBd9vg2lxAvNP46pjzkHlDwKFZ7tcmNVwy+6CjfDXE4wMls/B1
wthEPHpleB83mLzkmpIz0d9VxNBvW6nv9a1LkijiTPKVvzfyixhM3XuHeGniUpy+5cxTFQQVOUof
UO1fPC7Vr+kV75MIh6UfUg/GpSdYQHEXkm/0V2Kj5OpqxuSEUzMia0YlW6/I6ZQqBZM1TFKzybXh
pqQUlllfNJH1tRJyq6796vubAQsqQpqI/33eUpDk6xdP9rnmCN1pMKkqhheD7RAu54n/mplesk2S
rAJDUbyoGvpNg7i+huLW0BDW3GXEziV5Cgxg4gxYg2bmy2Nirz8b7gLvH2zcmOz8nBoo47SMjFtC
XUbgim6cV6rjcuaFUZK0eWhZXBWJtG3I6p9uCxRGouxVSNXTa69mxtLGF+nD0cCgzFCuvnsP0Hth
ZuS4izxll99YDC4Lf3Dtt4c/ZvslUvK65CevV0DYXMEGjzzRTLhQSoJpg1PbsnlXV42pu0ABeCHL
KIwv5MU3ZDJW3QSr3Zmi4Wq3wQN4jWimpnNKf0VgN1exkYJhhPIGGsQ5zK4lbcBQ4BDVrL5UEvbz
EyMks1kv/9cD1f3JV9OipvCxRA/0PyFcOosUb/ekoDLXiWBkZ8Zp/U0TFH2GNNbCncA6EWVtzwYL
ouqGPiWpkFdYu9OBziiSyVXPrMxrSvg0vmdFs2/cUgkrSgfT0W4zVGMP0jXNuhaZsjTsQuVB2jYA
Dojf4bwroLIjl8gA0171aKdptzGYcTT9/oUVpMuZxD6Y/itNsEYWz+Enq+m52GClQt/Qz7dmO89a
xxiB3jVUdOtawCHhcrEU1KSsozJY6iOswAY6ktBqCEN8wuTTQEj14SKTRQk4KUMp17kQJJEjphQN
APOZIEyhEXcnzMXFVKHRcNL+wERAZvnE6idq9XX5IcnbaKk9Ho3Li74TbKPRMfn55XxomBFaFDsY
+RfhNjhZkoZjIbIO34fdiFb5PNoZY0Hl5t4mQrDiCbuhRPQ2fW3pjpgtHCgJtjb51J5Bi21Dytrv
sr7NsLIQhKWbspv8wOstX5/1HlGjoB/cG78F9ptD703AqROlL59gW4TtFq92QQFfiU2rcrwoL1IA
rvya7Q70rEOVNsEJuSH+yGULuIaLa3vcAYSIrJONBTw1zwzvWwhZNl3pam16LM6u/4nhJ+0APRIn
XoB3F4n3HuRzeecuiPIZJbozrXXUiza5SI4IPbyMV0FtEYYIn3K46WjcTITEywuQKQfbDLb/vhcm
Lcv4CCr57pDolEojWlSYaQEKr12pJs9cpQKrV6bp7mS+L0zikvTHkTL+0FfS8eaePJoMTDZI6UW7
CJ835kNDs88eZKn3heENyK4AKdAENWI96pZAq86QDi2L4Nl1fC7WuDrwWrkVpvUXh4NTRo/zzhmR
ElOFBd4gOMnMfYd3xh43u85Phppnm6lo46db3iCt9XlAjfYlWEz3cgsJ68/XHuih129hA6duhxhH
et4MluzYqxI/XOhA3TtoeIUGG7sW6OlWmZ4gTganRgFqfMkmEcqfdjwjoNY2orBxVBVvdF24hOeY
W/3Kw7xyetq7Q87v4BQVWyJYq+P05dZTAo+WkLQIrSi/TaHcIqQasWAF/OI3cS/Hj72NiXN/ofpK
0OiNpOfiBDam5jBUxAOTuLoPPHnTZ8ZBfNg37gsFmrEPuMiC49QsFz0F/lmhvIrVNo9aTVTDNW3m
zwm6WY7tRcNBPJ7yZQQKb214aGJMFGnRahkqli3tPQ6UinFIHPO4HTCFL5pSEH1VoZ/qghLhlieu
tRdhWFLZxd8BhqiDTq5DXmwVkSq2uwKi9ykirF5CdRn2iQIfNjuhL+8OzUw7aXKNjka1DRDSJKcc
XD6xHHq5Nz+nYg1w2XvAdGB4n9NX6J+bM8mh7Bqvo1iozeNElO86FZJq2XYMoiSWFog1SmVdaY4H
3jH1goXkgwxlvBqwOVhBqNI4BNor3MHUOzaruGqJGJwk/F+tc16WYG93GGXv+6TC90ScaYc7liNu
i9Dw9A5EjqbEVw0zKxhDNN3moyAP1kxUaW3oE6c4vO4FNOEOW/7QG18WLyeLlRpKNm8CaOXchUF6
xQ+4CZ6WytJ+v8Zccr5LJdWfxzfF3g/kR6WzF5YaRC6O0Vbmrfv9LnT5O0jbC5qy4NXrP0MFIL6T
ERubUy95k0Cd+R5HYVuFPvrBp5QeJZXY4+vdu99CM1EcGewUGxvrvzIf/NJSOfEgsxRfq7kKJNFn
qDpxSvl2Pp+s5c+gsrxv2h0Gr1rtD+Ght9vSu9/b/xMmkvV5HT0yuASLh+mf6ID2f+0vyQLXw9Yi
nG0E9F9vdSyZzElpegcu82vjWzPno9G7BJS8PIONPMWF4lnxncc5Nctt9Er5Twk+v9mKblqcoEUd
B5E+Z/X9kI8XJ1ip7Nv6kY/kMExXSGx1eT3Biz7gwDSc5H3Vd7RHsHCQnUqf49jZzcNO3Sg7gV4k
1qsXOKnaOGlfOMQOMIkLF9VZZ1uJcIiZv/MHrVpdXO6aev3J54nubR0kRdhevgJD3xZivh+Lpf+/
ozPkfVWvdstyld9IPVmaAA+NObFXJ2w65FqCAVFEUe4f47VGeShzCaF3uOaUbmHkR1R5KP9y3nBk
b3C0meHWEz2gDKG8eslXGi99sa08rSp4LK0MjFl9h2u6T2n1awNkzPY/hvLSFJ1mwoSbVPN+gDWe
LUSkGslemChLkp/gkSQCkzlqrAbkGhnAyrQJrzTs9nX0qdA/UVVxAfnBCorEqzcP1JVv4kbtA4iN
sPnKGMR5yor9ZERviZeLcjHQ75XvqpfK87tV2MKiuBrMTDiha8egsWIua3eIWa/zGxallK7hvk8q
NDKApSZF053Cj9Gu+aTdUhDg+qwBduH1AM69mLOEyLEIIO5rIuLQh6O8TMrPHw6XP9+jTaXl6Yy6
ut+gVErs8wfU0WKSR+WOd78n5TRenSTJO6je6ckuccZi32LJpcqd08MSZB2xmm3R+5FoKDnRfmCM
bmdI2rfJ1Y66UXrw02Sbeb9Pj8vaEaiZ5kjFFWaQBcsHdA8BD0TgTwzCs16MFZgNy9zUy/qhZuJJ
tKXIUd6fHwecAcuN0LSN0tTNHD/Nx4DYymCCpPRDQZem4wgY9ewI6a+hdMRCYCgYFxeU1AplZTpP
jrcyvppfO2m71JafgOg8PFS7qBA3KUmwMXs2SUyyQgWCant7s9+Sy8FcyoZ63CDzCez87ajqtdb+
7uxkIxya4EAHDMxyt9LrpCdGbcmg45UHRF/ErRLK3t72Uqbgj8UCYvvCfnAL07Jd0o1mLkW8XmGo
1L0oS/L7qdvHYp7sRGstSGRt+Xwre9iALFzfZo7YOwi2M2auc8bHs+OJK7nXrFsEGYUYv48zShbD
4fbM26r8B84ij5PzAxfknpYrUsrBlOaIP3uCzPkFQBU56cF0N3cE+MBUGYiAWc/AXaRb/mVpfyVZ
WixI2qNttEOmZtM9RaPVa9JbGvCC5TbI9A9vDiUktGY05c9YJOhp8l1KJr0oK2I2S6FkOkU3RFIn
Nyu5QK5g8qvkBoFK84Ffn+qIxzrfcNSfZVLAglyhl6XVyO/74ILgRnmDUe+6fsabgiv6YSvwPadi
Zebmhvau48l1OAVn0NSf86ua4fRSB4X9r+/dgS2ldKjmkMWwJx0Yg5NjIe5yWF+5kToIvmh7gSMO
DGgGIuUsWxyNMzA5fuI/MsTJi72dZZ4Ht3iz3x16EjtDPC5bTpaMoR9rkeDjDnkVgHXKqDcSAvqb
cZjevNd8b7N61KwesRzQq9a414kgrHr6OxY7ECkc3PrAK3bvbsd1uwCMOOZqmGSJ3e9GfZsUii+m
1SD9i/ICk85V5tQPiTiEwDhdV2AeYsCWxWDAa4JAUPq1J5tpfJb5fMs/EfhK8gDx/yEdOAC6pByN
1PM9/SvA8TVTtzn6Yu8Gj3j2l/MLqAf1AY/QX/QlMuXHmJwYq4wcV3sL1hErtFmadd9O4kj6nDEV
ZFevWMOIa9vFMq0BFRFUzQvYX9Uv489/GLS5QVevBrxLCuq1V7sPUPDRF5BuGsmrF0EDZ4GG15JJ
2/PoJgibFmHL29nbC6XEYSmAqksrlDP0qvQHeA4/7prNL8cfhMVrT9Hl6JHAncSOtwknrQTvBz9a
PuD41EAIsXXM5LTmjZYQHC69DfWfrNWu2WxWwkhrA+2W+4TTj7jA1CiDE1Buh8qSPoYOS53+eTEb
Ahgkmr6UzWwtE5u72+oK8T58ef0y39+vcVp30pyOC+6gsOIdSr0th4f/Tqv3jrODtgKbAK70g6zs
2lzao/tsaQqvPHVhjVYUzrhRaCPR76j0l+SSBa/YE7c3psHLFQ9SBWPtUVruc1dbQcrUo3fKTQiZ
wFQeyspDU+N1lJIcQkaYAqPYtrNzEWJ8MEXjwuSpEy9L++yTP6gSIdWNbH4kK+DsdtzHDfRISPRu
3UHtn5UnoM0C+8F3s7sD5V1rjWDiEGbYgug26xQQ43tUwsSMBQataUoJDXPIJz0KCwo0PFA5aXy+
Iydyv5zxYZc/w8MahbtgDSiT6yUpM5m2EEyaqQeTXY4cei0j58CCyD+es0no/OOuGb2/fPpgWYlP
t37QITRnT4neb9hCYWbYuLlf+Wn3SM5SDDHpnM0+VlOZpanW7vgOTrmyVc2aRyoPd0TdKiMYx7RI
Gu7+pTLbPnVGTqO7u8p2UMwfMbDo2NFInf16c0XABJFEZT6VELwdKDYAUrMjfc9B4yQXpZ4oqsn4
dOywMm+mHQElg4mM30giBg8d+sk0v2P2nIKdQj1bW7uhhjc2pws2++jsMz4QmueKlpz6W3vSK9zf
JgJuC0I841t1EzwT7SNha9uO26TLHHKBf6tRzy2rvMkOudv2GP4oLur8ns369WtG4/i2nuXkU3hH
e8l/CcMGIRLKZc1lueV9vkQrTr6Vu9AcNyvutVWY2QXhXwMkxkVnLor9YYf6BqsHQN2fpMDRHLqx
wxJxBlbKhmgrSvmi7hm+5KDHYSMmuR7YhS67nUSJ7A+BVADstUksUOwvtlDOtUKeAWGOs6jQRmeE
XqcOv4PubsbaZ/dHEzRxracVfVz+vl69GQcVyOvQIBNanL5raBLomhR4psbnPyTFh+eMay69P/0W
KiUpbGsG4Ga+zWo24ynkAPJ2QllpTUdHEdbLOsgJZlRDlPxgWi6NzNXW0QMkhQ3z+/sDatPGe32h
WeNLUQlYdkYA8KwyojS2OElGTZTuYx0U79jiTUC/LgP4eJyv+wWqj5bzzuudTrqpuRjdJNPGigQJ
pVpinczhOOS6ELJuYrT5E4Bi2I5LigxnZmi0ZP671jiTTXseLgG4f55Pyuf6hj0Qx0qWODEQkJxB
PNNl3OPCWZc02BQAk/mepY8i73FVh3pjGWByawozZb1jk0MMl6e+bUyB8+DpUB7ZJblzIN6bMXvZ
Xlvgtq7jtrxDowWfzeD42Alu4HibxuG7ja1sZofxqTzv9C3ZKhbZZ3qY2LkNkG5Rl+jhoPfUpV8D
Ple1twJEBBMiNRrar32pf6L1ScFSqKC5aSEp5ebUf3l51jxa302MAmLzMVCOMGaLAc9BUZeKtr8M
pzokMR9419H7AbpSM7UmjyxNunHA1WD3yrSVf/chcazkcEWWYPKJzgUGczJJcL+IrKB9ueAInAfS
6/6nM5HXgUZAYjmODaHcq5eoeDoAhW/11dqRO0OiPm27gp+Kq3dceIvxHppi4CSoUR+zWn7ipcrQ
IPh/HAqYdEVhHwvkWzRWhcjq1D8D6hZtHpc6BBRh9GVX3Hib0GlIAHWCC1BkcAUpVi5OX+Ji2/p7
OP9LZm5J0HNUESVYYoIhYxgXjnJUJN5Ibn0xNOKpPCF2btDvkzMzYOYmPQzlRa+ZI/vTtc9CCuQK
NIwuHtBQa5rbZcM7IF91k+e0EqjoiFxAC2hDwbHKyzqAkdlOI5TfqBy0VatFGo4HeyyIJ8DOXDlY
gROKxpOt2EOlreIelBwJPy9qYRWcNjuxc2YClgtjG6qp8dZDcdqk6iNaJqyFBekHmeHGlsh6nMI9
qvMz5qiImiPEHYCbZCL7IaChldakJgRlzT+PxutKdHLE62fHWW8iZ0LPqL9QrjueCnsTw4qKGahL
wS9sMaQk65/165GBK0vNhNxkzJCj8dFRozzPeuO+pivqbExNhRNP2Fw2GCyP2zIyWa/QmhUdEolm
VCZWkhTWFR9C+X315u/tP+NhY6KSOb/noT8AfJREVI/dwMKXNv4fwZrawIXjWI50of36O5WyRNql
sYvxzOas+AH5mTqDHEM1pwnYTwA8ejTUOuX7dH95rZTFC9iD9QrKCHoEd8Bc2J3NHGJUWLk0kKZm
BfDeyvS4UWb9jtLcOB8ZyIFgwJz2LlTsQFYVoM2mZ+vYsEGe7wS+jTAUDWAnst0ah4bxzie/hW4i
q4hVcTSe3ieHSsHl9M94JtihI5ta6fzj+m6yi15bbDfmz40wCww4B6jJgtsWuhcvHbdlh6tbxsjt
mxpeFuwze4epNJ1d+2sYPEQjUI+PPDQdy0kL1SzGhuqkmH0TLl9qXApbADDehZawbw6xLw1kbtSf
RazbNjuWdoiXXhWokMVos64ZLl9C+ltEpDV07mEP2jBzJQKSOTzSaV4GDKLLQ5YfZdLPVKGeTjZd
vV8GsYJZ08elQ7RQTyg0Uh7VfeLo7t+YRfV5WfpnHseQEmws5UMp/vXbvYTpG25N9vn5frtgIkBr
qqQr0NKO8Ob4MTD+HLx99j4Vp3vBd8UXDXphgadtHyNYWafN+z8pttU89juIsAQy+SGi+I+vbY3z
EyKb9VKAeNd4vKvn4+1GTkW93dSQx5XGVDN/RNT0BFdFwO9K/CbcFnaSbfl5XuMKAP+efTCa4JWr
Md+NTmCM/bXD1EFHuu3m3g0XDM0+KDLI0BR6oVtNvaQgEOj0ZxTXgDyTGOVZpid6m3+Ix7JJViQ7
A1n9mOSFkquogxjUOpmTcm1W4HOsweUO6PyAKrWA3fRPThNtzbkVyaWgRwqBSjGqqPSm3NMtoNnu
ki+9NpwfNYtdP1J7sbPuJpOwsQPKK67e42j+qdg2NyFeUYXnUSyyon5c1lVUUZLzSQJiJeofQtf1
btGVcUcJimAwrcK7OEIxSwwmcaRwjMQESG5yF4L/EedKIXZl1vVjjWV3abEQM+UObbhcdsnGouJ1
wyj5K6K6gpbr/K2/RNHhQ3Y9mRhSW8ejDCC1lh2g1ZRUB7b7Y9MSDGZmzx1l5RDqH2T9hfbcEK3U
qX3zN5vcClrqlwzhoSgQsa0E30VTlLr/VeLgnqH4VSl+D6+4pYs0KSznhwSFwru704rXMgrrw7G8
DSTP0H5HUzEwEYqOMkzkYiqTbOUeEJLIrobfufydcmhL9K0JgLpP7fuQnhOge5eD/hZxbDOnqcrF
r0FAUtwkSgDjZ66G99Oo3Fytqtzg9UtGg/ds1Xpeiwt6IUZpkwSEVhtjptQKXRzfc516z1EXVP97
0T3ANcZ5JCFNZ5BYBzkplZCgf3cx7Ddp9UnIms1wPP/EKMHNUwD/F3zNy234Jp012+ymurFu5gTl
EAokT8mIVRROx5+RVLw6h6t+TDxA9NoOLf7eguvdqGKueySZPQ7ac9t0yZb2v6TB7v1ymyL90ib0
UhXnNRFzoRct4pytw27Q3pl2JZzn5jCVFcBgiCCVa3CmKz2OINtxDdJYvpDeLvBgD52j+iobwclL
NrC+TBtXSXjEqwy5Ja7sZPsOZoKVp3CTkF2gVsqfXFiOxnAcC/C2aRQfombfjapkR+KS3dOxDcmc
0prk7rIcc01nGR35Lz4rjd9MUCsXqn+f+CTUeVhtcGVfYg8AuRCnNIaFznJFDElfGENPSVPxbvBB
GaQImabWNTYNqsyA7vzMydjar+VLsST6k1DwWyq6LWs+kok+q9zbC0i31VjFeJ67Gv+JO97I9k/Q
M6SSmkIhUN+fxpvbCbwXhQFtBYfmzC74ehULpR2VWjd+5LtNWTOCN/fYuea8sTJN5ClgGRN329t4
Jlic944w+8EZjTw67ldlJFCL/fB++cLsGqt5Kbdsm2Mtfw/x0f8qvZcdesXmD9Nah5sP0Vwf/iZV
NvTN09G4CjvuP4YKo0m/TD3LrM2f9hfXsuHdGIeDh1Tq2KqOPkszoQMiA1dP0k7nbXZOv5Ik/scf
1gVGsS6mS5PuuBneFT4J+fVT0rIBFlHRz7f+U2jHzBW4p6zhcY8gN4L1eBWkmx/dqzfo4oT96Wus
drEK353SnQv6q4mCjUK/sWZgiuF46Ynqo2X7BnqYAtQsp6mmxQ3qIJEX3gpNnBgAAkEJCbK4ooYs
oM/gwKfhbT//BTNHBqiLzmqQG2ylnjA+76hE/UoRKWC8Nh+190txNhnikQaHGog1MDpIkLID+kDf
U+7SDy/ksYWM5P8KKKDenNHmxhq5d7kXX4NH6UnYWVwFtY+MAQUVjD7KIKoFUDNsg6z2+mSPt6L9
bzvddJ4zf7ChmamRoHsTS85Z8IpWO13ygFtu6BRcQob2HAmXmaEUG+vUWuzYv2trxKyf3TJ7zXUo
+WEfwlRhnwyzH4CihkeN3N6AYDCHjh2eiWbP/QL4a9CDdKeBTYPuLzvb9dDeq3WQz8C2RIcbl0CU
nMDdMW1fSwp1HGtZ8wXh6D8iMqLnnJY2Mai1OjJN/yrXb45FSLOmz8eEgjgdcTzHlynMAA3chcTy
GpaaknipOVMbWp9ySFZEjDNHrU7zUYyyUYnq40xk8+sbRximPX/3xagakZGlhpUM00owGJCS6YqO
mIJhqaRUrZyrBJvgbFVEtMUID2kXcXnN007G+Stjk9RrXgdso03zVSrplNCBqDOmtXl+9patBB0x
swvMlY8Pk3wr/+JFKWdOEANYge+SJAGvq0oGox6vYMARr0O/wc3z/kKWtT2KDmaZnsVf7fBEN510
ZCu+a4FvOaBd79YanTDARWrUtFiCQSDaAWX+u2OhKjhQJ0v5VH5Q0Y3mInvtGNKpsb0y5Mmany2W
6SS21E7rD+r9geK7MiebOmhJdR90GRN5d+/ELM/3unytmCuefe6rf+sJMwSmlXU5Tfa9p4G/TIsq
/MHOH3lL46mahSGA67ZmRT7zfoLfsoRKZgi1ivfMck30kMAnMBRMXG8k5urmPX20+ROMqs5gB6M2
eWz4DzrB4T9XudpOfX9whhWtlK+cRzZXXvwmsceLdi5WdOroIcTOwTy+CqSVa6LVlIxQIzXp0BqQ
V5SHJQaConkYTSVDxqGgFdfRqYdXhm5dzUdRAJaFRbq97W4oweh4KE2lLhUFcyTeametMyoF7Opd
PUvvKpmJn/Giq3l07VEUWPgHg1yNZDw718EUlwY3O6v1XfndxVhgOrugxcmWCryCsT4rmQgNxQC/
ZbuopLFB79u2eJu8j8FpEQ6+ohAFc5Gh2mCucs9M5gBzsK6ZNTcT1EXscZt0rlw6IFHH1zU/f7aA
EFcDljj1aha53XcRPJzQkuMJT+KMV1KtORNo55hWo4XLnIEvX3wBkFBVOolUyuVbWZcJfpGgK0oG
bDYAlEZlmpCRlGQqZRdbdeowGUiPLMKJY16quy82OcLUBN3jwAytaaD0JLPKgpIYWqh8m36pWPGV
DDmAEJzgbeJK340OT61DFJNomuBEywRGkUEZdHTKyvnQq6oYcDjkFh8glsWLFsLOVAG7WeT1wV/u
aqbd19WJLOZujxtzYSfheMMeQ/bBMJtFcVKf/N9jG4RvGXz1KQ9wtyu7Ek/SSCsk9KO+bNAgXTj5
31wwu1qD2vOT/xe+HCQJP/ubLigG6YwcRQDqJNDfu4W8tXR+zKtu0zDkyjL8kUvu4b7+SonCwT+s
hzVelotAdlGSmwVuueOb9PxzkzsQF1yzbv022j4qiydufcz6xEiOcQG5pRKVex0WX7ZWP57SCLtT
7hReuHx2Xxlq99ACSNHUbo7yBub10qBznhDfTXeTBC5WAQd6/1dHETS5n6gfPLIUc1vJOLCK2X+t
bw/TZUcUjLNRlSAgI7FynY6BJsx+x33ReOUSFXS20iuikiJXIyQk3oXD5tN1SjetePRFiNUSiOnY
7OHtn9Q55KfKMZGsMq5FN9f8bf7lCzbhDSL4SU6BoPAnjE/GZDEB9w8v3ZOY4ZTKn9QkKafitl+1
goy/AP3uakeUwcvT6AtY6HIAmImdXMO5xf+DXce3N1/nkToIy65frXTIhICdrfvBjewBCSMulYxS
LfXF4Eiqi7zkDIqdAE0OJ/5vOdHvVG+hDuJ8G0Yz6xX1VJ6fJHD9+H74pVahwwcMHMhzNV2uM88o
jnhsdGAbFRkPaSNAswD4EqONo2IcA+YjEBwljJP7GdDe+3o0Cy/tBe94ViDBkaLG9zqbumG51TkR
0qY5p8VTnOjeHidaH0ofQdK0W0sIGStDrH6gXlkJVt0omXRGSeKIXolGCTxBuJlqj7oOk5VRLMSA
GrnDGGRXNvPmgemp7FnvUsQlmRenSxjRcrR6+b42aHFyxYH8IzyYlVoGufbnaFaygk0bkP3ZTRUo
FIxKc+NxQIqfSoNr9Asr87tuV5m972f9wrCwOeESEIcbDAe2eEDCUSHJHC8xubdJXdr4TXx0EjBl
C1l5REWv9Txn07FhmC1r2VvV7HaWDrR6clAa3kVGH832gPe70kBsD6djpyaBUy9TSsAr5xHLhc2y
dknrpgwkDMEFNGKTHpdAzF5z/iVFSLRvs5B/+d5/2XqfQG4QcaDbhK/CWBbqJrYkg/U4TH+1P5Jg
gsCt4UvRhAUWnUJ2PUK8/VBmBFcG86tRgLmu1sh8L0wFQFAubR25Zz6etsfwX3o1P7xyu+925oXr
etgtlXlBiCkhKaoIAGrnf9dqIAQDpaRR2SndjxXRmVesE+DAU3xNQcEUPm3oK7g3rJiT9fHf4Ym1
fXf7Sm2/Mb4Z4m+wz1UUX6OlNxamZAmpHwkPjpDFbDOg7fkSZ8qxRbbUjQKenPAkEfmcnlRvagIN
n3oGGKwVGvlyKAIe2xu9KlX5DXHUx5Pre5xSAJvuHd+y6ya2LHitnoWebNAYbdSTHEGiMyYngBzd
kOP12fXnav1szkXTyLhw7WOljwgTIyi+EPHEyKLkN9feMr0HFIaSE+f8xsYeZgfQ8zUSQx6VMzD9
tt1il8a4tEX8ifSKeUwg3v18081nkjHWwpgU8shpNKtjJUwAG5QE7JbWS+mH72CuDCAX+TPaYUt6
vQfHNFggLBOc6FPzEA+xqqyDhsstYCzUVjmZvz4hCp1ej0dvrBBQF3BEV9Mo3lBmpC1ztt5mQkx5
6UQ6FnAnDwFnVrWsgJ7A+gp+3MCml31dJc2n0jGunppXHf4Xqsss8gwjUYysijTXIj+syIQ0axd+
t/mk/8vPXO8x0MA7z6rn4oDMem68TLKIFxFcKN1odwKeXisF7d91P54aBaKOjVt+0eLsx1M/xfOn
Mn7F9zvXbtVAxVpsEek+7Vlipw9b+1vLY+4nMNSUB98rRrcNBcLlXFPQJU23N0xS8opZhtHb1bVS
owtscOklQevK82pbBJu9h005DJbM9TYve4SYygUSP27QuHCNLA0GA01Ijh5FIBWt+2yUlGl//dVx
wb9kVynOB0OPcocgF2wMu+t4qBplVRNei8wRi2RLX0DONlBKkSyYOw7B9D+GYn8GKrkyvVfISun5
+EPmJhY8jtatNQYMpkF3eUd+k+TiRTyAzpyHr2Z7Vsqp6Yc14XXwgKN+RPPaPtikAeZJ1hI9HB6i
Ewr4WEKhtAfjoAJXQzniyl+KkeTMSjoZdanhNPxBAvbqtJgibLQn67JkkUC+POPxwuLLNuWI4PpP
EYm0koe2D9kPltB7g06BJ2CVh5OuUasFiLD0uH3iqqApJWM+ciIfnjwICp5QAx5tnsaKL84fgzDp
jC7pbFS5/t4ziSjxdtGneXLc0eIjNKU9jBbil/xmQ2DmKkTvmRiMw3FwRm+RSQawYu9ZFBJe5xfE
J9kwOHLSlmabViyKtxRFWqA6ovukB5uQSMf5LzH0/ZnkAzfJ38G+rjijDvG7VqnO1TTSIWkE1oOM
JG9vy9bvm5oT/9F823jGv0xTd/Axrwpl5ZmOJEC1TTaind9p8X/+pttqIR4e26lZiKOBH7vwSqdY
eQHo+Sj+8Z0OZKpiltPN6poysgEEzmaRiYVuOW6oxf9uOGoGFmAIZ+ire/SyzPkOBohIYxjEfdKt
u2EQVjzknE/ue+EqcPPPl5U2Bvpu77grboWugrsBFqL2ctdFFAN8f2/EuMYddpkVy2WoGf3lSzLd
XDu3fo81IkgoEDu7DLEFF0rcBd2FSI6SZVeXG5cuki0Lpkt2/uZ9IIbGSeQ1Plqqe40wgYLPlkVx
cUVhAuwjZa4rI5aSOS+erVo9fH2T0wNvSeUe8Gf4qYKwizMSiyxa5qBPcn/CMHBKsGocB3MiDoA5
A5W4nnu+/phYVsSEdo2D9f433qXVKith/RSnPf9mke1CCdimIGeT+DPdBND3jwhVav+jh1qkCLnd
yxSLHAgWTvBJKQj5nFvXr9+OhY63c98p78Z9QnyJESh2HMvkQWFgWLKaFJoj2FJiRnYpPP70pDSt
2j8jtshV0TUSDjDWcg2Ep7b09K5P42iW5PIxy9INKwlxuWY8Ojvsd7GDkf/uCuKk2CFRLm4U20QZ
urk55DKoApp0PfvkTLWK7OYJdOOFK8kVpBzF3k+WDPq7o56ft8X5umH7/CDhYiFF8BtOQYjJdyse
w5MjCq7CdcgmzM2Duxicq1QJzsk0gil/fGQ0+AChQt3BcV5LPnnOhvy2KGMCfBzUmTPSjN5+Ih17
G14xXwMXdaeYqZgRnOzWSAaKc8cp3rgn8u/rOUVSStOua4bhMpIWXzGwMxQXxv9fZHJbPqnTNoCS
CQTZsN4pWRruYyXaSE5R5Dg0e9BFud7s2xqO4jDDbCkX+PrQFLxZ8euAntoxxHrnzzhs2/0DFgbs
RlDOO4zSc8HBJbRkely84sRP8D/Z2971VJbo8lttVdr+S6m6QQSFGteQbwuYDPD6hEcM3Oc7hMGt
LlniIN6XO6m0pia1YTvLBFNUDxABC04xkpquCdcjlXDuafxYL/SHHTSZNAYCJoEb6B/mLJseUKKE
N1Ilsb+du7ZMmP2MjzeqHKDOK9Wv9BWJfgmkatkcK1U7a9/RV3evL+ZHZXEe64QoRbONY0nX0Lg1
ZBarNAVqUXJZr+4jXc5giswcxUE1l6XApwhpiAV3tDaPYQuXrVonpIm0eeZugSDAtthk9KEo4XZe
T6bV+pnRcaKMxsQxxDS62HDxroKDeSd45glS/MwxVAwdyA1Fx70c/DVp1LLTGcECQ5IV0+F+YIc1
+v+uMASaAy8PyyotcOzB0CoKUReIQ/PNfbGRB2cJC6nxxD9Guw2Uzqzy4zKd0BHruyGWpMVJCP6W
rkLBDe3Apz1jX/e0FK89KnMjYPalFPizcXlQO8bgbLXKm8ejRnPSV0xmIvXaIVjeU6bLdZ4j8Alu
Go58tfQmTKFJyUNQuUy872xLMGtB4GulHGurAe99RO2XQBQk2UvTnHYf9M2+/bqCEvbE9I/Krm5D
N6be/xMZREBHnT6e6NOrnJrbylnzqXG1+0BRTVILXXQqLxQmrB6cjGWAHEL93hP2AxXoQljPcXX2
h2gq0+5v12o40avgOgTM6G61cgtsPdU2/zBsBwSv4mbyJgspu/WMdqTijTv11Tcrz7Yp8LCdFHjT
J3qlsTuvJos5VyvDPcYvtDnkqUbKlfRWXNhQoC0RzGUPZlujkpfKi83QkDop8ZkK78DS9O9kKUnE
9NC2VZT4LmS8FcO+ASjX3C9Yla9oLM6pZz1UrlYAMD3/G2MCxUOBq/vsyDUotdTJBvKO58xEGIdg
aE36jd8TWK7przS5AMB9rbDzN9Wkea221f7LnYE+mnuwO4Yjse2fQeF4Q7em8cDnPfj4iIrP53BZ
HuQEKqAYLq722tg6Eq+NiipJyif/E69reRUwsiACYd5VjnQ1smEHpfOyuosd+KqZqqEoq/vleCKb
9mTuu4FrB/o/NhTEJtLfnkTrthwA3w10Cd9UAkXLsYOFnx+fWBTbG5+ipxFggAwONrugAnVncpvR
MnqjS7lZx2YS9LDIf7EKrkXIvlxnHQ3byvR+f5Ac5lneAtCDr7Ksl2R66NjCR+pBkelCjekEnw+t
U8CrS+gGXd2y6bYUWRGM3OS8+Zj1tRuGVbRS2+K855eICmQa7UcknK6RUohjtXPNAY3WCCq1uu9q
xJfh1fcqyFx7xa450EQCq4s24Tyh2ui5aSR5zBRU0Euvs3Y/YrLxnAKRC6VHsi2d3rP7kxmPtN/l
Jmf6DrM21LOgqbz65bQb7chCAHuiO1RuuFWoo1/w9Y7ZK/S3Zv8Fug9maqtIQCRMbTDoIvcPVkZR
KzeVDgPC8USHNjkhNoHPaCrauzT89hr0ogk43wjwPYEcxOCFewJSuYhSMQH158IhEc6+6wyWhzuK
I7XX+QnTn8dWdMkgBaPjSgi6gsTib/6z9VOeFJJF92HyrA4Xc1Bo8zBdiaxlnV0ffDciEoPBhdwM
IRAG3YzRqr0Qbvp76e5TAQQ+kJi06CpDXq+HkyWMRs5avv35zlhYNMU71FZY1G2p4yh5G+nh7rJS
9z3I0vt3N/in0K+eANdw8bA2sRg0SyPuUrCIhhv6Ql2qSg804Pdyh6H6nk5ou2v5ijfzGpdEdwTs
8Xou+pcqOMZgEw/ZqJ8Y094YpqIBSRfC/RR4waNbMp6X33WI47hUZUd6hyzEcPnHULoHUQdmZJEz
m+UKGk6tRkRzs0hw7fk6SM1TqIfY3b5oHikJi25PbeaOb3gCtM0o1y9Jn34NVoR9lwIXtZ6kue3C
GEw19RdiBoVMmB9vl25Yy6yRYlNJA/+WlYNbJBCfjiK1H3tEwXGOZjcGL7KtEOE3fcUZGfiKQQwl
r2jtL/okhtpIMFS8jyQbzhTJgH4rt3+r2iLs/SjA7LnfyWx51V1+nNC8dc3mxRsKcwzSi5Bw1Z3B
mdKlNIuNQIupByWlIwn9x/N6M+AAwpdsJRXOMxWxXb1t5G6TBswutg+737OWG4HF6pIdE6zSVb05
/R0c9f4+kd8yY4JWzYtJt7GzUfB9Sk5x7y1SB4XST9mqOZgNjs4qrymfPRDtxb0mmtvZyL9zxFCy
VdtYzO1ERVSeGky3dytFhB/BVBpcJOyLgVPor2v6mOjjCYMVETYOnOV0QoKvjQWAGV3U4a1VIDTl
OYG/9tLLfPnXwISuBdd9epOp0Z3HB+Bkw9jVkutvMIjh4mFVqcNyDXDZHBNgTGznCWc/oad3vWfp
xE9sWWGuC9FZQH6ffy0SVrG8LwUK1MM6Ezyh9o2152DYtC80CAJs13z3tVauCKOfnCpPlM1xzklA
+MFpEvjVvBXCo2N1jywojHDDsBc7lOfae0Ld7wBAv+l6q9xrLLpTB6jqAqboXV4EKsx8Zqc64oMx
9Ibzi5VQcEsmSTMrVeqlPSJwo4Fz4OS8HrnDacsYvvQKTbmiQWsM3tdlREpP3Hbs1tsyX+9VEty4
5Y+JBf7ru263A7vfGrbZZydroLO1TOo7nyZF8GUgjDtbmMJlWDkEcGZPbtyKC3xWxBycZpKMRRmU
p1gd9+Zfi0gzlkYu0Ylyq1pNz2Pf3sR6/oFzLPumLpGZMQMFYN8lP3O7i+ESD2dPfI/riav93iP9
Gl5O5yJ4ONXWg1tFpPW8urQeXUJrBSSAdVxlj7WSIX9C/zg24K2YWKy3Y30+/ZiT+Zp4GaA5FUZh
8znAVUqzVgOy3IUXc0DX45e4Uju06bRPkuR79Rw3DMEzCmQH5lC0G8bpOzlyN3yhNy9M05T+lwT1
SSdNoOtiJmUq6H5oS2y6v7tnNH7g9Nih/e6HKTJuoKI7W2MWaB/o4UoOVc1MbGCJlNe9dZdPL2Wn
36Gl4shM7lnxjRmNZeqzHvlbavbJG/BcwWHA3JMr4wlPFqsloqleRFPq12Hfsutm5OTvVIawN4/M
vUTClpveeaW5zCRZfE3J2XVX9v/ybx08y3/GrDcaZwyOwpJysTEeEehYNsp9EtbYREiBivnGfI+C
i+wN/3v0SodgZcrUU1p/AkZHDQ2Uxaztj/SjtosSLcuivRyFpf09IvUDmY3u5ONGdb/v/MumOd4D
adWOLMs5vOo1ToLQvguLGH4pKgXRfrm+uWmauVq3fIX4Oj2fkm9Ut+Asho0jIjUDEDmx+y8CQ5au
pi7IRRr62m9eMf9Tuj4Go0xDS0zXNziZVqSHMk0qHAn66B08VHsGr94yt0MmQK3L+YTRMunzZvux
D2a0dtJIijgqwUdodBh+oVFdov++pkU5mMQioIPrWJy0QqzkNfhYgwuNTjVLh8Bynxghmfktjzxh
fmGNJ6aXh/HvHymf29EAtKGMpL7db8+bxVbKKeNNVmpTA1hR+IuY1qFUdjY4T8cl6Isas+FhRqvI
AAF+fTjmEXTjt5j2smodvvjsVNPEmcwSDz0/TNqbmwXKo678ZtsfNEaUvnDY0MihJ6Kx4eNe9brF
DdkkEPPWOE5OSiZYNUOo7KDxDJxEhNTMnGWAl+7eD6Eq41OejWYZIdoyw05eEuQBMQt/Bf6Vkjwl
DNlxvws5V4kwaPumoAC4uENVnjWXumGVMewNPUXuPXAiDs1zHBoCVM2Sar2Je49PQAiBCdXzZQg7
73bu0qK+zVYPDIX6fGrAVsFyCwCzSR7dtsLwT30aKqxzmnC7sX385TslapSkQK003uumURTouNvO
egsa4KFnvOX99hNwIJJ6NQE0Q6Tf+YX1Tm7X3dnQS1XSlxTRw08MYVk4KhOA58Ixxe7yJpCR/U5c
GMmFFFxPop0Vea6pkHM4RgEAXfzYr4rx0MoLUsKERiNimoTORsjShzPUUtd73V0GZ/lE11vr2WPn
S18YqIO49xsSpC9/Vgg8LMgKJoh1SCZE7uzOWwROX55GFc8cf/P2KW/jB6N4BYRxQsVs8Vr1HhvX
83kuhHzC63+2zN/c670mJWXyvHXajb/usNlRNZyGRYPCy49m0iCJKW02Xo1c39TNWVZkiOs/EVnG
BAJDTZ/G4NzsCQukakbt7072JPxWbPKly7YP0A9mcMfjWJkyK6t2C3JPPnldarj+9+qd7Y5vVcVZ
X57Hc2xRiUujIthJtWEfAP3xzFAzFqPzV6JMCByhs7bb1TscyVd7AaBWBJF9AZNA4RlCwN4vbo1S
9LHZdaaIXPrj0V2z+x/GUcDUGrKfzUFe11a+vipr4Rvy0RhGPO8XQVRsPuXuMH5iS2q/7c/LAfmT
AOSEehKU1hwUdAY/Z132dpXqE+nH7kmonif8afwdHKqrSofIksyGHHI0O7rPqsqtDo9VJRhBf4gB
kyVpDg7PuwOH5GuU9iJFudiya0SmBKYEuD0NWXi6jlilwCRiLnEV/8zBOmFDlKXorgUIXg3cI1up
rMswOE42WAjTW5d97vsD2omwSYrspsCYYeHnXPQWzj0oPE/AQPgUk/suF6zhm2utTW4xSOZRc2ZW
t7WVHZP26XMG0cnp0wKW67EvQlGxUR9t73wMW3G55UMsqMnyTY8oXGKerI4tQlLAzHxZXGmX6cE+
SqnTuRmBEfHRV0bZJY6geAW6GVneSYT6Ie6gvDV0iZslXVHguCJlvAWVcHlYLLVmK51NOlfSLtGz
G07mHO93PpDdBAB7b2vKAXYt3Rna6hawQ9N5MlQeS90JicxH2dwtD4jIrcD3SrSG0aOlxYNWpsLO
/L9rjQwRh8jcsXbOT/NBWAD4Z0wSlrTph/tbnt/X4zugxBmkEfv8h8cyR7IIgU5jHrjtNTbwyD/j
xn/7AY2cabj4nL695UR4hE2YPQApoaVxpv/5Pahpx4h/MaghHkQlCtVEF7PmmFsRnBvOU6be1uM1
0CMSjwZ7OiWyBvSRoDYPwofoM7FZ9mCqSk73+NP4h4/I69kzEaZSRJWSWk8tCFFhW7dmuwiKrP5n
6FEcQ71LfnRDmRYttGeuVb37VxqE9ehOr9vG7ynAo28GqUiXkMG9ynVr+bs/oX8vLNdyXEN7zGu4
e5jlz2IRNcs+n/MOYFymNFADgtRfQ3XJMSEnEdq/uCMTV48pbfgSrMeZ1E43Bowok4uhq0xaTyIe
YeD4QFohnuoflE3CbyCPvzvh7lbhkD3YVXCyuy5VzMnmywJrybhEP0kMfSFo5JmfvKvYluaz1huC
Oga4GavxKoT9ayhd1WKGPCSd56u5Y9jLvDKHlcCA95969xH/PM02ZzO/YfTPRNgBhNh7moCce2yK
cLzHcNMZshes0KqEnWPc/5LDqpKw6hHiggc8mY9OmlNCv2zqlsF8+KiM1//SrO39OUTsSO4oxPvN
5bpUb7NsnEYuP9R5MUhFl13GpKn9e9O69kCeFocKKq5/S1HltPAbd3R16uKcurEjIucmeJyAh6p+
eYrlMN/7Nw6i7JShHVr4UMN7ZBuIfYkbn5QqVLjkw3UYs95a3ITGQGwXZo9pN2dEh270CzmfgYF6
he+zNtSoyxPanwLBwv+WwSpS74JhYxTP1doRp5ZIcaqVoyM/C3zodijonkhLec4DtoDMpAJlYOq6
pfDK9Ka58Zr2Lcq2LYa2/T7hVgjgRHwe7n3L8q73hB27FP5CGcwt/hwlbi2mRBLR9MWrJLWJC5c/
wLg3kJSrvS/pQSow9qEizwF4kHlxgutILJQFgfLElvK/5mHbHnUjegJMCqSldM1onnIhBzeuYgnZ
o3VnxGSORHJcInzeMdm55sTMuVtl9R6Bek8/5KX4Ju1N/g3Y3gVbAOXDv0uef4bKSJQq+YGYH8ol
4anQtkRDiY4KmCyN91f0KjZNznZ771KjuRpZJVn2HfOswxjnN5BDxLDbcePd+4Kh0T50JB9yupw2
Acy32VbVVUFVS7Dx5Ekzdy8k7REDx6OG2iasv4eZbNj/9sa9hiLNFJbZjou866D8/zn58gd0JPpW
Ujajq5j9xAjF2ZbUeGjdfMc0GyDaDAEocz+2ZOP8kN2bRHiFx4ABf4jPB45v0bU0v8/vqvA9//0N
UnfvHsBiSNAZ7t28yvFNjNMdhROKHM3xGedlWhTwSX+y4dVEPDDybzXIeMOJJ5SwtV845QytDJJe
II5scd9NrnzIuR++BhqPpUbTPFK02jwgDp6RIN1Nl04wbLDMjW8wdMSvU4vivIGrif9Ivmjl/dIQ
f3t3RvN2p9m5AKr9OBbRApNGgZm4n9mKaE6iQ1YZPGmKSCjPBGOzGPFuh/qiLhjEOmo6tGi3Z56O
Perjt8D5pmsp6fuLXSwllsy4m0aU91p3IuO2lPZx+5OOn/abHR6Z6aO996W288B2Fl5chiSiQNB6
ookD10YfxnLrt40AjV460hn5ieyV4CcovoRHQtM1+8mrfADry/QWPIBUgLqAT9siF6pivIUrUgpg
70XGegIPKUAbrl5H3d6zY0Tw55xB2or8mXO8GqLDTuYWTzL24s3Tcpt0gp2XgASDFaDwp1nSfIc5
sCADRk3+uVRs9HZkf2Ybik9aaBe1QirNJnKHslKOGNyFPEqMKhonLws1BSeV0OeV8g/Bq9PcsEAO
rtvPXlFxSORw28vkCjtzATurW2kMTjlzDlowea1uuQ57p/Jl/ZVIX7rQ/wihjO5/GIXeWF7JwYI0
IiTTHKGeuLnsgty3FCRi6iWMXhM3lFa4kTEQtchZLVeOAE+xwyGU0Fejy8gIK+mmKp7EVO4+V3gj
IO2MPzgpLrCqNayAbku8wYE1xCKG+iRpGGVLo8MvBVcAu02sICesqZ81fJSXMxZNW+qoGO2Qwgob
nxaYGZkXl/avC5TVSPJ0My77YV/OGi3ODIjHyj5DLnlVEChqfyDPwNG4X3LKVgcuOoXrIrjRu2no
sXzfSl1ha6PkW4gEYghLXXgrjngWeBphESBnR/6K1AQx2qsEU9wCR1+Q7sKi+tChCSA5boviVWlG
sEZIR47p3hoOhGAwoIPc0HmZZ1+c7XZuUv7aHwbBkeilKRnTiEkWL2jFX6DtYLI5PAwOFNgHibi2
HcpDceEPD0kZpUnGuqmJc5wDoDj0tzS9iu4Lqazu8Y8ShF/U5eTSus/6KPQDoehbbr0DP3gSykxO
q1UCf0RVu8g6WkzXISDFmPzU3GlGk12SmmbOdrSYosNGLCL0fI2rM8oTUaMziM/0r9DzhUgni93c
WjpWbHlLFmkLL1SE60cavbNGnPMX17WRLzY3/ovS4NzvKiqJIOEUI3H5MqhAsAgQ+Yc3qEWdrgd6
jJ8AJM6v/D3S3h4g3a26+Y8lZkMMWK0NkZJ2vNM7IrlMlg+CeVY2f7A0RVQMCH12OGwg8RCFp+66
pZGy34YR/t+3dtDCLXMJTyd6192N7CueNHv5ZC1FHvYqYwX3OfxltMOdRBBQTBJzRP56gZz1FCvK
SXSv+P9dNW9x3rrzkaq0PjpmKjU1pb4ILsy9iUppXuHXRDjR0581QVtLiEV8IGdVj+pmAG1IeBum
REHkoUfyG7VfJyj+jya1zhMM6Vaq5wrgBAKw98Bcq6ICTMUkEmVc9ysqOGNu4c4MkRlI7Un+6iGl
5Sgoje72ituSUOsp0Ckmj1Yl6o+xYQXyT7vVGFQe7MVCCCU1T87z+8LPX7MukP5d/D21zNYJcxP7
7h4aE7w7p6pDP0eyGmd/qE/10GoHx3phYP2aY1SETC1HoRteywxbh5vwNHIUu1dRSEfEKWKdxfhI
Oh5+LC2T3pMheaKEt02Y7bemfv8rKia5S8BFV7rokI8FEnGV85LX4pk5UuT0tfZpqXxDB1enqjWn
F4QrDlbLIxqigKT9e8LpCpY+Ld2jRgQW/cQnNiw32urcnLH0NdISPWRQGe7dxZXL/9Otw8MZrDBY
+zlKT4La4lS3V6MFmh6LPPCOlbx3GNcw2Lli0Mwh0l1TO/yT/OdWpuepSEgvcRRPwTvTRAE8ogGz
UTe1Hm6RSTIuh0h+6STzkxj6FaHU35GKo4NR8c0mOweYFisK0cS1Qd20koYcYdGcEo7GgZmQwnEu
yA1xNIJvwndLSGnEHiyqYmOEOtsZJs9gwLRXotW0RU/udx9UBxwB1q/pAPWhPg4bvkODZQV92N9c
vnQEsBGVOvq42if5cRQqxPv12gMMYXjFG6PSiWToMo7PLm+tkpjN3N3IdhEUhH9x6a6p7ZoVN9vY
QaSy2CHDlW+WFSOag04viIFNTTIUBsSWufajXl1PNDO8l39gJQAjUaQSQUeYItpVaTc0iKrEXOAB
irDwFQTGcFQZFH9+FGxfUkRlDppribh9alMrfuwZjY0n8lNWA83km2StISAgLuZZ93EKupc5ASSt
lr1kXeZ0PDcTPqMZVb5Dznb7KYZyPG0gC5ocQRo3takW/p4r0ceovPX5EBdsJNaMPbu7gOJxpbg3
3WDLIGlBFtWO9FzxlWp0VvHnoLQ8e9bNp8uAWJasulxgO9YGFOGjql033WnH8cEe3x0YHJZqVv/7
6p0sLzShvtW2hXuzBZknd8oNgkH4ff+4jTqrNi8HMHhWM/1gdAPWHYfOpWRejELCoC7pXkozSReu
4S2GDUZnyCDaPVXH4PMexOsZEBSHOme46aBE9VghYOV9fBT7cS/2WB4z9nPQ0GsvhZnTTdQ+vFof
bIH/nZRa7x9OrNMUAdriYKDgDbzDgBubjIFgBz6v8Da9/vr/1VF/il1wEBwSO+ShSQTHKXdfoIE8
DpYaYESZsm/9FwMY+rrR9PwDVRjeuHW9jzENk2sBpNCdKxNAunEaEXszzol1NYPlNKZSZXle0hl1
owcuhUI5feepbcOpJ2kw1S8TCvu+QlEdfeZgmyQASbiuMbkXsE/osuIHp1w2PRw2k+Z3dk2WeImz
tekYd3QI7hSU71AfaxkZaaSzduAIytk4NuQzKtKeZD3KpiHqcbjwxkwpGOOWmxPVaCPNIg6kOGKK
/0gd3p0VP6fR/IZR4Vg+z80oQc7MU4SRvC7PqOGFFtoiAqrK87Tz/xM9S5kTbvksHAPwhlyXQY2F
NFW5usaV9prsR+Uumg4gRX/ITpGtypxOacBmjQc9kH03LKkiNqQoTmVWS0XiQE7wl8RPBRajo2tf
6ACBYqZu23IImeNSQ/G3umh/dRSnXigmwed2Cr0v2IocDfTsa/3OvPwH682Uu61I5wrC21TM4lli
XSFJRCBRUG8mgU3GqKJJf7G2eeFxT/u9QQCVLuIBNotCa+SSXKFahq+HtSDk0lGNIIVjSWJCWfqP
TffvvV4YQCSmyn4Flok8L3WStTmuqWCWP0TvGuDjv30WJMEoSikxmPGqTEqvEiF+9zm1rrwZ818r
eJ8x0hhjcAanJ3slZK6TIE9iUxHHUg08TAGmDCf/QYiFuVTO0lIebjDHWcvIggQuxh3UJ4aFIYrc
mhkkpftNx6Hi/Px7hy6gRZhn5LzCjZ3GBvn5BQGlzJfswAjMLdQ8ECGw28QkmH0NJkg936mRe0eU
yKtZVbOmq4llqhNjyAM7hIc0aD6YxD0667raNBgPMllGNUVQJQrwhGRQQvDR23z2XevJ1x2RmBsC
u8FJXs7WjN/pFB8HtSpB1G0VwF1CpDI3Kyou3vwpcIzIktJG9VbeSBVB+yPitd3LDGz7g+hmGvh3
BtqVDjcYjWyBGQvzIdV1ossGpjWd7xmMK0HpgSXgkchsV3NF0AuAqZPYUG/qA5w2e/R7U3dbs/tg
Jwrv1KuUkeUu0ydU4d/3MZ6a2dhSaBX+I+T9PJiEHctIgHN8YnLtQejEzGlh4UPF6U5RJaMkKIZ6
GcUp4f7zFC5Spwfq1o5sTdGSmZNwU9bQlB52qc8/e2eBp9W0ev8HvplpZyXABHFnYNgoAGkr4egB
TOsV8hRlkzohN7gZPrFaDV2rXWhxebnH5WpezNLLr26L26iFVedwlJlZvyRAq4UI3G6zFHdHPlpE
i6eXCavdt67qANiAUEwNlYbrD6r6DCuWnqaWKRe8fWsnuFYlwc7lzgB6ECUObBI3qtLNvLK9aI0o
oRT+iJF5hm6cdp8iQx0nJg/hAt5rnwlt/5eLgxisS+hmQ13K96UTc8XsgpSYs7u6YhgC3LCAcFXW
gHyEGbdpOHR2HVtlv1M+2+Wog6KPx0+IK72AzdVo6+ucjLJO/EmYuMUUuhvBi2aX/vRqzn7EYoAD
6c5g6s1dI8g2IBOYhb/PmKMFJuWzuBKaIiYbhFrsJCmyA5NEWtt9ZFaWwlFtaL+rPP0GJbSXzjqM
8Jo7K1DZLeQa93wb6InA+kaF+4aXUs9JNMfoWe4ijD3OngvszxElN4kb1yT/DOw3tbHXnPE0BhKF
xf3p/yRvh2aVw+PoZzfduwjteT3h3d7jI6P7aCiH85DhvHAQA4zKrbbtpmF8R2v/QA38fUFF7U3i
73ry05OLtyfRKmXEcpe998eDKiZk+g48pdt6EjG206JHmkEa/nX05d3hHARWJEQLx1i93tl1qEno
J4tLJpRXw0xiGau/t3/vASxIbxRq+M3z43fOx+3FMVqUow+X9K0szbsuklRj8dzOULBDKqll7C+x
/86ayn01BjtqTq84ZRMexIGvLU9VsvtA6Ehem/0WAuTkwIVWBV4ReACssb13S/dGuxqOtkVqJZtJ
k12+/S/fFFuEse9n+jqOtfmIHVrAa/1QWlFCqXpKHJ2SacCaGomOpAluGCebE75Ly+iVbUKcRlU9
jgGPW27o6O3srAp26WkxtNJGindqasPjoJkId4vHrjxzG0DCwNElrBr25KWtcpiALzokdaI1yBXp
iJ6rkZm5Wc/gdnFQBYkQO6gLwxd6T1V53IhB4A1AeL4kyeFSqqXyNMJLPLnfyqntF/LkzML9tV2G
JElIhFLiEZYC8CL14OVeMHlGNPp/nD/h+y5ZjQvg0+28U5skg6YeuxbZtEL3lX/gf9ABVb0QBXXg
f+55pNdNXoV0e4GQ1zRGGU8s9I+pCumPg9ldrgd651JItBwgdrF9sMwjKP4UhEPuou/uvPPbJaih
t9QrWX7Xc8ayBOfxGNX54Skt2gUYgM3RRAQfud6gFNsx3kL1eVSQ17F5TxoBQ8FMxk4fGIQ/UnrN
5FVmalJ3TwfsRy2/qUBUC0K+B/dRR7sNIPP/z6yUWsuTWjMcG11IynH9fJr/l05a5uPkiIediDBO
1cTmyQtfIYWUknCy8Cy9aO5Pdmj+215evlBby6b4SvPo2nqy8Jiflonh+kaX7Z+noFk6WZIpQ5GV
U0D4qckeavG8CWXhfWZw2/d8SAYVZJWUo0nTAIJFrTMC5IcOF6+avXz+Rhj5CAKF+yS4xKN7XUvi
eJpa0ORSMrfOZmPrTwtrGTBsxTQT5puNCXSOzeUNOPh7ngUfs/l3LGG+W45L2X6Q6vVGFdfMUoOe
G0V5oJSPHLnO+Q6L+s/Y12azE2YBO/ey6e4zv/URmgBLhR6/kT+h5ebKJoNA7vVYLkkarjaL58Gk
O8h4HHBqKghZlEOkZdKdebDmqTTXa9WPgROifLrKPtC/um4DW/TbnBndX/1Prz5a8WUUPf6WF0LE
LAQc0g+us8BWCmSJu5HblzIs6eGZjDRCFBRDIUfZTobPBQxYTRNCSdOVcf6MqK8UuplMjoyWrLrS
RTPIxcSuARqUBbOQ3JtZaReJTmL+dFa7jYKhBbQxzHG9mAyvhCtaxbdQbwX32bVXrPshPWcBb/X/
dPvOveAowSrcdd+rAdQtjCO1IfAd8h9dXn01tHOutsnd9wv2i6WJL9jK+rsLISWmXrPJ0oYQ90gm
IQmY7IKwPoVtD9QdyLizcTPBOouQJ1kOfgj10KFouCiIeulW8X560HJK6kAIwjZU67zarXsmTeJ/
SLPTBXTfn2pByAPe1lM3j8cS6NTQyVocgsSMKOH9PlbIqWlcJRqdzUblhAKxvbEdRRH+h5YplA+W
7cZF//au7luy00ZNFtwGdPnPlCr/28OHgJYvB97uiSPwsD41dEdYIKYqXJ5Ri3/Obitawe7Xp19k
XJdZw0FXmsl0VIt8ud7MLeQgLfTslw95rgTGu1PKLjHLfu3HRTRLP64LZU4qPpP80EwRySlpJQK0
ID/hxiTC7dZrZ5MOjCO0WEl870wZW7IlpKVAdtzbSfbRivVFNFeUrxowi3GvuudN8Blhbr72cnIM
pM3Mwfnt1XWL7wS9KHrYXhoTivgE3UNNVCVNrwlC+osL+V8SWYebIWzgFBae5iMBMokywBA9TxHy
ISs/m11qx5t0b5C59SxWshjMrtf3C5GoCbAL961pW6PanlO5Y4Yhj279sMVcri2+i1aq+gBrNJyN
vAQkbxsmremjrBitn2k/uWEENd3yx0TPe0BnrOXIw9I1gpL4IV9nfFif+hjT1aajqP5Dr5PiULZH
cVDUpieg2f8SOjN/nvU7ZC4lAFIMLGvdi59uik0d2c0oXaOIXy2x+b99SF5loUJiYTWENlNZTHyJ
ChvMOmr5K71Mm/wdfId6cH46l8foLzIVarziggEA2HaOOw8wBDG6ljm7/S9ozgPfky0XBzVgKPsV
u0L7/15GWDgyOReP0Nsj4RnKLtleV8DQUvFtEo/K1zyJoscGYyMdlV8OOMrwB8yoYqmspjCn2uVM
FiFRrJW+znGiIOZ6zB5gHROZoKhE5i9pNRsrJp2dxqmRdt5wjmxXZNZHOemXzXg9UJPhd4hMdpz3
ZRF6go3rfDNJVLPaKAFvY4DB0cZVJubviBh3HxCacM3kXx04VB+ChK1fNAHuIStnamLEE6kblrGV
njXDve3f5qxqQfoeTzG4tNWsmIYjIQBNAKBsb8q6LKh/PX8ZEr8RK8jUSkQF+DubuMPB5Muka87t
g7ptsOKPee9pWxiqmWbNJdENUjh2H03mnB3OOz3ynCp15X+TfOO5hxPNnOFoP0CxtbW3miIGG2Oe
QbX7QMFTK0aViyP60z9mZbomNA753FrqpU16TI9t5khRQzwiFVMyDeoLf7HcROU7fDsolT70FnTQ
NjG77qAF/tGqPebeK2hMt8+f2kE3wz2ae5BBiXntW9iAIQhCgjZeDYwkiEpgg2kQ4UBrWHBMciek
HC203QaP2VgjIrxZBt9RFtfI/8bAtS80Yr64TM2X3sqaHw84vdNtPtTMWmFanAftyZCiVh8H0Q6s
ytm40yCQ3HpQMZX641ETqh3A2moN9anHp4qz84QAORTiOL7HxT/D6J9HTrarWiEAtjgl4rwrlbVz
5RIX6n8ZknrkdTqaIQGxFgUj2hkDO1vtVHkTyvQH4sVrz1/LzDEFK6tSoUlEDMXmgcECLHLI3BWh
jZ1NNWAkFGDgzpiaaLTjgIFxgOp5lINoyvJO1H7zh5zausmRiQ0nlpGYEk+2ZMnI4buW6mt+ISBh
wI2vGDEDBcJ8nPjUxern40vQf3UwekfqOG11CDJIjp+QkKNpB3/NW3H/OM87xkzccL5x/tzZ4g9m
TRR0crC/AHWI6mw9VVc+B2+U3gXE/ab25Jfs+XvxhqBHCFujKxe3h1H48olGFDJUMUkRON4perE8
329/v9pSw0viWmHR8hSZMBRRGUqkbsqhF+RgL4FkXSgBwusEzI5hFIkIurkEj7T1yU/VLchVuITa
3Wx4WbaqrPxEnQF2cIgic7GrUOswDhIpurph4qPQoDShxO2T/Zns+aake2v/6PBBqzwYhNiCwl8u
owAPzEE1ycEBkPeUgM0eICVRKo/3b9MKgKoWlB+xFUY5etXus9+w9voalkw4CoUsYaXNwF2h/pmE
JFTkJRz1di0EYFaT3PwrVTUsxSduqMz2lxml34ziBE0usJamQqTXJ02WupvnrPXiPTGp7ePkP9u3
a2FBxnXnarpyVjo4ekM2pHwM9ksb+o9plm+f+QGcSkkR+3mm1NbctDZgP6SMiRNFCOtT/lUQTdi9
VMxQ7f0z44uBWblsG2F32k931VWajQyVRHbHHjgJJ1D25j//z9Tl4NX43FzUyw+Zh+S4xqopTv6Q
8M9mUaAi2TRhOwGepmVdlrBja6bhHWVjKJzQNU9tH0u3MXnsEOCPAAfpiWxdgJbSZE5xe1hAKL/l
YylTZe+R17DLOdPqye3XnRGPlOv2OZmrxakA0Q3t6nWW/nCAY8e8fs+7AngDQsVO3W0zEyyr9aCd
1rjs60IemETnXTHBr/MBbyeuJYeP0uVt8Ptl44Zr++RE33mFJOTeVJyd5kRMIJyiKA36XPSWniE5
U7lqWHezXyox9PLq9zzPNqGaapZaMKFutOXXAg3j6YLD7skD755qajsMSPCOn+RFXhw0iLB9TWyN
TDecrMMT7KRZPQy//Cab2Ce5inWgXYoN3J4fJjHYymXBzfgjic0KPY0KEz3+20kuLM8HPNEuwL+Z
2pAcxt1u0LRGCK61a4PkUWQvmMk7FU1iDjYXpAw4NMQ9tCjBidk2v1Kj9vZP6+31Y86IAj9HvH1A
wmpJUxhsWOh2dP4RQ4vjAR6dVkERsIXnbWB1OCmsmLuI6kY/hqSLFqwKLHLbpSJsB3/ST2FIQwfU
ISd3cy+2T2wAhLWJ2C0WzpGaWqgAlpGYSPMeJOMBmvD5cgkjQ0GH4LTaBZSEnbgSyc5jtonAVD/P
yo6KuhfZwwsxzYCFJ7Y1lWhpwHAGXNC3VIb0/NCuUcdkM12jor9pqR7XtIF0LatFlzTwQVZxHJ2x
Sgeipu8FUANneVuYQQCUC5N/wTNQ9vBnvpro1gUXw8kjYV6+F4wyBEJneC6WOnxFmZBVrPf2zrJE
7ztrOeFSqDAXt+F1XF8Etvus0jH1zqK3n3T2xXWu3YMgwFv3tAsoa3M32XTjqqhvlewJTTi3SiAb
RrjZaPpl1GpeeX/yfpCOjE1zIVV25xbhgawIGV+v0py5kHnEC2WHptTt5/J0L+jWq1iu5WaGKkqe
0m0LN1117k6at01tdR9KzIsOAX5bdd7Qr3ANsYr9th8ydQgyr9NtI4zWFV/uW1SV2Xl9P3xaS8eO
e0BhSbG927w/sdpSjwXPIBQBkE412iOc5PNCPDDd3n8auWxQFpk9BxRkwRdPvNkgA6hBbUQKcrXx
o7oukj/VZZS+/9gTCKtYXBB+DnNwh4SjK9zbTdLNcmCQ9KP2xPujNQjgzrLqKhIlpI65do0kSmgW
HBokqnEuI9EhdLSL+PJP1LhC3PuxgbVkFhi9GK0bqiaK5p5GJiMo1GecImlqRGCCmOYY7LkLhdPA
HULYrHzwYX+JBOV8uFFSzQ1N/u+HnwbiHx2G1JNErd+AieJbVhzApR6sFh185/W2+CVLPqX285rG
qNbbZsf52OZg99D68dqLU4/B1coLGeYwu6J9uIspXq47Lf3JNFOvOtLWzlPShtxAPq0POAu3pSZo
eDQw/nQWhx57ch/RTE3AOodqjAOL7q5FBLkH2tIIzmvWEywnGZMLuLZ8x0oZI0fQWdSR7f0ka/4R
5SVgLOwoeO2CyvE2EpFHr8mZfJ90Pm6txs1Gk/2Sgi7O2UtsHdf3aQxUMiMvPljtN2PmFo0KpdIz
5ooYaajFOfMQWuv5QHW0YITcWosfA4u0smbbHJcP3/61Mt1JE2ggZp9rRbfnM3L3fPycO8pzSbmd
kiS2L1AZrngcJ0wTX3Tb/YlK5++7nyAOvn+pRY0f3guPW+8uNVtsjGixt1G9W8Iv2UFlF5y7LOI4
P7WWfGKwl4efvhx6rwjer/7G/htZZdilxsSK0WXzmbDet96KF88/0pFgj9yqrZAZLBf0Jc3TEIWY
40ujOv/ZwAYf5NuvwEWUFvATPTMbbGoYrGsno2WBa4fsBlAQI10/Tuhv0t0zk8ROmzhS/wPhl4ew
QOqKb2LqKxHEfF6PqE73bEs1dElE053PmLAlOwAcO+0tpNSz724IHgKbze7jQmq0Pt0vCAPZgbUz
af6esrvS0X9A3me+p9SUV0DEpOOTmIRMNuJTBghhUldW5IYYFwEsgAvK6tttQHns44F4BIG4qwh8
HmhW06nqbCDhsip/ilAP3r2i5dtsJvxoCX4cnWdTAb/8L1UC56lXWhmuGLkDHb1qrp16VOGZRL3+
aKE9WWD9FvV8uIP7Fz/nh3XhSs9GIVbzf/vaCvmPrRGCw9GmyJAN+ylxg09cb3KQFriHjGJWy0OQ
8HYUP2QlZsXFcE9q1KZj4V8akORMPcyNx+6hPIDawYUg/qNd+hF6wam9x9akgdgSIbQFuNMqzjL9
Dj7yIgmysM3jCq9UGcCZSmhhUpZ6J3Poyca5DKTrECo7FIhHAe3xcyGG8QRWXIpD6RNirblJtFq9
jPqx8X05HjOZMA7xfNV4bO6wDVqXsUeGgugWtbkzZzIDTtwmbvmZPYBj5/EHprUMzVaUYjT+kwRF
EA2CnmAIQXDblmGy1//28PFOL99QhcMRSHtmahA6Bm3zQnMKmTqV1pNzbGxKcFzb9NUlbwMYrm94
775THrY4uB+VyBsl7nEiishppLi3WHnpGGYcOgHxCNwv3z/NbR1A0EcrHCK/D+c9skJtfjpCw5O8
P89yhcHsjrrmf0uBXmVxIvMiiaPwjY4MpDTQND1sTHZDoN8vRr/aMM924t/GuuUu0CobpG4Y+7Q7
Tmjo/eE3hKGCY49+X5ufOr71XkktKzjMqAE6W1+gg8aLRUMWzalymKZykoXstTE5ogly0ab6Wncg
MLQ+V9TfHlN6oQwqg3dsviYPpTaPURLMhh0Pheu8Phlfrs19gZdJL5l8F8XsyZBMNA0FSK0VL6sK
dYQstxiRfDkyFFxfIO6nkb2i50tq3/tXw7u58li982xUNZowRM5+WPRcnq5f1m8SU5uT3fxpPA4P
5uNcrr4mOAxGBLJqNUm137EFNDsnhNgKyWP5UkQtL+mpizg8GyWCEtyZhjx7h8xP43MS46NI4pFM
c49lmAeA1JbM+6jsNSxIa5GunnSnG25laRhPCVpmvE6EyJX6QOKIRkO8v3b/mzaUKaqUBaiXCd3Y
eMnlDrA2Gd/aBEAHc47Er896ORc97rzyROgTcFs14qzezeIng2TXIpQobEZHyKTrqwyYbWKEYWzM
Nsu9TFn5KmwyeKMVxxIxyYhdRuIX8D4AbA1eI+AeP7Wz70edIlznEoH6tAofJFT7JpwRCHm40z16
WpkslbgVVBGu9w6BaE7LaJ26mBU38MnYMMf4Falmy5uYQErY9pkbgZTHg94xtAVWMtsj0N9vp5Uz
bmWl4Lu0tDEHnHlU9N3b6qAjT5JMgCasYxuwzROue3+ceFmxOUA8qfYiLhwWKp0UHM6sTXyt1D1d
of4npKDodv7VJko0WDXECA7gZbGGNK/HHy6tDmm+UmMFKLkE2u/cOu+R/ItFPmAFEgwD7vPJ/kWr
Ij8Sx7N0kumRh4I/vhR23GZlqaQ7D18ot1ovJjSq3fbZWj+CgAm+aaxcGqnBCxULc7luuSSzayTI
ddNtGGIwgdlXCe30Sf7Si8iXUQq3JPmmocxtESRavEZceRMyhU15ZC2wUL2U/CpNllWm61PyL/8P
s/ch5sc4i/F61mCFCLdavzfgf37SiwvIvKbW1dPx0vbSr9yKKwYunJAYXPySJnlghT/zEqilZczU
6Fy045DNSU7/72b8/oIG5D4KYbSTsCcEjBs61hsJoTLA7NK62xRKoePhdD/pb3VnIuxpYqs4Pg9w
GLKZ0iQ4sIlHIsGGV8U7pboMp8KI1kZdxAUfnsqS65Nv/h0opBsUkx9Fc82JRgvVtpDFjOm7HWRi
WBAv4egU/5p936CZYht1KbFyaRMB/blrXZAxeJbwOxs+cmTZ5TnSkAhKrb4c7t4I6w1NaXnvEhj5
oCjeSh1cXRVsJv6jLUYu1VMrZMLqIuptKKMa4O6sQadFqaetgcDBctMJOgnCog7lszY/U8GqTP81
qNkFAZVjRPYPw+Pu44Mn2EcSXI8R+Pc8uAt1F3glJOqk3u7EVchcb5g6FuySZxVEGQV+o0JNcN2z
75yY4ofNiUoc7pp5Tbg5C7KUu8dOE9GiE+Hadzqm90g3t2GxI2NwmLSo6iMcrMyCnoJHWs3KoMfe
arMrYQLEddv06aX/kX/oR7o2/9zhDzn3deCHXWNKZhCUKYojou5AXMNxa+is/OHDQcZPCHocqkoy
m+us1nuFl85D40rq+U9R8lv/D0MVPt70DbrEWq6ctOJCevnMouGnRqywvDP1lNHGSc22TtunBTnN
yf7u68FiogPi/i+u7nL+vFCFzzsxFX/LAw7+ZAlTNBd38NocRhwSU51KDUoTPm3xTH16o1nXGF+C
ttqV+i1z8z2oVF3HsuDMZwB+OqZmeC4HK+cERF6svTjheacIH9E+qE8YxG461naSXuqr6roWuX4H
nWScVrkQj+NqnGlnq3Y74xb8HysFCqDPpxkf8oNMKKpD5T1pIV7uV/Wh8MJ7opt8vX4aoeKUfuqT
x1p8svdfSpvQmxRWasXHrx/YuFugLbIEoDGnh12gw8INfPJFpeOKBEBgHO7NiIHJHDMOzojK26XA
NuUNZ5JZao1Qtkmab7ZHS9gN2cF/lSTtR0LZOvAwz6WBgaAC6zzaUWptYa5Q5PbIcMB943Q65/uE
R7DTWUet3/V21tcGA5N1sHd+CZb/jVBmxK03qai+P2GTgt4Ml1JVjWLlu0lJEm3WjwE/NozvPhKF
362Nw84I4hrOjMAeU0Q0p3PcdAWfS6kzeeGMdlT/fcp5WeSLeSLjOV9x60Sym/XfZznB3u+NITIU
xQ9j50UqEy5NwiFXHSZrhZApZWA0kWR/vMXbC2b14yq5KLXXhVg7eXKnYi4s7V8bnmzU0Vg0CDUa
vZv3YloIbzVsDzPvIUMFI5PKW9cc7f7hCjTNcEM1M4z6a2TfGLW3+69FQGW4lZV6a6KZxRBM/7Oh
bSiLaU4Ty7eMTis3rmVJ0uWrOh7nB1rL+dnU19QG6+aReXNVLnkfgjBQBbLBlIph0moQuBMv5Z8e
8OEdF1HqgcgP8FaOCDYSoEKpLokYKwvSxkEp/WsDk/issNJvb/G/8iVFQSR/bEe+mR6YVRA+IcqM
xP2xzTTloaN/s+KfmMHkNDOFXvFGhd6suiL2/NePHA5IQJugOTjmZkXYMqInO4ItYYJMkE/cY7lX
sMYlIYouLxLj/RpadQRbxAxO0e1DlGgw9v5mgeisew5RperedMXQDe/OG7xSeun758Pr+ps2AlPb
bCIKHoehz5CxlafadDWZrG3IIp8Jf9/hXty47ie5DJA3WA2wSuUCX7dp68rDZaDADlT6ttFV0rp7
GADXAYVThKqPPDiX0R+r3X0ApRCsMwzWxIbUjrHbsD23SvwVP2o9OUF8G3OrlimKUJ8cfrN3m6Ek
9DkaLQHXlM2MB82BlCHxfzJPeNOSeGl6VTxyjh+sy4X8hf2XyclEtk7FrUoQVUM/LU6WAX2k6JlP
ibDsprx55sIirtU2Hq9k8FlzmZNcsGQfLb5kwiVbxPJLgCl7G6IDXZJEbf+mpOYAgYH+fSdBSVJq
b+4wp/P34F7+Z/akwPhrTnFTbzoyg7q87zgyvcLpvFdH5u0PJ67QCrv66cq7mN6LnMdyd7G0C02l
4Nykph+YoJ1ApSfnY+k+poi9vvHMLQ+qmmu3K/W+hIL2zbAojLofVmOdfyzIcz+GNE1HMqlQ2gfz
5i8MFR8BOGZFteeKLBh25d1b7pI8g8ssWDL6jissIJYzNW/05xAQJQm7FAKWfZPGJk8P/aMujSTi
RzRrVtOqdlWAvi4moXNeGPxZLB50BzHjsRpe9suD8vuEeeRxo1Su2he5rf9XSL4pir7r3yELq9af
6HzhRnLDyGLZNZtTyaISfZYgEDCMVteHe5HDWaVB4G3DIW8JfawsF8xHnkJo2RUzrm6jO6s2Ipok
wreTK+30x0EhmFX70rJCDK8uQlO0AuzoKKuKZtFZFZ7E8hehpAhzHg4IgjZ5wl0m9kBDjagNU90Q
NR/7E9Ix4B1hD4YD5/pTax+AWHtDJmTQVuvq11HzZIOs1fY9Glhz5zMdWAfCQqksWKL5Qz2VTUeO
S+rwlGSbIZxQHGkccASNIV19yv9cJ6NBRh4fL2xKB26XOuNub4OrYWdZnuJyc+kSh8zj3LKyNn2j
J7yv3egYQuipAsZTD1WfNfv0GgvwDAqxa5Q8KvWSmS9/CxkPLaHjZrtaoYAFms873GoYS0RFS3en
QtCsLPpfSETYQ8W/qwIE0WSaLuCzqTFjv/Aao5DQon8t+TpSC0NdqOv/hVKLhgRxS4JThQdKTgiW
rK8Zgp/L+P8AJyhC7IaWVoPwxAW7fvjyiCwVgtyhHZidw/GkSh6XuN+niiydiU2Qk0N0EM1uFtt2
0jAaDRXHkQC7iNvWr+09KZXxTmZrU+i0/PQBk07BYfoQjcXF07IKEkD4VUlptanCXHeWh5rO/DZE
Q/RzFG6j4qgnpSKc095WQ7aGjGb6BQFnJ+XhaG7xxnppR97V4FIMsYMsvkEmv/36KjrSMRsc6E4f
b15o+NUgDYufM5grqTDm39/GeCRkGIYRXeJV6i75DiyWuul2vORCqaoAsujwbnkKbC5b86JEccuB
5MAdoVLQw/nyV3/eI9NxzsVjE2I2rY88VpKjWkoQbCTcnBDFMyrjWd5bOMu7Q+7pJmGJKeimSVbn
5PXScVXlYKZoO0Nf/96uKp2pgnKwc32Q+Dempp7eg18iUNUYmM/nNBokGvWl3jrFL29Xqe6myYDc
2it9zFbuiiKbtF4CbRL7Cya8eBkwYW41BhCUEbryTIuYtt/azcPLa1z57G+CJfU/xSiZmAW2Aysc
nsO2Reb0R9r/2ocXZsTTf6awitg20drU15FG9YIbhPO7uLyJAGSvhQozXUrmBFn4Lq3j8vjcaUjv
jE2DK0oljCCXOlSlSYvIfz2OSYCM9uLAAxKIpOWHtjQNpOsdWpox9r8CZFQsxP4NCJAJw7qtIMRY
7hiHFvTdSdEYKgx5bkjN7VMbCxTlCESfE+p5rrHr0dUequv7wlcxT9wrdwC9MF1dwht5XLgsP06O
au4TQB1kyAKT2pd3xnUhe5+A88QTgJFDXPP4nJwURzDdgjr0ZVGHSjayHNFqKmOfXlfB8ZnpD/s0
GXLaSS5txzaRjN9EnTSaXXkMBWU3tD20eo7mp1rkOEm7VPkh3Mlh1db6n+TUrZbR/uzrxB5pVo+f
AkLBEDSrbjZP+BtAr35aKV3lNmhOc5yDDukHnvoMJuk3Z2u6neclo4XWkOjaSU4mVKgl0LqBV3Sc
rsXed/DHcCiyWGLi3VLjz7khE/Uai3gLwAD/rCyy38WEm0pH7x5dtw18o+m+zYlbD8lnipUaBpvd
dq+nvkqaNjh/JWfZMu1C5WvUupWgWLYNvJ5SCfQy0k1uc+g6Q9af12RmTYtPqJjrlq3ohRYId4aH
1xR2DvSOejqHJbKDOLLJWs7xLUHpxpIKL1Y3fmYl2W1zW+91dlFPmTBVE8mgsxy7biw6S/yF5ziw
PsemMi6gmZHoqZrODnG3IA3rmBdHwduQIGTIINCOrKVTPDtBbE151Visd6Uy1kEvkGEtbICKvmrU
G7WDNrAP4iwXMAKOnSd8SyKIf8EgcL68tEN9gUPMTNRBIQYWqP6VyBbLVNp8bAGAnmCrJt6oRle7
gp/8gMEPBqJfQhoIs8gK64xf5vjMeb8el+NDpcGL04qaCqOOu4Nckog7WSVQSpLm5GYsCYPJuPC3
s37uEDSZI1ZcXTb5aIBEQqrMfBvPg05AksY8XtplOJ/3EvdYyhsAHDhvtGKAC8QVaTPQVBMAXz7m
rted2T6LbhM6Dd6l1eBFCBR0wWwZyxBRigkE0HOdVdUjbhR+lu8/rYyHLnXclre7+GqGVD3cpeaa
8vqEzPodgTAIOHWdilehL/j61JOyhpVP8XPxc3ecRoxagmPpO+DzHPUEjDRFWig06r/FolqqUsf6
Nqw1iZJjVynalC3k78qVxR3hgUnki8UKjHS9AB1xdlJQki+P76IR54T3oS00j5Qt9DrdYY7ktr5W
96c/F9l8aAFqsLznkyDh2D2zzz9J87KD/ySbjB+c9WEDzK/tdVN2gq0py96HM1zfC5h7pZM13Uqv
it/btw70zSv1T5hZiBXFtBBFN68Kwy3JLLYCuUo41AzGqPp56DsnYYqb9euk8oqeVXi6yzBL0Z2Y
UF1G06YczIdltawzdhPQUdUPMCXnRcQngL5CbK21QetNle8DzY9RKS+xYMRTddyp7x8FUWu9fDLt
iRDtlgNmPCJh1sZWCLefmHz0L0n1ukekZk4jKtSfDxJyzZ6icvxdsDptCZNceeInESFipk244Ay+
KS4zr6Ow3wqpKHbzTwsQeeuMwFbSUEm9SHatG+3oy/4AQTAaN9uFM6frHHIKiE5xaX+M1BPkocLH
0xPYLSVFvGAFmAQ0i82PAKD/nF4BffkhPe5+Hnup9ER8TWLcH+kNHpmUkuc6j/REmlNlU/myftLv
F5SbbPLIIC0Y2/tuj+btWRyy7BXTAjTi9gTHyzzmlcas9WAROsNpMfjW/6z3JOPUeUUtBoqjEHnU
Owm1bcC9O4zd2OXtyD7b9ajbBH2tu6U3Mw9gYznq0NOj4xqfDvpKSBd9OnldlRWffGwpNKxVeuy+
f4Aca0Zr7H4sjjn2YvYwo55vMSqCIfea0ncticbRF/hnuRqhrH/nFFtjvz2aM6zpU5Cd3peFZ2cF
ZDrM+dtQYsr0sdsLv/zEzxC5BhmUt/z+AwEKedCGO4wV0wI0nZzCRvpFTIgojYVN/0Ubyo60Rk7J
zWf55W0CNUzT8HmHX+CxBWDNVWmO3yIGgq6l9/dXVDisHUwroC55WfxUbCbp/677ZgT37vzF8a1T
+8F4PhntxMqO17uGkVK/6xNCOj8UuEsUj3cpq282+rsqj8zxOBqn7rKUdOE/FZ6fWHCfG5NU8Dn7
eMLjZZdG9GeFEYUCLTO2L4UT5fxQWVEpCD5gT2HLvsqWSkJ1bayWXsLSnMlbfDOq5AfVhDKT0NeH
7bBwsXHLAfhMwPm7pWW1Irk1NGxZ2JC3k35+uqR1ZJJqAoM0eCBZrbCiOTCVjMJY4w4VH9wUA8JT
Lt6r+6XEs1gunuOmFekJsB9Q8H70SES8OGMOjs5NaX2ox5BTBIAO2dluRo4i6Sxij76G+D/L1ThL
0vTOLnKp3sIv1U6WtM07OFhdtQlbWXBGmr9p2f+GfqpxqPBIQyiCzYRb1Lc10cPNdh4dXtfHJKEU
EeRCQ6L8/uv7QOli+qqciE7e8Ep4BhiSrQNPxOchSOjcpk1bUMGiugSDeV5Ff9BDJos3lkqLpFIB
sMzC1UQNNl6MAyzLLPgUoPIl8uzELwUdxFzlHQhBuAdJXibLERGMgpfGNEDkIRUDtaAJ5fSTD/NY
xuWJydvWnzdr0PNKycOTMfAPITFXAG6QPZmuIRVfP51dCqpJwRJ0pusdMjjLOvJBKzlH5yY8m6Dy
NoKTnnvQhikzSwbmVSxIG9GyVw9BMQ6k+m74gqxtPavU7WHGEh2bLP3qeLhJOlYeTAgcnpT2waMe
FYNxVEVG4iliICmntyrTWztIqJztFkvMUKAA8hO5aaaUdKbkkYT9Yyj916DlyL/hixmRzWwm2r8F
hwqxpcqi/xVWtfBvj7Odi/xEqC//QrDVt+KAu66dUWLQxQ3lHD2s7b3zelmMRvquoDvfLPzLhPLI
DjtM5jcx5LLkOCNnzupH7FfhplkVsa0Z3cV4tsZyDBI+LOfj5eyX+QeIdpp4GfQjp953k+4HsgRp
QO168AuUqvPFzTlLoxfxgXYaYKyN4XdLi5X/Wl6L0Zt5No43SV9dMsrQibWOhslg0A/a/9US0K+Y
AxI6VH1W9IfNs3bNqESNuEBALn1Ye5uIXGTPLGu4z0oY0KTT/DnInXfsEpb4O/hnEuLCR7GJAoq8
nXk7heoj8WBFkn+HZLCozMnoSxUUHMG+FPmRIVUVN0iTvtyNNLz39k9isl/NGIrp1Yijt0gdsQns
JLnVFyLemMU44QmS3FxRrokS1QT2fHgfqiwaaR1sfJDk3S/ZBpgo/cmsF6V7G3SbTFwrztGfclT/
w3wSjYuX9YW3n0dr2fbnP7vgq7JzerQzyDvk8AM0JMUnXpHo3HUi8CS6r3ACxODFm528WIUKM24i
8NF0buVtCd1FFESI5uQngYMfJydGMLjorzzVoaNbbFUQwEViGCURFAf/k0pxDdJ8uto00qjHSMSm
ZNwseR5A7QD0iayijm9C0bChFKC6gb8TGz6kv4CEPb/F1QQI8HjZPht6II/m7v8nY9LNgr5mud4m
tUyePw7EI1BtiswgPCAXyR2KcitSYaXL/wAoOWS1wCZuBxZSZZL2Z0rFLv5faMR1dpR0zT/fSTxF
Tl+wnz0tEa8ZxeTJd4oFWRVLf7cSnjr5sJIOsK//vq3WFruzebcUf40R4xrRDKV+OOGpfIKHnx9R
N3RZzo4/znAOj1CLIKWdyvjbI6KoxgDMuk9Q5xgqM4PhWCxekDVoBrhCbtUPKj/MsKmkr8P9WXVP
PMmJl3FpEPDqoyzCE9Y1VUO8NzDTLUDs3GsbA4vJlsTXMLe17d9gStQs/eL6resElkhR+I9r+O5i
ryALZRtZNmCxnA8oyAiOYCGYM+GuFRF21JOUjKlqQZ57jmziK9dSdnYcdbU4nxsPa98YsIIs7tMU
C6/F+VuvBhSitHllYwVsfm9woFZ1hFH4FBq1HFIPR4aJP6AhmRHQJeClSa6Qc9pnjYJ8EWWctQZ8
MueaS8FotACei+CPmNF8/Y0WgnjYmSafvrZ9+u8/n2Cj/E+b1l1c9mtE3XfjHZoE1RvLPUv5tv0s
/vdCH1Lo0yd9Xx/zE+tZBSbSNOxqjg2hIk7Exs+Svve3/L83kCbVdBm49S0vWhysA0W8k+m3CCmE
HQyrizmqIJrcqbTnwnBisD08pBren6K+ERW4mIejbbUra0f0fa3xWaMdCuiwggyOVcvRfbiuPpQg
tzKj4qC/elMqa1pJIRd9Whme/efoL/8RnGEVo35B1QB06ctn+S7K4RC+ywO9D5hl8NCJyLbPGrTE
pJaiIGh6ZlhQmivNwpKwGTum8DqM+vPOpXsrBAHo5TMehbSP22tm28+JRZQaNUjnI2C9I1NGfRoC
DbP/bwwTG2JNzBJaGRk6cTJ1lOjtudJAh/ZydkXkzQQmCG/e5TCTjbRtxJM+12OLV/ScmFtv3Yhv
vd4SCqFv34cl+P6oJ40d/YbmJuAlSSKzvaz6BDKDMHmnEBrji/Pw85Dn09LP3NprMaI2EeQRN7Iv
2SP6FweTrsSAijVU8yn+9n6eYD8EanapcpLWH0thW7oHooUgMd6qNzcQj+uFDJU1EB4kyhdjMeko
jkO8LwA8JKxyr3rtK/yGfn4mqDGi3kIKySIBBYcRckONhSWTDgffk7eWql1eYnRqVK0OZiKMn3+r
XPWbYgYZ+rjsBjMtXdQ8cyMYOE9TNTYdsKjHW4p8quc2vNDTiHyJxGLTIb/qEP0WUI8WwGvasNQ8
GyyR7ukoNEIl2Q3xPMDnbTIzlj9FEQsC06AMPPqMaHY2LCt1nRqiFB406Vn6y23iCWym0yRPE+NU
iDePYaM1vs90oOaaG4c7I5WVZLBmOTIa3WXcckkD5hftVPxlhg7Jf7ZbqKlfTYJCyWqJtrTeeIqf
qLnCBYVZ9AbRYCZ+3WnKfVII0OklmOwqTE2yAko3ZXn+VuypNt+TNdL+4V/EBgKCalpWTmb50JCw
a86RP7hryb4S6Ay0t5wsbHSQ/EoYKYnKZzZ7FU0gQyZaczElZNnIVuDTR8FjDf2sckXvsufrcA+o
uiwP8wqpoqCh3fvjN6I2KyiovesMl+eUxxy5e0T8SXnLGh+giAVJ4L4NOtMJykfJNtX1bogsP3GR
aFHZAvigz/NY66WrbpKPvh3nrF90+8Ic778Ou7ZYVsV9dVBoDG7rgFRkxkPlwVd9H9J8VQXwqskE
y+OCUfomT399voX8hL/Xaiaf333RblZha4JzKWVd1Wz+YQiDd7/fZ+SZ8qnVfPbzj+YyTy4UbNdS
ef1qpp1kZql5bZWUyWN73nXM9/O65r2KoH1blgPeUdT9eMccudlyIehv4LUMq8i6ZuK4e4qkrHmS
2hXZMqNYVdyWepuUx7AAgzTzmP3LpZzu3JZysP/uCcEk1HMLAp7VtTkJe/i917QA5px6iq93s5fW
1FaZOfZCwjAGSmtVIfLT5gGueboX6fyBs+8U+olJAxtaiGBTYyGFiJqvGDOZ4tN9gAq9V53HZUBr
5EfU0BmJKdUGYut+718CWPMKmcp3qVn0ZERSiPvjXdDO4BNw21rhctyKnQ6rnb9OJJQZIZCAU01j
DLp5/zgddyob8DIbnSAJC3LgUH3eLGXiBlL+zjbO9D+IL9boH2RZwVwcvq8qaVtb0b4cbjYMRjRP
qU3VJIeyVMqnb/KHrzAJtjw5N3vub0562/hnAiI5ic1MqsWPemPeP9NbZFHLk38FjVhdvWxhaL+X
LI8caMyh6jlVLABHNVCT+SpLPSuxkNXUd7grILWRDRUvDFaedkxtqL7k8AbnXabaR1qo4uqlGE4a
j8h89+0qFc8uUw+6rcknuli8mXxsOu+4qJNp+NOfM47VEBIoAf7MNlTANpRKK8Uw1/RpuUJFAPdy
IQbGtaX2MNOk5JRv1vzIHrNTDDsk5fJsKm0k8hnk67eoSeCXFX2iHHvDc0fEQCECohtp+3HKH4dz
yvaicmazu9aHVcd0VojyXFNdTWU1FLOaN9lya2V9/2zUqkQrSbhsaC8dkFGOX2euF1LZaiZNYghb
ekP0E29zSEU/Kmjgd8jiTfi5EinnQwT7Rwbz82gxwY6dO1+TS/3Dv2Kr42IjymtHMfWYNSdT3lmS
+Y9AYoH3bwd1TecXtG6O9+aPBzJhUj1uiPiP8KX/6VH5ZWIwlnyIhRie00mkWz1ktNnLg/siFfHC
Mn/N3j5WozjiM1OTY57R+3ZnDzMvsFcoYF2T4ewPBlV1g4QPuT2VAh7GnInuBQPqUnFjMifoxDFI
UC+ZRFkqU5vYKpVpqSIsrU/8+lktP7pOf0CgfJLWLpIJUSQ2oywCIWFAWTVu0mdUMomnEi3BoFEP
QB8SN55iQprN14P+Ij1+0lz4AJZB+FW+01omRz6eLvdGK3ri1Guq/DTEIAmkKyi+dIpPDPolmJft
diPOwbhCoE+BiQSBrCkufsrhKdcxi7Y46gn5/iBf8iUOmO0fnnYj4RG59CEOAQEe19l60t3hF9FW
0WLFmRCmptHkQgqweZNmSDz4/7fkSHF9fv0ASAfEgWh0a9xL4wFZdxES2pGlbx3TkfKo2FWJNiLB
1wl4w0JHvVHT3eSYIDhR1PN3h0V0CbZZ8y8OkxVvEvm14aasfvHYk+BcmJfbIqTbzjuwCn1vK7Ry
R0Ds6EUiNsBgG15t2U/SHWnghajKznJJUvxHI5JGPrTu/MfmSgWVgY3Vy9w3nvmuENii4hFxBAV6
heu1Z2T7mAhzJEubGG40WhoFHI8BYGAO2lzAfvbhcjpTcdCJehdnReT+OslNfKtRH3dc/9Emqs98
+NUHFjLfkW6oXmqpio1Qw06gkJoa0PU/c8wPFEnwPCurIv5J0eSbbmkHSvJf1j1RFy/g3sDJsvDm
sDJaAmPSBPFXzxlaQzGj1aX954BZOusrZa32kF+DZVZIo36qlrZLK7zxZLgj2rYXxJn671yjh2XA
qIey+p+oEnVPdXRD20coAVLEyKEccGxNBY+8BTFxnRKeYaVCpSkD+j4NqbFuaGHuYMFfglhJBvk/
EJMHtuSVVFwzI+6kMHHvZsyLyHRJv2U9HNeagFTUf/IGXi23goiHeogC0Pn3BORH3c0qi6CdA08m
KINDzi7MvmMw6e0MvdbzL2dmNlvx5nC+/DxfKqyQhxMt8+/0q9KaZDCklsr1M/zOsTAizJzcBiD2
2nvS9TQeABMATZL7VoOFlw5gUcZzN9ACdlPUuT9jSIImKuJ11nprFlm7pVC2aaI/iB8072WIkqai
toQiRqb3cN0BWe6QfF/FKfOxZ9mTHBssYK7dPmPfFZxneoL4IOF+1J9Q+4Fv1vZBTUPq8EV8FxRq
Sj1zrDAMWZv70VOclrrs8WondoImcCFvsi+S4VDbLDOcouNbOHaCwR13Py/QnKZG9EiiVDnlFeRH
MyIeCvxt+ep776jnd57tnM3Rru/QQ6HpAmEWrT9vIJln3f/Z0Uhn/VSwdpSMDkXxBRnAeCVWicKG
3nM7YxCBve5Y7h3+D90QzT/PmNcHuQbC5sWbedok2dMLcduTwimtHwjq+LVGTRtqjpISYL0uhPhf
hk6hvi9X+ZoG96ffc9xHZ6oyXoFIJ6Zw/380+UYVDgosxDdfMH/ReJ90asbkOPqqzlG5rOZP8c2e
F5X+UKGYDAsfRaPeTDKe1dZCzHhF0m47K7vSI/Zd84TkOHOxutmfHezRF9tzjmjk8iqawZmq4NVu
GZuRPBCURtq6VHjr8V2pVv3RPGCnyFRgtO5jB1agiXDSpsEqTStlqizE+zbOisAwjvtNVzC0XPki
TRbb8inT21Tdq3FaEnD99ejzkv6dBfCOjGHsTs2f4VPS5I+/OdKqoKwpVmS9jHkspv1hEzCHfG/H
3uA9KosXxlXOwSZamSvdHPA9QmmtTUaq7jzbP7O+N59sJ9DfMA1Rd2xOnu2eIuhSpZqZDVBnIraY
0plIXylwmuhXBnfDJNLEcyD5NEeysExluztmBanHhMLJdAAALZHH9t3lBuSPIyaWShvNNbuioDMo
yqcl+l5Bk1ek85JDNF9dwSp1GsnTw+nXJ22HTwlD1FLfV7/z/4zLj4cKN+Teu5FFsU7FlFj4sBT/
F1wxZrLCM//RW3mFOsNFGj0bJVrR4Q6woDjS/Vekk617TYfBC/yHTq0U5B/avX+XVtJ9wwlHFJFp
JZJjXu9aH+Y7k+mB1fdfHzYzMV4ZFdlEOmWUBZ/cCnoVq3yx51Ey4YbFT4eaCGiTD0qJ3K5n8ZyK
7evGz1UuzALaFR7gdU+ovlkGJ4gBntxx0mp1xJjore5gH7jPz/Ycef4E8myO1Afvp1o5ur2E9ETl
BIT3O0Ye9v1CY/+phPLdzVuSIUo6bO/9NUs9j+B/KWovrtzCdnYawBmRDpze1y9Ujb037blvHXsq
yQca2eYzqg2Ll05fDALxQzDpV196PpT20WN4p4r5VNMJOQwrqjlk+AptPqgM4HOY8RxT+k7pdi8G
2szZFtPX8YQ1UDXzdONgEoWZ/Mj5QNYW3dFrnuSKiDkqqN4p5YEc+KtVIE+q2sWGa7ToGx1uTLEF
hFGj/3o7AwlIdHJQ79ivu/zD0D8Lv/dftAGmOZCEIapBi+wiWmPPHnnuN/4WklOdeOvDH2ANHHs4
bSNXRC+J3vSAXi8WcGvAbUC/RyJeG7kPzGooBArcb1T+6LGzBeLa+knrtQRI/l1cnP3yGP3CoTl1
Co8gSBOiAKRZ6ZO+Cuwx/Yiy0XxPHHTMNcpxGmoGs4TSrVBS42L0KDq8gNKUt7BCScDyw8iYQQWH
hQCRmoje2I2+CEWWb1JibTxwKVzVghzn/idOx4QETkf5mvapxrw1p8NDuxkUPapqs+AmNpyFKcWQ
YL8XYQTvKwEvo5hSwrNGiIGAPT6asSQF46l0b579IIjleodyoQJCGaagXA+O5Xu4q8H/IwxtJQYu
BvtSgXdfkzfruz9kH3vKpxnqcmn4W8aJ9ETw+dA0tXopRy3GQEILdAlclZu8yi0S8xHqCHJiEUC9
ADy5ARcj3dGLDSh0V9HWWcZAbQEMbr5sGRFSVAcfqaeOgF+dipSlewx937zblQnC9CNIVqvCFsEt
8ssF3W3UyRjFfkI0AbgomFzWD5mGfl6jkxQZiFSaxZj8nXOHZQ7QlWN2LLv92dNsJhBZTkz4ILyN
Dy8NVHpcNT1nr1gBm7yO1V8cmopvCq9LWWFPftgx2mDaOHVPdurUHLVPuwA+dhoRqgkDkFavIIU7
1DpGeWzKRkDc9H4TdkyqxjwNGbZjrXQl9l9F9xqFGGV5TqtFAVwZo3WGtVPE6hXElUNa+95s8wiD
e9f+LS9l6HFP/IiEGdf0mFnPSf+zdnoHFWTWwcCmgnUTMUmmE2ua6yfFvbtpAHXq3IMlwhjgLm+X
Iw51G7ND8++PkO09+GbpFhhuW3CGGxdOmihLujqEgllmvG0WqCQxOXVU1fRi1Chdle9Bc2CLR1ja
iJxucocue1gXl3iSiAVPvnMvLmyjd+odA12pLmA2Ddk5h1Ccl6nLLh0Nek3zwKQqo75AeSfMQjSv
yIU2q9Ap6xa5HacSHzdhN+hyEuqmVQ8z2VhWEOv3+70lgOSD6kgu4M2f1ZeAI4qZFByUODVdQz/2
WHy4ApLJxUrnm7JIbDbYHrVGomvGiegZKe8NjiLNb/sRgG5yNAwoECoXIqP9S2CjCfaXIMDLlXZi
1TGQsNqQxcvoHgcL4URK49grIUOPZIt4g7nR7VUehOGoCL3rCLuhabTqOVBlBqRoA8EcMiDLKYIz
VRFvTZhDFA9rEJQbPlH/o7PMte+7TEcZKsvXhCPWhWU5A3oNuIBs2WL4YCcLxiDfCjDeHkn2jm8v
9cVKhYlu/ptJaawT8n759qBiDWHcPhF/reJS6scxJDbBfdAUTnvUkDO3nQTEIrUkQLvKiXqkaWPT
d9nhyE+n1eADofKtHnEuXBd9/oj5lr6SuBXlpCmjD2DuBEaHxxXtQox2J46hmTAv2CCwo7gsi8V0
te9mY9lbuP1hRcQ+VOCx2e3ueeWAK9zTu3DqxhsMjg8ppT3ZesNLiHsXk/BRknrLamiVhLl3Wms6
ixT3wpuS36HZZL2INDngwnF/piifDnXVoem1wf7RLCRUNWJjNrc72GDu0Rrph7R1aLSRVJoFwac3
SL9N9q70lj2VVASFnxMcQFlYrq0o1HlLX7LcHiB0BSES0Uk2ErqpGqHIPzgPnV7uVkziNr/niENP
Qy7VZhr0514pdjDtZnSzBJN7U0w0mMmaaB5JQynXNMYii6Yc1cHvmx8giN3BX8UXdkHN07oNifAF
nYmgCxGian0DbUZfUI0LupRu80VOSng/XgL1nN9VM/VcBmK6TkqXVZu0m5Ua326QRsPS3FC3nqOU
Qcfg9kjPhfqTbMQy5s0Wg2xAMd+FuKfcOydv44lSRHKBf9oWs4xhWPBArDYykhuVunEEHSam0R3C
uSvQm+DL/wwZsY1gLW8NNL9shrKx68M0VCqJ0BL4eVf7SIQ+EalV8mIKldxHpYXzCimuIESJ0mKL
ISTK+zgNNsk+hdozFhW11lzMYabCQ1wDPw8VPFLqphhmcjynrSOU0bM4T5Uu7vhs0Yh/4fBk3mLc
zr75XggtZIoghM0MRTvyp6K8ekgbrV+ZZwO1dBCFaWf/GxKalR05Ng7uQ9E/6kJACiQT8Mk2iEy8
IrLEmgyC6NR9woXa8XsWis12vvbWA1UcaD0djVlsKaSICsxhx4kqZkXQF5hzD8Szms2Fo2YidSkK
OhDgclJLFNWqqehrjDK7BCcqp1sqqQ2rOhMk8FeXe1UbG9jHJa8qEMloTHC6rcBf2RzR65m6kMPA
cgcJZCVunu2tqzq4NrgTxdzX9w84+m4xEznHQ/jbT3gs2mGeOMtls4f/3MSnNIv90JuMZTgdrZVL
uN9yQrfcKXmLkBbiYtQB4Dcg1AC5NTKErudR4j3IihRKGtbrhCBIP6BgQfB7exl96fl/cptaM2Y7
DhB0qpyl+aPdR3B5JMxxoV4Xc1P4t94gG26/yF8ir534j6Df1K7WWCmZdQr/kUrArOyrBMy/H3AC
gN/hHuCT63EhqYvWPrZdzcI4m6vR0rrC3ilEZ0dUio22m5wkMthr+EqZo3mG/tO/HZe3MZs1q8Jl
VZYT6xeU7oU/yEGaUPO+0Aui+b70yPZACFXia1t+6j/KlAJgtIhPo3T9pY0xc1k6KlmstjotpsnE
wb93vYbBLr1DZgdRJRn7U4mk/mNB22tE5IG+JZx14o57deEuy7awEJRtjWg0MAJ0z+5QEQDRY82z
88JJ37wm7+sKWc6Rdj+7pQYi50SiiWz+C30Fr0i6hAxHkp6HIOJ+7y/yGdoQ61znENcFv+yAUl2X
sVQbhiXrNF90tCKTc/Az/y8R/oNj85wHwVmrDOtECeIVZ0aLP+J4J6bJc8SrP7EbMAU3mf6+w9+j
dYpb5hQQgOXJDmxd1mgSE7fBKmC+KusnH2MpsZMjHG9LdDVoozkxvIJ+YtxnJ2tfPijcmiV1nCNb
sJ0W3hLGpiYSEYA5LCXfDgB2J17C4kRorY9WfFudyfuOKSUrih+uSAIXAwd+lAk7ldBWbfDilOBb
9dYpiR832Idm3goDOq8b8iu82icLduYcjiQ9/hd6fnXet5WkLUQQDSwQRD3GnuY/bWlpc3gFITLF
OhyR1Qcc6RsBDxVBWUdFLLFqd1GjcOSjhseXskGroOh+9cktk+KYS0audsTSB4fvS4tr/q8++EbU
x+23EgfE0HqLk72eH1BjfbE1qWkxc1LYAiF6m27U7/Pi5yShQc7lEM3J9+U7jSYX/OdtW83896Gx
jjWgNx7kfnJQU2K8uekIw0zyfHqg1lFz60MinPktmEQNECH2qQiJdOyoFYPg1rCDmMAv0KarpwXl
bfLf+k/dkkEHZmtkoa9HgGrMfDsq0jWHBYTGZVsrbRGFv96BzZbTxgyjoMQ2ShI8oYvlvB+PaUMk
BeN1WKG512Wo2LHamdldIgM1uqssIUB5ghvnU1RC67YecP9/4ANlWQCkrV1sZasB6+mvNN8MTxnq
zjocy1eWETMO7qEoY8mppNGYe/+sCBV9UGBZS0VIn5H4Mw5HLJYF/dREOS0boZYgo9ddy+f8IXmm
0Oz4et1w6VlAhGrIL90wMhye8y57ke09F2G1JjOTcT0M9gask2ImsxtBHf55NCMDlYbpG8VjghdJ
7DMnHFHtpLfgMkJOMqa3U0RDM8BidImtDYyypWZ3RZ4iJslez3n4LHw8opIoQkHNbeZy5bgwLQah
kUOjfZhtSGjOF5hxGFH437wj0p3UFcZnY471B8Qgtze7xgJ3LgpSttyVuVB9liBlfJP3l0EotZlx
XRObENeNuoqmMomrN+YAlJ4qB0LAyC56vClQVJxF9r2phXO1idnm6KBBUZwSVQ7DnJ424sti0Vxs
0wteLxUsY3IVd/2N9mtOPzLuEuNlAM6iMD0rMyJCFg5hvBxQsimfnsj+U/MJhuS80qDz0YyxtXJC
otjvvSj8tb4CEm7pSPsVw9Jz9Q9Z75ErSqxN/0mDK4A3g+zUsVaYdhvvKSkcUrIW0DLrcuNKEmrI
C52UCnXMfA1uHVmFkmil+zZE342cFpRNop+XhOgh6v9pJ112kZbVsV01Wt6G+R+NRjznrfVa+HeK
lghPx2YLBGqI5yZcbIdgOxv9/G+5qWgjS9Pcq2igf4hZD+f9iPqGgnjvjDY6tNig+Bec4uqLqFvE
9jOz/FYXwR1+8Y1/BRuVlMA7KIwiJ9nto6TU8joBil59QCqsDMgrfxNJfNpXYdhFenfg1h+xgzzx
4SOnD1JgOQ0Zm9jvysgUH6H40ASkxUF4Xea+CfCAn93EWX8a2sXxYnvc31WAkHhAi7Ec/b5xqsFC
rFs9m+c/IWURXxmxa643hZhhR59GhvLIWnp8plKWNdXN8pBA+VTMMsiqzwfs++XEfvjKblX31KaT
aFzxFt1rQa+bmTiU6yUY3ENP1RjWXYwoo2uyYuermGqCkfqkTWQUEtxdk3a4qLFyXSCWFgAuo2tD
/VHzJTDF2psVuxH/coBdlFnT/5SuQkWK8zHuEEJYRirHJDEvSy9+zXjfUrRxNG7+tiD+prambUoS
xnRDnUzUi5eFwq3cLHBdyQapJqonFk/5LypcQa/+WfeEW6NDsfvojWPNV9QRxn8vycaBAGNSIFZa
6/hJFTdaAYo+vy5I752h0Zs7KM01bwlpqH2VeWnzdV0zXlqhap1GTV1cZoegRxMD1VRycmHwynjU
BP4wdtswyPM2fkMzZD4LBQvWQ3kbsvIbohvC5AOoxpVJDRHLwUWSssHewDw2hqaNn0ZT4qVWNXTR
v1pKNyXnz6VcgOlFJPfO6XYdETVSgOiJ8cSXNQSAuzHZHiLiqpon5z+96SBvd2eLrDqQr846skjq
0WMBphGsHxJZ4b76jrHr21XqHXciOkyvItDuCtVkDe3Gydt0q2OQXywgTHAXqzjXhJ9Bai4Pvmq5
rRcfT2VRlfAwbVRBZXeEIKYkprf6Bl6ZOXdbxKWb8xgJfKqxqqTtU//PREusezNIpNb3PSnkoCRE
eZwuZpqxcPhiA7Gx93JFdG9YHrNSXiysoCQjh6YZfL6flaQSlA42y68TSKEYUMJYD1Ac00hua7CT
AKk0JGP8A6vBNdUKZP0SouDTWCDem3T1G0plmhRhrYbvC1wThBSVsm+eXaD3vhGGKWLhWmMPVeiM
0prDuMB+eFT1KWAzt8F00awl2obw2GpvgN2YXgghu7GR8qqKOMKXnNCqYMXPwyWNBYSAwNEbRGIQ
XKaGtkWVZCgz2AhUFzkrc+7otmRKOSBMnn3zWBAyvrIU0GcUBINO9WM/lO6rOse4fQtaqZykkVzk
ASBxLpqTwHv18/EL/JFobkR+b0LXwyIxwHm/YEALUZzcabw5mFYXGixYNLTwzCJLzMrHLzmeRXPk
ysb5+a7zxhMaOTFxdGKWmj6F8vMb2ybSxglQcQu/xoD0OKOF5f/A8rhEjfiL7PDzhkL5p9aW6rdw
g00ynEJps5Y3NJKFru/pIs0WtYgvCrV6xkTWam6erDAHnARKj1le22Ayhk4NmBcmBv3ocDjU94iv
8zh/HXgS+mgoL/fgBuKV3XBJlHUXblcwVgt5ua1aCDUXYMG27Dqx3SOeTGWKe/Ws1ONFCfX4xw+L
I0jVKwrMhgReHo2s6UDYHtSOqTpShQgqVVFvdoCRVEOYT83kqIHpQojTbZYLY++IbWDcFifgeXYj
cYMdYwbw5+2/0dZ4OdYs4vOF/JHygG+nN9gqdXZAKaugiKYa8/awJrADfrKNezXzlNQ2s4TysmMI
RaBsQk7tC9uHJg3rOCnUYwz2cA/nV0Vz+ZYAxotZhFwGWQXOa1LXVwsslrgibPlKMm2WjhE5iq4A
KTnVncR71zjV5wqQclzN/Q/TDFQwJDbihrE1PHVVltjiAPTacP76vn1f8n1k/o+b1eoYb9RA5mbN
H60HmqjWpSm0S3yaI6uFzqNHVwnU+/Qdtck+KMA5vwDZJiTYmO5IZsd0pQIg9iUS83tKBmzj7eTb
noa+mhNyup9X5dEKDBsBPnSLe0MYLBKoFaPSJ1bHqHWMQL3OGvYWKqxJzAl8eGFJzCG7dRZjEYoa
zfsIwg2rTzDWHzDUH8myPPZQI665ykffqcEzKoGrqTrrt5AmsieylweW+b9QTkKYEGeRXy2jUYOq
SEDXJEyGWM9/kU3Eh++5Q5Kt2g/h0EmEzzPxA98Im1Pz9w5MKyGsqZXAZr9p5OsHrZLJlIbKMx/d
r72TMWmv25tsJdVAZfIsTiJJX9YEB1j/m732voS2Pl+VRtkJXMMWF2RAYjV8q8Nyig3beqz3x1Re
lv9Dmk9uX+fsk076L9iUyif7p05/cQTz9Bqu2j3FGRG80V73zxEgf06NCucaIXl+wpnyW8QJkYXD
V1Bp0g2bnjqyR3pFpwCaakPLbpw88CzRH3huDAHxP/dPXEcMeNY2eiiin+VRtlKjGcoBmEOKzIHC
dKt2sjKjCKKIIiFGtsCqllHtZd8lmRi5o+axddAHWP67W1XAHkl/80RT/1GgPg8MaNEP7A6LA0sP
vdPfKBTCLbeqHL2ZeusKQLXIsdBEps6mboN7TeZEROy58z8tzLDNgNVJaAUWzDx3xdJwJ2tFbrJ1
9NbkIQ58MCwWu/+01bSUJumTLrhPFM8ywiTZdDJwCMZ/Ryn1eLHRuDSiTkovUeKWRk30ut1rbAud
uLG4GmEfgvnY3nUqMgcqK4zAaYD2ALFSw3IzQRbsnQ2i8ngFRZsDD/wTcn2lTBW6tBvCxgxVfKDM
BYMI9PQrcCovIyWE8GVUrRs0GGdxHJg6ASp4J7XhbZvclgvnsgGSzWn2+2piFT5bpgwV/DKnvhj0
gWw1t52k3paMKMcNcprBdgSDq6PJ189orobX5QmR/F+8rjI2ePNSFaxp36OWXbGDOZyR4w9AffGj
Z5KUgxs/qWP5E9Fjnv3J7PZpiA7cPqwOLIJb7oZfvrAGLUc20ZRv8Uc/rq/MO1OWK8rDkhgJB1Ar
Yn5VdofLncOY8P0xuEnX1enJohK7lQX/SfpD+FOKIWi41dW6ZQ5uPCi9K+IKBkKoJKlf1XZcjA2L
38SSsUe3oVYhzUUNHNmr8Bsc+SYbPfj8zTCj4lzDjf1/yywXmG64MUsDrV/EWmBeRoQK6u98AM2I
0w6xyo7HouxEF0Gaf4zEt66u95tlAulSFC9qakVhwmvCX/UHMos0Wn6e7/AmfeuCT2jGSzoVD0qh
45euYLGtKcGw26I9GDjwVy76tShz5KYcdWVBp4g6xRKpk6pbBblO/wlCeG/IEWC1j++6oYHahVxY
ce1rAGo4gYjJA4QHa5QXZQGCCZ+SZAAo6NlP6TU0jS9bS2tZokl7NATQnpPM/3S8ixlxVyzs3XiT
ZOLMyIHEdXRyb+VEzLTmRk6S5PPPZ4XJpoKFHYV1Hy20B8pTsvk3GpFuIUccJPJV1qwmCgaYZRfu
gerKRyMw50LCO31JMocFPwjeBJKgCQYFhTJzSKK54Xvuo9xObKXdIs3XLP9bG54nG9HgdfonrLJ7
73Ed/a6zDNGHotI77x4cMwyZEV8StfharFuAmpXMZlz5d0MkjGZpR9KVUgmavd/mmQnC1qr8PJYT
AuxqNbD+PawUE8MhpUeBVbw9QIWTgmFmM6gZDSHRcqH4KerpdpnNS8rDa+hbgmdRxEZ+YwCgqWaK
erxy0BcxU7KLXc4h7ze8X7yt7UBTqW6rwYBLQKoRWk12nduu9lu1PT5alWPmrKfMjzgos+9jD/D6
emywrAuEy+Keik/cm6h4izGsaUH9S6t0MKCotIYLXMhNpYfuURomvKlrGbF4nMblZCmpxloxE6ut
vPG//qxGcpUsCo/0jwuF4qjx02ixmV1Myq45M7PrbPnen/Jd+iad5bLjPLXkL8cA3FC6+7kV7fVb
aVWegDrhsUox9oqMNgmAP+IMsyFm4PIUm9BGDpXckcpOT3WBzIZZHuNhkCYQwdY8tGEuUeJQxlzp
Yht8x3u/LEs3ZMxE1Mk13S/7FSlyEWGw16hAkXiLq7uA/pJCopSokyMLfML/1dlQXcGHjE3VQf9N
Ez9zxNwDHCayiR/74ATlMTK+jryJrQ+rcs7IGAa7kfwKjLtvrcgs+j1sPkUn+tiPutp7VKmhVjlf
JqMrRBQ/8uBqtVFniox9ez1kPMSwnU2LHEjpYKLL6JPHhJpVRMdzoCy2GSkZFYLPEI0UhuySGlh0
yP3s5TbVJYewOLVilWpsAFiH6aPLllULz4ngERyrMRQvP8nEHclJ1VEc05YvCDDphxgzuX1C1Pll
JXcorzyFR5VZG+9w3ERosNf5RwPdvAx6ECsJgpAfF1v0bF1uLbtJkK0DpylkngIjoSAvxsHePWU2
PYGGtwj2p5H4DyHI/m6vNwl6rhr9UXOVugjEGSrlhKCul2bLaJZpLE32qQdAoy2okVtAJDkWtTVS
hAOUdxdBaj0YdtSYjQ8jd6K8OAzlrwV6PGUSsejLiBoN+l6dUxveMI+u8QCgWR8j4GvQVzOw4K0C
oo9Xd5L1b+4V6l6g2Bb/Mm1s8fwEZ//5eZ1mgIBG5J9AKUzi/cSMEj1AECpDtbeP1Z+O6xTgONkv
au0cLgApKJqegOd4rIc+1L+mnXatjuZnUGce35yGG08IJGTT2pvt6GpO28CMiXIUXrehUZE4MWut
lEY4wBFB16xlti2nQBzJjgvjliWtgzyeuAq1mwV0w8mJQJaM47p9oW6j693C5ncBpm1v41nW1pCX
bx26kCpefDpgaDne9R/EBNSxEbEgOk2nGYQbRr7STXkkytkHnC1CoK1/8CD8OuVHCxBgh2nQQPZ4
cx84O8PTXdRtcioHAvwDxOYaGbyKIA1KzDOqs9KJYcl8zJHUVxpeyFr3zTvMXCu5OreGzNYmlFU1
+kv2YBB2ZDJaEX2rp3Eu9JLK41dhUI4tnR33O/q6T9EZJzLJpvN/2Zt8HQbKTkVpQsrOxPUKnPRz
Liuo1vTIuFvxAcg1Ul5LcHLzzP1Hz0xL8FowUx1kusRxJKqmwbrAHS7hbs7ZxZKBze1sxLnSXTgF
qr6LqDewc7RyyYG93d5+4wlzqJjMN22wymh2q04eEyLyJ4yNA5Gedc9hojHuJuYabw7Vv/URhgWn
Yyd5vHJQVURZnuQOcucdM4tT/M+bWzIktNILKfUO1zvznakFzQyqf9iuL5yaqBQ297mni+ABRJRM
p7a3dQnw2RRkx/fQkzYiGnR9HooMMF2Phky0dTIPHi4rk6I3/MS9etIiGJiPA95jAAx/3PEH/PAz
oietxTvdqj+y2+sKObpV0mw2o/rFBwhukKxqEclJh+I+RSfBVzFnY8v3Z1KkwODZIritNF5uZu/m
3JzoObEB2IKJWM271eP9M1KSECOMV6TF+3Ln5fcD0nDs93iS02N+1MDgW6IP3LjOZrswxnDhHfTq
OmGZwYT/1sA3Hzu61yBpmJHGCdfUCcn9W+2YDVCuCbH269MlaYPzWHhx+GLieqfVuUP8Y2RNhdFM
5Kq4wPv62JWKcwO2+FHmf8kRNZTUjXHOBy/QczDtHIbMiBpglGGROleJHBV9L5vhhdHp+CZnJN2I
l2BDZqmdMQMaMhDfcQL7pV5GFBijhPjH5Bt6vw+4JwAm0mZgplPIVN19kfDn7C5LMneauJf9IV82
H2hijZQG+ASNmZ0e6yuGU8uDjJmaXjOIPf4lJihEQe7HvADhDqKM9wGstzkHKUaovqy3ty4lR/xg
0rN6kZrpxuffrFYgOF/7hFT7w/ZXNHyJc2MEhgm8uRgLvUZvQcpNhRtfiR+hJwa4Yc6NAPf1feTr
I3Y8ZOUyalaKHmrELvoLHBAl9fEfudkzvZYpf/I00mvnSUdAnXyYNvrbkrxwsjPHzVJlpHNhs0/d
4RAbyk9sTEm+gM8IabKG2Fcz0147mXnlvmeFWOqwHsRN4mIg/8sw8WoroAvhjjQqNfa4SwIVT0X7
q70Bvk/g+ffWZq5MqKacfiOwk/uT5tCtGZlrb49wf0aEzPMswagRgV1D1OlMexVbGsj4SU020RoC
IOv+WmQ05+uCYGTqCGGsFvC7GKgUBEDMzlKvRF6dZh0zVTeOb1xn8Zdyg6xorHONXI6yK3ZAZbed
uIjSm4VqjUFX1rIi/UlP8u9Bz4mBUCv9tqmNJfoewEYGVbm2iG5eqoZKTUr1dHnWur/b05rT6quz
TvXDAL2xxq5o1UoKT8zPMlka37YeMquUz9SJgLXjnMPpXf0CfQRFGGvyfmYXBeOFyl+2ng8NHf1K
duDEdAemu/GKefjQY4yOLlQ9tu2skNaFB3RPzzvN/z6e8ifBXyuNc96t5cfRylvTeoriMGydUA8y
8Css8DWxOlv/mp4f7PCJJRaEbSBkmnybr6V8N7nTscr2EcJAyextAa9SoWunRgoojvMF6eluDBxx
UbcYMJYof2FHWCK2iWLoj/RGRXSEwDMlFCGQxMUcBp+nMU2kvkmWugSNPO5eJKT564H+0Hz0gvzK
dNnWpQQO/upwrQ3HzicO7sEAZYWNoRuNjUUQArIQ76PrkpiHUg1EfSp3nSqOHomalDJcmXKorrAh
TvbEyX7FDfhfMhJvW9b4XPNmtl868i/nsLb6RGZCVUIj2uzxRvuIAjYdjMJpgfEvCx3epvnVKMut
sOxTWC0bHGFvc1FBFzsMZjoMbuSzLkfL8mFnc7b08Wpg40YL+h3qTTgv0yUxa38hTxqTSPxhF5Si
/bvzE3wH6oL9/moDAjpn2hDxlAzm+ZiqK9vsU7CRW9CSeatKFnJS09cOuR29OrKu78DlmJpFVlNS
xt313GY8iBW17hBz9SR9S2r5OPlP8YP75WZThb5zO5K/jW7gWub1yDfdnK77ioDnc9TRAS6MEYP0
bXsfDtZjiAlUVI4ZdwMjOh72pTWVv7Idj9zywahUBkqCIgAZFQaPkKUTUWYqptYachc+yHBWuxVb
+gpDnCzgtu7BX1lNqj5jSbVGI2FtuXS6fBwOHNBby2elqxpFbmFBEko6aqfaTcpw9DzPnBL5ZEmF
cPe5Ztp8y5czX64lhu9a/DSX2DaGfRwACn5ACMDK6KCKVcx09xnTI2aWP8Gtrj2EB7ACQF1MuHyJ
+oGzIzxzn2S30rGkbeUTzf0beu78sj/hbpgzuGQfwNSN+1wrNnjRBFZStxBYUMNKGYjP60hk3dIp
GAIZ4vDSSV3WC8UHTsV0O9LHjgtRQmxJtmWyIGB7FJE49r9ZNUpfTzb4JAp5l8pUXDhV2GbHNMYf
s1thuoww6jgLM4xkL6mdNEHBrogV3ooyggj4vjpIj1JMw+s5JifXn1EqiFTBrkCyjbrKeDAs+0+O
Ub9ygSr71eODNbY6Xp6CYHJwbKFDXneyt9z68Yvcwy2TonYC/4qgDvJ8VGGs2Sqof7Sc4nF8BoyW
V5HSIBIsTcfMB79aWhSEk01nCoxFKh4FUtcSjCg0gdNcvopXi1/aXgm6re5F2evTkasjg1Ap9zkK
bk6arW33wyYVLEKR/ZfqeBewpUyNw8bgni2j41tRt2sfKSJ+0SCjDSZgF/5RcS4vUbt0yJDIr4MJ
rcRVRG1ocbdQnsnzhSwi4IbkSihlsQdezjlu2/KpqB2sQu1sSBp7OXRCXWpHzRAx307jGRU0pDFK
FNjzKGa73RkIeiEZx6yU+Ufh8qBGTbx4QbJBh/UDyaTxwkQuhn3YfjZE0G4hhoM9k0D6VfJcHYqO
MG6zQ38MUvM4+t8Kyiy8EJOQucDKJaSwbMKoyOtB27pbb+cnPK8ixcXHzrN7Z+rHOLOsqe1TCzAt
JD5i5sSKlipzXaZAWmewlpb7pB4zSPTpSAYN1PYL/nqjVCYwSr4PUWBIVMNSNvOBBBrARfmUlHKr
Cw8EoJbLMRhKYsPxgPGHjxAkIHlChe9co+4Q6xN4Z8zpwpi6XZQLX8ZckJFCzXEL7tGtwIJtxUnM
Ftjs/YLKfyLdWRqr455zR2wkQPYkr8R/D0i9riJuEf2OfkS/iVG3QJ5/tmf4PSDDgDz+Ll9RGu7A
X16pilBN79byTP1lpEyUbCE0z4M2GuiLEj/UVKab9NnvsXkWIjcJE9LmhHvOR9RKDS/jfwgDMfjq
XcVoF1n1tw6grwnW1TKb8Kk/zk2bl/mESSDNAW370x/aF5gKTNxe+kb0Vq4Txg0v/T0nNjXUAg50
sHX4Wo1bY9C5ILHttQGOSvdYOA4NlW25TrOQeTXfx1ZzvzCPuZo/sZs9n5cKw9A2NbS5xIFSaJ4B
fiO58aaxfuf2QuA7SHJQkOu3KSZYQL3nmNKs43XVYOE2h+XUeKYwTQo9GUgW5HvKyZR/R9paLEhs
FbMDdI6eN05SSKxN5J6B7LY3PTdG3i8qEBdZv4jfTQGHIZd1Pd7092AsG3V1vs4PwJuZbpFv5ciN
cDaUJxqDr4FTbmFaSeQHfCQVsYr+TGC4H9KiZ+3ctzSvzYWnLVqc02hmx//XbAynoydgF4xqvs59
+/OaweKFOZJEflMK2pBeXTT1b6DaGjmvVvmkM71Gh0VY8pXN3M4z8fwJF+NyGof2qyN7Z/eVllRK
odfK1nhL9aTq5gyRDUtYcBo4Cm0WuUciqlaCAEJ8StJ9KdnXZJna9usGdLGZ80TrAkzfz5H13xtH
CIzCKDnDaEEYR4DFBcnbqYNEjI+9r66I9pcKmZrMMdP6OF0tA7RyodfSEOXjz6ZEiTZlRXChT4iT
0nOn4jyUnZEk1hDyW+5ysdMcLYNdv7q0PIK9BvGbmUP1gzXfatj5IUXKimIpL/mPY42ijWBKHrQB
9H+Zm59CBD1mtfXEbK0arV6E3oPnpS3/z58sSwKzmVtZ7JIfHg2hqNAflVX6m3/OYY7vLKt1gvDx
OQePYDZIZs93RZRkORSof4ZYLTRovhYuzIqfiCGtApm4RP1x+JCW36k8FaUYavQLAdU13i5tGNqo
ziLWX7xk8UrI0f7r6JGKcyBsFaUfnfOdQo8le2IYnI6xcmDyXMttoS3aVSt9AYaVoO8Ckvwz+3PA
FnFe6rwme5W2fOGw83ZkbTUEs5zZZeti6pw8Ri3T+dfvcDTXdPZolB9oBSj7qFbUZ01TWKEEP4Vk
Uy4icUZe96VqkMMpcGJkScxJhecDkR8lDI+ZNt+C6784ophgD1+qrlfgwhoZJ6LCGGOBL6ZKDqI/
TRHt84PNzK/BJhZApBvyb8QCUbv47eTI6F6dx334Ro2V6HTopyDYOaI0AcFnVl8x6Hd0CjSvWbLq
l4NpwBw0TaQDhsYDXW+nyjD1neDoX2ZShzjQLV6F2PcurAeAk/s1ZEOSTzzt/6dwifSfLvcBerWm
HE2GKVvW6yhOYxCNBuG0tOweqGRJr9VS716Y4iDA1V0ltfkpUDX8R35yz9NH/nnEwXKUn50nehn7
ittGPgyYTwfmeu6bFtS6dqBvIA3sI70WjH3S6RgN+mr5dKTDUrSnO+j5Dy3qGFzot3qOulho2GOs
05j+NSxvAndAxDSdUyCO4DUjrRyqNG/ZIsE6fX4pg6CDP4z+6rLdVEix0HIv3BPom2oxMjpngzak
EVr247GY1jnllKM7/z9EbbMGUk1nV/G8GPBZ7U8ddqOC8rPvrgCtsEquDCB7g415lvzL6Wyf24LC
VVuRsyMZW5N1tZnGrdU1DAlvOigAOOFU/9qfKwUsf24mNIxw10q2B94Il6+MLJvAEpwKEmrLDMgF
5zB2XWMB6ohVqp6kmrdfUUluwG6CJz7nK3jzS2QhWwqCKZe16z1qs1J18uFDNHCI1L8od/4yTGGk
RHsTL8tIzHrwuSLk1h6N/OFexdKTNWRR+HaD1q3PU+uqu2nel4OXO+xgl+uXNeD+biPhq6HZOJUD
Ii+n/GqfXha5i5gBgn0kahgGmadxv+3AgY5WsV7F5WNCu6x4Tnw72cEcBqgrDRU/U7y/Q0wASyNI
e9TzQNAboOZpNukD7OJW41lrECT9LvK+6LQmvjycJw2VZFxMf5uII4skSCsJklHjbPUa2SQ2nBDj
Jb87brlbjRv20L1Fj+tfZP+1xxbRaNCPYUii3ykWIy0FXnsrkoiPh7LpyTWz+S5Iz/Dm9sHMY57M
7ARpcCobW/Vz3i5fd9yRjpM/0vi6AxVmhh/mKz+gi3wytO7iUjfrt5KtTccDMOUQnd3Bii5ej4PD
gmdhEdb+psc15odZR9HWlEDczUYoWk2xCDcm5GlEgnDMHwHbWb+XvBQmuM7zCNT6AsZzrMHPqgbj
nen5H6iIQ4Xfd+7y6jn0bYo41XlzB+Thgi9c7W/GxNI4ELmZY5NlDIGxbYYLxloOh+St1jkf3Q9f
/6fW5YLxLxNLLAG8/It2ayQk7JCx4KGXa3kLUm0S9AWW6+VGgctO5voFRNRv/Ku52Gua/uvqceuG
8fx2GpCGASDxGjAt8pJ/payB4RujvHoFCTfn901p2jVrHToFydnJnSSBJuJXK5hKNho6vxUPnzVP
qIwS1V8ATABLvofUU5QPKfPOD68zjloCV2AUVNgkO49L5QYgUX6lra00Nq15z/0z9kI3tg5B5aSP
NsdbD7Sxm2ETvsyGNF8bj4pQGGzir8ME2wFVq8TsbifBtNn34REjiP7uiIScakv9VhbKMwB2pCsq
ZkQ98bY/Sk/oKz+gNuYlguoZT7gLJgjDuZA6niRnz9ff6ucreGCgZE6E7otwhJYcHJ8Y4xpqGxEX
4E+6hdnf5NGmKuOAwRxHe8XXlNIGPaoPTZ4gmRTZdOcqnIhwVHh0kZnGVPCteQ502WUtZTdclBJd
dpe5YTd1Y6Dt8m+W/rxc/wV84EITSJ5xAiy8RjX/o7aQE/v25FiYU6dU51sFglZXKA6jmv4gVcbx
zrK6uKyehApPEoUklnPOeaBr3RrH5ZDm+9BwTu2T7JijXONiWckrA6x2vve1njunQSo8wPPyRQzF
j9bEmq7WTh6phs+22UcbiMhEZMXfkMW3UYRkmsZpE47aJxvocPKKuqNw0sIxBVsKJkUKyjMPZArC
H/W4BSk+jcxo/Plu/08+CV9JqdP7dhL9aqSywOo0EGSDxPNZJffzFKm8QU2GWJbyz0+gXc3+y8aX
WrCSQr48+I+FUfrEpgEO6ID1ShnQSLTuc7StwMUo5Ye9Q66DmgQ41s6YGMAZFyZHdJX2aYmmatlb
1ieRpmzn6NdLvQ/l29uifAiMlfpgKDnoohwfSB7nHW6ZrslYyBO6hz5kn/cU0pEBOo+PNxO9jfMP
l4vsp0e/kk4uTMryswcFU42l7hS7+mwll4Y2VYl3G1TIMq9LlU2rVq7K4gx6jkuqhzN8YwdqUzts
awgwGo8ZnEntJMoMUI5qwVpLWilvFa5zz1hHxIVFopWZuNGWmD2G9vAkFfb2GpgRlJXSNl+VVfQt
2Pm3h5HnYRRrBiWwDc876Xvu1S+J+UQnt7d6Vxp3CBsoYEd92QLOharqpCvTlPC3cU+enz50YNeq
12RQA1ZVYtiw+k2fT5i0bDniWXP14j2WoW6r5J3Pie+EE753W18c15XFRzq3Hd1rWIrZtySvz/p/
Aa5IKanYfidZVkUqwSoi8yF6SrRt+FusSGWpUMfSVcgdePJeMgXMOgOFXP+GauuhKwmGZMHkt0+d
b+2Z1+xZSCanXUgJVkrSp4FQWExDFP1goRsHXC6/vPXS5ISjYyLWIIHlY/8Vp9O2CmI5nkdo25yB
0TYMloMAZxHx21Sr/CJVvcg9c+9IUiJcMRVp/OPn3Bg9kWJTGqvW2w+gJCWItLGjCDnGlWRItYb3
LTTPAW1OPR9o/Whb8HiZADahBMJQ9LhuineBDttwVYKuV0BdNjAqkw06DlwNqKDYVle4ZSQIDL9N
WBjF+Bq1jBQXQ2KkeGp+OHzGvNt+XtFmVMvQDLMDIRTdvmtfm8golpusqozwrWWypCgaXhn5wS3J
x93xx2R0UMU+CSsuIx873sGRKU1wNBjNwGjSZfTdI0iL4jOk2n7JisBzreCOXSOmH2qxwKUOfKME
t4EQa3t81Y9pNb1zYUQqdkJ54sqgKIQ+BnpQkzylcHkVssMF3zPMdhI9DU0hNqO0Q2pCUucJRTlM
zXx6AZYICBspjUbESxm3CTXIfRf+9+R0b7eC2SwKxyKmovidVphGCHnpIjfxT7DmJXCNLOU9/c4J
yGQk7QN+6cQh3/BOG77+ocBXSL4J+uOWD0VyXSoCDsY1hX7JLv1gm5+aG9bIxW7NPKas235IeRfs
eQn/bp3ma6t+movycZDmUwmmbWIP9RqG4XBLyK6K9III8M3UAwZFTARMiD/BNqQDXQj7fEMKcZPg
JEO7iNIaZD59rweRtTnk7StM1EbpytugMSaRouP/lckhHxt1POEzD4De4dQc6mbURUsCzxddQd1C
XVEMG1QGmQUNQi3FVmzVfwMJGxjyhpzBtvIbXkdy6tZaDxKU4VuQIzS48D7TCbqDiBCDIJLSiGFL
3M6bDW0Ks7awu7nwiggQd4qGtmsb3BxjMFNBMvtbocV+akvh1NehIU/KDGDAV8Gb+wWbgui/yguq
AN/WI7CCYi7RupRA0TrR7zldYi0KnLaGSDtCZH/xpoJ7ruZq/9ETmgKlSq4fNdJYEBfayeZFCbbN
EfAVdvsY80a8m1qEcdP/AszK840rOnbDz7LSKt2+s2huq547yqQvNZqVb5WNjTT5t0gMdAHgohpZ
KAegHJA/Hb8tlFilEz78ett7jI72uqgY+8HwDy0nV+S47DUeUDfYYVkxckuAxc/kZDWReW8dVsbH
UqZ0F5G0gjuQRUJN/BOKw3K3drGom/xaIfEFzpvDfTmZtmi6rEtnjmtkZEz/XIxxxONvkqwTT3Nq
/WabQczKDns33wEtIi8EJtXVvcyiH5dCoMarhaL47DecrPZZ1cpYg/0fNXujhlprQzjtJeq4K9Pf
xAFrw6PQqb8AWkwVUfd003k2qi0r8iU8KNCk56hjkTz5mA6hbBT8EmI61Ss07S0LJ4Yx3PC/Txto
723xFEN5rRatXF4ciIeFV7Dpx+uqNw619eltijwkDugAfZEuVxqee1gd08KoClazQyaRR+LoDxbi
HQo4L/i9bP2DqiJXZzjPM6Sz+GdeFvBqugZvRgVO3m+Fq8sbbRXlIqrOYO/W6eKwTcCT9vaoXd1Y
n72hgCxvr85JHO7cW7JqL8Ez4POD3z0RQ/+vC+F5X7jcXEfkkpiRhtHlafkYJmSVGRIyYkz3CEuq
psR/qCrD9wwlKC9T6FoRigRKes7td5uJ51sfCb9bMM72GBRRqJkPKEI8IqHrxbTobWbr5ZXF1gDt
ozzPls142HJTwLa5Z3+2eICXB9ArsiOJThlglyhU+sZtdPfMnYQX9scKz5Yhxp3ET7znUg8qU96C
TQDZFC/wY+cVl+8Z/dIC5Rpf6k+zJjQa1NXcFTC4WhBxGaQghJN+0fOMktZadX3jd0B8OZ3LV/CB
DiaVC96asHFlZfOL0Jf8w1C04T/d1xMDcGN5Dvi3syeAzOFADKsuAajshYNTtN2sJ0wUnLAUINxb
G3pgCi8O2lm1ZQ2cb0EN+emYMAn1V8aL3tP70hhaJvDw8JGK8kPk2LcD9eeOCF3gJfKE5+MvMST+
caVuIZTlR/CC9ZWp9U/h/wERjhupYUcqsZVLDHcgd93iShrE6DdTq9fWAtW/50Q1iP8aYB3gopkQ
yn/RXyvBfMQRH88PeTsjGMbRAxthcFGI7Fs7Z4+Tk/XSzAAh7Ujz3N8dgBy5H06thKdGOjhiKuiS
ztI9+RbWUxsqBQVda7pA6JqTHli/g8QY7FDIvomEF8ht8DkyTDYJ2Od/epTrGnHIBGSvuuG4udgW
Z7pUKBO8ozTl63pMC21TxeoyttdfxY9P1VgOibAo33iuR3NZMr+NUItzXY/aKhLD8TUJohHE9P42
hF0VGoUiwKM1d0+z8KuyYhrKsXck9Gky/LPsMv+bz7gKk8zvjTngZ01ByOQBYJJVHvhEHblXaXw5
tRB+cMfl+6dBmlTmujJz/JJL0+kOvSzUsTd2Waz6bqcKH/Kg079RKSw18OBklQYigXDv2skvzWwQ
N6CG6kW2TwJohGpNGZH5JU4M+eHGHLq3U9TQVGaFt61Xdqnr/PUMrVg8PTW8DaM0nFaozPur5T+6
x8jS7kZZrwlbc3zaaiIXLFzKXT6aOyHrhfD26U23MkDAnW/mo/GishOghPhf8swKMaEUjEIbdhfw
N4LZmlGEeRde+VJveW7pyJ5g3xJLjyS/HhWFc2DcBTrSa+fz+7sxz1ZqRTZm7EdgOUQR7aIFZhHq
z2TRViuJlfbk5e5BbAwX8/TRwUC6Ps5GQbEctfNXZhtVMNk5uaevJ2jzqknjfLsH0y8T3a6p0qcK
VZalH9TZV7KeUl1VvLZlAriWgfiHszFizaus5gtGjRly5Hzjh/4g146IAs/Q1zTHsUksfc7r4sba
gOgzwgJeOuFQI4mtxvWObPTn8C3JFSPdW/pV9DmkSrHPMVBbLicohH1fdCiYXHFj56m1Xk134FBo
4AEmzQeUI4TxuB3YE37IAg+R3YK9oGLWUC2LbbuvXwtROnW02d0+3Wi5YO2ZNU9A4mq8+Q3gdfA3
Eq+V13kr3j0sYnT3IEow3jcG1zyKvLchPsJfBzdm5HEMBHTpaP8Z+dzZyKmF833RBED2zWBmxDJh
4I1nopPvjDUc/p0gcn4/vFYNiaEjD1XLUaBmqRZu35KzijGLajgCWtnS9xghlF+P3APBjDcpznYT
Wt+dCyyXsQ5fuTOFOhac314oOSidZr0mXxcN9q5ZATo56jNodUedmYZ55n9wRGe47mc8FyOocZbB
Prsti6Q/R2JUMz1qWYlR/gZY4TFxzguhbeDaeBt4QOoGb+axwFgPVqMmHflQ8s86Py7DbHEuj/XQ
X7hDytQepBfPdH+M61Wt1/NAr6mbYAPgji3b8r1+s6Wk4zxOjI3r/R7XAyxV3OJHgpwD+8pXQ78w
7napRoKLhwI0UAk5v/CfZNBmWBO3Kwjckx1t3WyH1pODsMcQEywBXKQEoNjco12jdeQc+ClTQehk
I5D/IrdaPMItpFmiA8nPuWHoV+RITSIo8vMv7/8u5oLjFimeb1yDzuTEh4e3EbToZnx70wqMp1nd
SwXKrhsy3sQ17L3VVgr87hFuJY5tm83gycJamALirR2bCEQ2rE3nKjs18On7xUGo7jPs8238UtLq
xOzYyJF32ewg01/H0EOCsLH6eMKWMn9Q9PgSaWPLxJYfgDagwDus9Iz32G7Lp8WZYKy+KQPfE/V4
TvaKAPtGV3MPsQ690Xto94JtzmNXpLdCAdNhslRwW6uKVPQPFtP4RaHLhQ3jO9tu2jDd4FGXyeoi
CGveC2WAl7i9nxWRGGD7QGCoZAR6sdf4wOhoR+HEiTRZ1r3ChjhKGVJyab27Yso8QcT9Vw+aFyJX
GzVf6S9AV1/co7PVMDj4ZC5hEsOa0tM81zfAzr5Qtd2ckzh7tJ3mnJ7J3kaeoulO5ELB+D0V6nhf
Zva+LFEHm7i4HTqDUaD6O6xLUMw82keTRZbfCupf/oyFHXEy1wrfIIARfgaP3LGw2riWN42Jkq3d
bEg4h7TcJBqAnlAODNOT1OGmO3L02janp/PYHlw9nW2HFFGyOTDBqUyfXmsNqQrp4u/R8O29Mzmj
jJaS8ATjGQzTeZO9pUX/wkLgP3uXEzUys4pAX2ri02SJDW4WCBJ06OkQVi4n5S1FG85TtKUAOdI0
tm4MGuvVARpDVdTlvAbf1kx+B/5efaNHDMs15EQjRRbvZ675F2fMS7V0SheGqKpupfNsUUaq6S9E
/2pYaEIv8BGfBiGiSzWFV2g02YJxObfSYjmb8CnUxWaGwFrEncnxiHdzQqQWeH+PYo2JB434MD4J
IGKCcLAbxqEKZq2sFUeuEB5/6qM27d4tm2vyg1OYf0/hPO9H7dRThTwisCTqzoYiwz5PCKTgWpzE
R/xg2+uxtmVffW1sAfoAByngsd8ZQvYBs7nkP5E4yLL3Oer953Eq8SGY6QizrZU6w83RLE6h9XYw
ovLF2Hf5dSKTa8GvCxDBwnbk8EzHU0bcdVjKtqGTJqmz+Madt6IKr2lsjThKiQ1Me7ryMRYYlCOb
eM25g6ceVSfkWIu8GtmbgcwLVf03oJN1JkJmxKwAAXxT7C8vn3+zyLtCbvarorurMriVBMxygOsN
P/BFF4P6NrVsdP04BnB9os/+QvAQ9xRw8PLXumRRdbb5qQlzfm8jL6y//ASELBiKK1nSN5Dljq32
0x9MKNhq8BVC7U/BGgclF3vKf6agn7zukGznM3Iq+wPv49xSL8x7k/UcwGBx9tF9Gwf/XazPwSWx
NNh1W37Iy7yQPIhokqetXTUn68MzHeUcaoxByBr8ZBg2fWjFFGkRO2GblrfFK0C9lQpbi3iAkk9q
MumZtCNaKuivlvpfclEgGWZWH78Tbbq9W47D+yIXSyXCrCN2v9+XUi9Z6KECxgIRshjPKHZvtKHe
zER8npaa5/LCJl7zZGEjMFEC7RvI1wLTk6gse9DdzyzLf5J7W5kpWp/hIX3Eu5/dkZUCbPSywfot
Xw1GMm1vveCYbrvqFx28MhX/hnWyVSirZC/q6NyI6BifCfkhlF6k/+S/aTpz66fbqe758YxHPucr
iU6QJQIJu3Ttpvp/KovM/cFZZEBOGCtBodZHrUCqxxS4xrKWRA9X4KqAl5cEFADPv/u+MGkh16Nq
vyanSg/pBnh7uyM0PxZZKgSl3sLYWl4RRAyj8LlwgaEKTSdzIEf9LLIlYN2NdN+9yZMi0JR9H+/p
3bmIC1l0vHcMVykx+bHbQmiZKzl8rKUd3t9qeeyhBWnyq6hRHO5QMgLwGQxuhlhR4RMBlSWZnVLZ
9rQaaDCnzOC9kdxGj2/6RGRu0QgOyE//A+o/wLd36UVGM+KxiyqQgyi6dAscJSyveA1wAuyuXAYx
ewv1095HuciDPC9Vzu8YpvIs1MO0W9FTIB5BfAiawLqMNDhdblyXUc3yhhqwccgfSW/Ks8oeRpbo
jSMKTeIyPoKg8tkFVcSF+1eNhiNBu3Xtxdo6Z788tEomLQczEOAFXTq804301SvDXiq8Gn5BCu+u
tjKZFvPtiY0ptnWZmWE9GIn8ZG3FdG+FyFNIQOp4CmQkKNrhWHmyQPn+5Hn0TTFsFVeaWMmsGPFg
9xg8GeHQgPKyAwjitQuqz0debHjrimDGCNFnz6T98Es++XmQmANPszRmKxSyf+qaq2tRgzB9pwOJ
YcOcVu5M5tkAxs1wqAck9KRRKjJfYCwAKkuRKt8AqgOCNpf9Ow2joeG5DXOaj+8r3EDpVazYml6K
ni012IjTd7j7GHr0R2wTDImmV9czlDghknGHGBVfHQKIC74VyswWp0GopaTglURVRRq7JoQf6aMh
AkMpM4A/sJch++YTG+ZPp57Al/tFQqAt+nvwu7Q85fFj2iMDkqNyINJxlCBORYalW21rEBvVsQye
D1MPb3go9djHcXCsrhS5E1q/LrYWwQJj+AoYKU9/IBImV1RiIAJXESnYkwFyRmseLrs4zd3BbIzk
HcTEdNAkLmrJctoDTVHbbv/KJoOVn3HkJJdwa9hIpjtCduZYSwvPk/eisewstCs1ZtwJv9lYE0Lx
yr9H3fikOS3Ht88i6lfh+M8GWTjETFa7d9eRekIfUUTc1V0+zLh6ub8KLCYNrXVcx5PesMNN62pJ
Px4BPiG50CRoya8armV+YwrVISZsKZE5/BsHKe2mZ/V3HAxOasU3BIqBX00GxtbJfywvT/Jb9jc2
dLgwaNd3VDM2bDkUrRMsV9XFaq8c5ol1FiDRr2Hk7lpF3HKTbijmqMSRUa3d2z4jo1i4LZ64+QbA
9U0oGF0RH/GNrwJIp93pD6iUWUdUbouoaTVw+FMrUS50bEzRLFw48ZhTmK9CVkRToOgpSQrKdwa6
RPMB5pgE/NWlrJRuKnf+6dXtZnkgvJ/em8ItOesBMd7j384pw4RkqX6/Cc0RplJp36js2ag5+9wy
Lx+QZcV7+c9XP6bJjHH9mIbO/1Vu84nP06Eqr8/3ImZXqp/Hx9sVRCocoyVulnSdiYBxYX/s6Ljg
yqdTBISxVak6lRRy09O6/LMEIF1JpfrXg2oNeeQ5Rm+GkkuRE8aEGbbLQv0w8VQmGDooNXU3ik2m
8rLlEPJ8FfMCjCVtWqhc+lOr/z+6cja9lv2HR2pny5P0x+KXwLM5gbAiEqUoQTP6DdmaL4gw8EkL
GTCqwUmp/HqvEZe4dSCz+4XhnbscmtRq3TLWh8J6K1gBH6gfijhPLJNfX9bT1xjyJK7dmBJ8sVVP
f0SlJ3/oFzUfK5JuHjNT/+O3bzm083ZGZNReYIGne6Ui2VCsvgibCip9ayjJX/5YyIhOk4+M56u+
cBKCDIlWHJqT9UXEARqqvMt43gSSBjX8TE8FRq0j/yej4nvNzzmx9Zhwk6328Fv7LzlKR6jPaJRk
+WCjZtc+8HsJ+tXzXZQQnhISwIGBnjf/w7s3PddOxk33MnB1MZNpNYuDlb1hG8C46Ls+oj9agW5i
44r1GjxAUdk0W4KEcr5xwm+SVRLH4T5+nok8u7Soj6FiF1lgj82ufBuJfrJJwuGQNr8QZYB7aNe9
g7aHgYDMBld/wgYxRkDG1pTE/ejMbE4xFGLUm+4Lp4RenLbEHB3aT6nQkkCtaZOBi9BJw1XUXVfh
NwStuDBCW9zzsvSX2EelkCLh1Szp1vs84yjmjUMMmHoN4RVNcNUnsCRi0l8Ls33cPG+1A5AZ4euK
5ocPA9vyuhnvRFk+IXGbFtlS72CoG0v7cxreEjoeTbLZTo54hHYcFrKOe4cNflpLRIDnePWdjTmR
lDjRS7R7OaUHtsuf3GPc8W2lLidK40DBvsJbrEY0XVfMolYJD8ydRePks2eG15Gw0K5EcK3JaDna
8tcIBGl64AZ8jCnnaCUn77GQDhMQJAbUIeJP1ZXMBHfIE/CClSUZ1tnE4LBC9oL/p10C+NKjNBWI
2vwP9oc9jgaHZfCXry0vStCXEBU5doDJAb3B7QlzDxzhh2P646jNN75QqBnbNRAOJ9+4HIP7nYdr
PvTxz58eWnK1JmXfd0MnRJ4VhQRwv45o5FMl2cy+hbOups+6WUjgmEWj2F6ixYWAhGC3OvRtY9YF
jrnJBGiMnodhnXC5BX6Xwfon4VRavRNJALx64UUCRKDx9fHGltw3H+IIzBWjyxmGItCRFREffNsU
YSIAZnwRKD/NIa67k3x5nTjoTrWgCw0myhzzjqs4cR05ZKcP41JxuE725npLeyjwxN7xV6K6Etv1
V5LNJLp3/ScZovjXgjPvST0Gp9Dyx53XD7rI/ogT4vRm3rNIU7J0OMPo1VnvvuFPOFmhMFRmPPn4
qZ9c+exa/vVU9zH9KJYvfQovNC/286rM5fmUMbQ+QrTNuci7QCex3XRWvf2QFINJxtCp3H9582fd
YxTsXKDDDr5+Itf+KpUg2q5Ur9MDiq0ox66vCM4tLlQB3g2UAjU9tE+v/HRV1RcggQwOeg+CPhc6
Chm6GJUj15uVGDAF0iHKBRuCl4LtJJ/VSrmajn44HdZUe4siOQHPjUcQwl4Qt2jpeWuIQLxREftt
h+ltgki7ggogGJs/v2fX8Wm4ZMCk27iloDF5gmvnReSHkrx7SDp8GtM36diSmiTlTdDuCY+rlltD
z2DQzlQeqpM2bdd/sj98pW+/hhHlfdrQx+AAC1LXyhmjBdoUmA2qds3wTEsHe31TjE/wuT0vuZin
Dtczoeg9R24CjFP5zxQwb6DDreGQxNez/puYTndTyeTVOsZd1/oiLLEhz+gSNfnOHFS6BeZK9/MA
5EsroKt46fftvSZ6FUae6eWRO7tzIb31F6DDXTCaun4q6b5iAxQ9f4mXt0wvJ0lRhVxVFgsBuxtA
YmuwSgkSDoMkKl/W0eQLoXRc72J0BRZO821ZB8j7bRMe3sqA72NpJAKSDM9QEkmGfDnJehXJI2yt
noZlktqAr/598GRxyHc6NQDS+4dG2JkkvC0gajwKPFYiM2Xepryx0zsV946D7kEmu2O6VQ4roR18
QWSY9jnjNe+dcXNp6+uQCkstV51yEmjZA/hYF24nUvl0+5ekKZoZGCIbJfesbB/Nt+s1LsGVk9Cc
Z4Tw1zEEVm4Cjx/6KE13/hub3UmSNMxQDHkpRqEDmnM3tfYBiQuTd1p1ZVll1BEEbYpvYwhDurd2
bgCJNyC2TxE1xthrA5N9NUZV4Cl6ThDqgfWlopqcUpCcN5qGXvBg1hzJfvx5HfefAT7RC3Mehipb
hQldjfX5PhoBHuJTwN5RKunNF2q0KALyHuRRDrbPSHnSQZyTNFXblqmC0OnJ4NM/qzKHvxPSrRQ9
Io1iNqKQ/wPtdyF0PkTaNSlWjPgQ5RTca+JtMT/PuHaRtU14SXSChic2vq36V/gsrvXlMrCcKcYp
gkHz9dsiuxH9IZDqSeG/yFu3Smls3MwBQTyswE48UfNm9wg3dgX5s0Gc0S2aAcNN91poPpzI0l5r
s89yRZulnoo4pfmVe1L5RcrTyU6hZZ8o3CpmJC2T5YNokrkd7gIFBO1Z2mv4RnznT2+qSwX1aNqG
ipjPBcY5gnvy0a6vvwMx4gYaT1OiotK6ljUL4wnJj5qMsXwQk6sl08DBcOThbSbH3ycC6W48x7up
GbUOQzLziBZJGRwWeDuhZIE4aB/5BE5aTvWbGHp6I/H89wQsdnrqjztsCgD7n0XZUuIvB7/6v57O
5ig5Hm/AKjn1NNG1RPHbIFSuF7FSKoJad609m6UbPq/qdo2tzUoy36yHCX1VzDsF1OBurIH9DQp4
JunjUsr5YByLbKRvWG+BuiYnQNMJArfxPC6DuEheokoq2w3lS53J20swtcjJjMxlcbMIRsjvD2wD
BlWlFakwh1MPZfT/6OdgV4eYXsOt71VoNJbn5FuHD5/X1L1YtCjyqUEIGQ40qhcaJntFRX9TS/HA
yHdkShBXUFGYyBv4M8kNbwARpfg5cpqc+U+oTDXuhmJTcZXj0PCNW4Myohw3/DUjS+EN3LlP245K
UbWtNP5jI+5LbBopfFLootI1cI7ZUcAo340OebVfoT2s37P82vux8BK5RJp4JOIPs3YYYAXBeTmU
PqAsKDNbQ4iLJOGOY1TAGsF54ft24YZ5U6v1wR2wCGnctOl0+T1lCO2FjS1oQjj/Mf+RIKKaD3fN
9RFKVN0BUGHDaAZjHBMjQszOiq+yAW9v3wrRgjGDcX1QcwCP6x6y6U2MD/qFUEj5H3o7WqFbAH75
b2bM6uP/n8TRbho1zy1Ig9/2dqCrggFuJNaeaToZiwW4/oXtFWPqp7Ifa40vsEeR/1AVSTYweoxr
4CtesTIZn7efSA3otX+dRfcBgcJUGhYpkRehwdpQjRWEjbJNox0hoxfYmXiyerLw7kLgaGJRsPLD
h84s3ZP4bUle8xI5UW5VeLF8C2WggmOeqNsLsZbr8/lDNTohtwqYU9+R9sF/SE4fZUK+PT1ggZAW
8iKHdfU55wPOAIjsMrI50RS8p7bzArf+wCLfG02BPTAY7403b98t5/nTojvfAJ/M66dHAhuTyy6E
tDSHMDxKUWCOircCIro6b3GIzWqkL/pIMjbB5o4vA1Zn53K9c9jSAHVEuRiJhlwezuhBNPbNDkCn
we/dNNSnJ3NjoAIuLqGyPF5AvcQ4/rsj6cABoORfrHhyxXweh/RDowOk9VvzA96liLC7nys9D3MF
5Q0t6k1mBr4jNRuivCihoRrsYM2ZLLHCa8cpikVGHG+jqVxUlSwZMhPb1lJcCh9Hq9YM5NB3xK7L
VTWobmFc8L7KN7rl+OddWiX2zrLtAgk5/L6DH89JbpmqfuJPmoCQjBHTAIB2SuOi1lkyjXTgbk1P
UNzQ+v9iFT4uD0AzXmPIUT9fvvUCuE4LE/5QsuPp3iw/E4Ax8qT+vDlboDd+GJ/jNolVSM582lO7
YCQ6IKgAXVD9A3GW8KbzBUS8XCfeCnhf3IKoRxSBN8GYFeTFUvFsT+f8C215rcP2ODFx8Bc54ktJ
QyR2L7A7r6H0dLOqTXDKtJEgSepsc3dElsVI0wddjA9IOwpi/JrzjGOG/+wtPjCJEjVCFK6g3Us9
op5fuAvOt1lXJleBjgV0fd4yqv1CSoDQ2iPeRqyjoXXcz1pm4UDRrNWqIX3FIFxREHV8hJ9aXGZe
5+ccCb3XZpFqli+oBXiDj5LfQ1kFS3J3uSwPwYJrN5FJtrevfksGMxdgu9x92TSFkzLRb5TthFE/
7AtbHnPSkUmWW7tyRiNJ6T0hZKhB7hYJP7wzDSx4y8WQyjIqko+Go9FTkTRdPyZtes37IDc9hxaT
Lj6/5Vk/C7mkOIN3QxpJ1Uf73OZGTnThv4O8fARUCi8suUQNwAn6sbPQZn7FWuZiFUUybe4EL0BQ
RPqUWnVXibHi6mz2Fu4yMNAZTRUfTKfHGP5O/oXMlgOu/RXTEFGXJV/WmRemjNQufm6skJqeQ4zd
3Boy1LbKkoFgJpgY24ziD2bJHNSZS8hJ5Irkl/4rG1QLi+g0AWcFepoE8Lvm2mqj80j7ysIxTsFq
ncneDJb25uVTzUn7qjV4aNTvcmN+aVnwkCYYNyKhO7Q5xmLSFpx4956TqFfKLGPgZvPs3KUEeVDx
ezRmkgi0qriC6V6SihMoQzuCWBeFdNNXEmSh2VKg9vEaFlI8ZjpWYxPZCe4xB8Zfo0Sy697nGgsN
bYp2zr0+9C0NqL1wbvd3TFcMekPWLc+uWbbtXLdbWekgGlFHYMfI0XrOvVJLrOTgs0wNnuIqDcnR
HMPSETeb9iP/yfC+PzhAA1Un7iepMNdQQlmKnsTFlFGBZWDFszAHiMiigD/yNfXw1gaAUvejAgF7
A1TDCkpF8fe6eFdCuGvowlHD1Di6bZqBFG02oybwA+RnwKaxXCWzUGvNsfU/mS434OEtvJpOeG+J
/wmjkdR2OLeRO5WL0dkrqM8pvFjdeLtbhyxfJMfOPlC605d+RBF+YUcke+eKDghPa6zjq9NTj9D9
S8hcmIYV6gMrHilqQZ6S7d6O3rPM/O0m9NffqoCR9TqYrcTCMzOtuuQlqKUFdqO0Ns7pj/jwakYF
tjPm4ZRR0mvjaBiyDaTMgyCZ+er06ptkhS8/POqbdNWpL6WWvZWyB53tu29lJ0pdr+IqLR1QHbp0
o5MT1JJfRbscUn933DbPcvdAJ59GG9BQQ0OT1v7gOCqbDYN88IUPSYqtTdlRZLdviV2fbjBlqBrk
ubx+1dabou25+kxx2bcJUNmH/0rFVIi58wBoUwFLtPf/EpfYk96CGLhJQ50hOlQt6O5iUupTlGhd
KvPzHWP7ossn9M8hsM8IidQ/7vLONUBSBcIT0zzSzPefYTtmx3qxAL41OwPcCyq51ReFW/iW6wGJ
eoV8Q0hvoZOcJUdCfoTcEAXfyGVylx48Nx4N4ofobKWDG1Av2PG1fRRk0E0RB34OT6jPaQN7BLje
fVgcO4unD1SysXLzrMB4GnOB5gyg8TyHOk8Qo3r06WjX+nAb3+OL5FVi5TtGU6ZKAISVxU9qZh+y
qAss7mZI3rR3Xz17fU0MQS19U68Ewpll9+X4YSAEb3OZRjHCRirXU7u29XfbpLlwgCFzYvyTIwlD
mXzyJVEOgZgGEeHbLRhC0PFqw5NRGhUUVXgLKY71lQ9k/henlQmP8jXvXbyv327+5xZx1/T2cTha
ZLbceTJ1nfE9w1BakBtR1YjosEZiSkZZLA3lOvqZmj1j3zFf9YJ1VfZIa55ANWdYGYA3cuTRq6oQ
yOeDWqJKnBieBmyVZMnPgpI34M/Ean3Lm9e8I5rF1UlHncmJF1HF1yHO5TKiohym69QCHN2a+Trh
AnA60y5gSmQQeKk9nN0ZkNe2uOFzxoRTTpS7XbmSqx1MpiAPnGDVb5x1rc5zWLEddCNTDTG60/Lh
FPAAAgPD/4sXiZouSWCzXZ3GbQPGNDTW9ACConWpfbrXMqu9D/ifTgXDTjXUBx30PwCt0MEaAP0b
1u2ePeNFK7CVZa3JRevjuIkeuNSpHyHcaZpMTIcjDDwqMyJNrFyv6fmOw3PCg8610jS4uz/mY/qa
wTS9i/Sw+/GbwDsF74wiA0UqU6v3MPWeYmmSuADLnSQVfSQgis9Rl2iu9pasSgRWXulzCJtY7mN0
XBvQSTUD5EKPxwNYAwJxUtNp2ybxnSzzq4n1tBKuQhxpc1XveuHg8jqbMcQ7lC2MvRI7UUYkU1lv
jqEi347Yj2Lf+kjkB7nr4XKJK80hTvUevA87Dgqk/+ajtA0AAZ329zMMVFKStN7FsUdfE0Hxy1wK
yE7Ik6xD7PmZl/swAZWqhfuUlyiyrgCW+uB2PaRGN3a7gIr9C5SjBjHbIswJe0dMJVKR+xgKe9Jm
mjfbmWKfgDHydrQUv3xuleS97DNnWP0MGJBAeD9B8etjg9W+9G4il0z6Bf6FMHoNqreFEP9Q7tBz
5klCqXqgQ2SPMdJoyz6/PnrSKFV+5k3+Nn9FUWqTxRgPitsEUvT6yzb+YTHItfDqfWBxnXtW0ldP
mvb2SInp/vyPKq2BHpgp7+Y+Ij3/+dqZNCOB9kem1X2IMKqdYU7bJaZ34DdIsnM/E3Mkc0+e2nGM
kJHGmYFHFFuFJKAcYiwFiptOJ38C6WXTqlZOLbPAiwWYom8hJUjmeemwU5cfQaX+Cn3omOBZUNfb
zqC3/dgGfqtXF98Nz0R7YBkNHbJSC/DjBoJztvhqLHlYyU7zpsHPCEeiTpVUYPrkm9yEaix+A8H6
7ylbbJa/sWPQzRezq9kOkc2iqMGjjWq/kMJEudtfDuFkzNT4aNvYR3aQ3PIAau5C361iRVoPPgoG
26BK5JVe+bjhkk0XqnP1DfKgzDsDI5ooBfT86ue00r+dEPiBwfl372BsRnrJ6IM+4iy+G5Q5RSdz
Y1wH7kyJo2odCNoUPYzlSBEEQz49F7Fduh21fuw7SwbQInp+nw2egkvjxei9qzoCFt9TINIDxzaB
30219036Xpj6BEmtevlDmQOTAbBIOQPEd+U1r93kJ+XAXSpmyrReyarzT7TXl5KqTiu3ccnmYx77
ogYb2FnLBNZum0UUK/rwzf1gyeS04yDGWrOcz20qQCt4t2C5LoGT2pPyCyDm9NXkQyVmLV5/VuRQ
UBaUScmJyVX64UNTwqSSVWs+Ujkv8dMfFNQu5TCgHpwTyo1k5i3VOgQN/WN8bzPMuFEJaY1YuoSa
Alkjkzg6Xamq00F0yeDq2uaXj4du/+2/LRAFLMHT8Al5PPxYt4Y3zsI20q751ApYaNVUqoCyw10x
sA20ILWmtzQKPf5SMDNeFBgB4pGzryLgez9P3LIqhMdXVJgX1QtFVAP1E9ZGxdqP4fglUBTpb9e+
UzxNkjXONwzAVw1jQYNncOZV10WnVZH9/CSlBBFvpk7oHXzzpyxyAdfvKfbn4FHk5oGii/9+3YKb
8t5n+5fG3X8wc/ii+M7rd9aSsVgNJQ6cYpeDvo5856br3VsBbralEeF0v6apXjkm3hCDhh8Tz8g1
Bvjooj00IyIgOxnLidNO9pcojkGc8qXo55h5Da+xMX7uywQFHkZTOXd81Zs5CmmOjZweMI69I+Lh
dNt6jXY/1+QHeJhkcOzecrdO+iZBDh6EdLbTA2uuMdaDtVOH1Cj8Y/iO9nq6+47YCoTe/d8zKHDZ
PMMskuurlLkQDkYI8B7e+uBu6ChG/UYfqwA52V7+4HuAxHJPMWd2kulio1ye5xMYPBtGA6iWPLdR
KHgiD8vimRBmw7vBZtqpAE0KQSzSJgWI5KIYI/EVX3op0KrSqGuHNZJfuDeSxFNjtNnG8XaZG/0d
JDGCt3sCBNH09ZCP7ofPfmq43AdxXKPOmYNzaQ5qIrAIoGY+sMsVjlg5Eypca4S8Co9xRCoENm9a
lEH2JLLSNMcowQ1tmkDOoo1TUQrWlHlzJ69keJSi4Q9SkhfXw2uGULFLDm0lhFTBHvgKWxLvb3X+
miG9Kt/IzcofwCUAQzANsFsDoB7afmE5LDZPCQPuxayV2sRB87/Ndm69RmcnoD5zNQZidYkN2/Pp
Z6yzP4Q242qH0N1m53UqZJ0BYwO30VRwe+iSKnsyKVygd3MROlswMoeDZn6OWnRJm8+D2bLeA5w9
rFNNoOjVmPeT58owTSNZmSKD6N3YNWDa5Za7z3hUlhT6ZbLQY83zak0whwIV1YCoju6He0HM8IDM
7Zxp4QeiAF4LDkm3Yp1+xagoxaWwOPLqMJXLRDsMuUoH5uhz6MOY4QG4sjnZ4aaH73GxbqgR2B/R
IjTNIYnVacGU0T63qwSBUrMpxIsq0sOBg9X12cg4bBltbgd0Ao54aDytf/q/d+0K23YgWjb3aWT6
uRNdb8VX0cMxVE52qKlPSt7ft2Q9SeJa1GlW9yAir1AwdjFQL1d76Otjn4JfvM7Msbs0eAJKA6kk
Yva0U12tVxVamfS1WZV2sUq0jZhDvry3nbSciAzzGtmZtJmXivpml+oWUjNB0Wr8Le9W9EeK0gfN
glYuTuQDmwdglPlutaQAVc2JYrOdQ32zgmQyebrKbUN4pxi8dQY8j0S7hugNRAEUjGhE594OZDvz
cRRb5QX0ufjKRsp43MnIKIeKEbtBKmY0GZDBAayERcL/Kqkr6s3N+j/1u+5rCd9egMXJg0rkoUce
kpK/XNAdrcE+W0LVya0d6Q/4Ovxq7InpK+MzVJlYioOSesG0kTkx05VcSxQNhBIBocoWtEiyzpIl
C/coJ4c2+WJFQDMc7BMc//gsJpnlL6UdRrkN4w9zenq4fOOVVU7wTfgkcbUReGI+feN31Hw4PDNm
Jc/CKiQsJ0Cu56WRtBzt/0FERCx74wWyzPaPRzLtX7iV7MkceUiH4BVN7hKP1ksVH9xY/zPy8g5h
cnm/BBtUbxHR0tfLT0MAnUEXm8B6EnkvgmdsafNSx+rr/if/dzyLKwrUZGpGZeFOlHt8R61+MGlD
Z2AOwk9naxyOBG/LCvYj/c8+FxVaGPXDtX/TAcJfTdYqLP+BQ3ooWSvXUF42CWDAgR+cR+ChxyZc
Wd3hiJz1coBoroAnbpv3sFEwOcgSwy/sBYO/rKPjJqbog05t/ciWYgvRvDx0KbZ5Q/sA6jN+b2C8
PZAPMPP9vQLfsTjfghKbNN6S7eoKfPA2K2DVO9CPt5/IUPvzjQoqiB0srI8IWVYtdFL151op/fPl
L8qlfcm6N4yljxNHrkl/a0Ssnh9JJkAMY6Nkqb9n1ICS7P9weue+9dchnOGCZC/dCR1EqpFJ++3j
DsuIg28u1euLbNeV4T64g0ghpCA3UJxmG4x0rMrG6wjJFmSOZPJGVROTi1CkrnpTqGObSeGTGoFO
Y8uibQnJRLO5+tm8NNSMsTpotfR3o9i8EH+Ns0ShCKJds/ku4T0nRWQqA379P+PMMfJbE1cETGw6
3DtpnePacyLVrvBO/yQefEq29idTD/ENrP0fLStCtJvzbtXZm++kPmOqfzpKEUMvldolSxyqx3WQ
ELV7kMVlFZZyA88Ngee9a0got3kL+gd/XxzAFGrFHKK+bDftUa5QVTgfT6gTiPDY/YEscVgmoioq
amPQMI4ycEXvi4AXj5/kuhPO8ss1gWvePgeO/n77IYf+0oYduG7AZMhEPyPPZlpZT3Bg8q7+dsVE
ArvnYgp2LpXeT8BaU/3p9bg4sgk2qWJBnKNbBcH+eZMb3xdMBG70Oa51ED70RSz751A1YzcVny7f
I5AhaUEjn3g6EnMxBkVbifs/RQ1kGcD/ZrNZgxsl6vTawi6d781Ln2T+A2Iu9iwFs4epFmxYeAR+
2ANwZzC0RMLm2+ya8XDyMMGnb9+SgxX6rCOW0rQUI8cUqhidCFl2IMzZH+Ka9/+h/pn0bKlHJfpD
WxCGiuL+YylGXj5u3x1Dtn4ZxCYVFajfck4fFuwsNEO6LJb/cdPO7K+SJ45etE1beTDthqqzSGGZ
yMxi1Ez1U0tc6kijv1B5v21Vzy047JBmbGkbGWGMAWZ+/Z1Eb6Md3Ny3nGDntSAtqhdsH2iUsfhR
FyzD1+QS9Sjog2mta4C8XC6CeOuk6067tG7ngRhB4r9/bdCrM3C7NG4UsnOODOlG5B+xL+GMYuHE
qX6z7cDZhcEjgEWQTiTGIN7uwiiIizynrOJ5BVEdPr/Cwondvhy2iowAEeKfWj7dgnoeQuVD0GNz
JYDW3VEY7DQ3yxivHCSCeM1Zx1clnkxdI8M27/FNpWN2xpXxrBVW1xXRwUXofdM2STapuEAgPAz0
wWp6hr840jhAOSh4r1YW4u7jU4jDuhqcniBp8j08t5Pa6rX5Fpto5ZIMiVyZPouJ8hzbxFv1OYC5
qHcSve2KV2V/Ul1TzIcoZow3g0ie51PPFieMePasWrSRy/0+ACNAFQOFvhjHedAKQsNomkXVfWWQ
bJVAVxf3y10IOkbYZE9IC+zuQXIawruUOzQK2hErZP0u39uxJgFIYfHnwUtiaTx0lEvqdGXv8eNl
5oEEr0KJEGNd9XBQ0aqxeiYn8ykzR6oLCuJ3HeGtbhOKWDJ8oaOYpUfVCgB4ijbZ8Png1H2uUgbl
yDBQPlDuw9IHTIHDJm1Is3JYboCZ79vrmMDhR2jpt1KYaV1oSAwL0z9hhlV8fDng7QCxyjFRz0C/
ZWyrQ4CnTonJbedVKrgyl7d+9y2EokWbxmblcZbTdhWOOsyK0881JZ18cgP4Rk5P9SK9OiEmrncF
yfQkJSikVTYEhR3uAw/bK5aunscAQ7wnnddS64PpvBJts/fqSw31sEcwO4EkQ7A7Is+fXPJBkSXE
i7HP4Ui0JOepGosGQ8Y/A/ow2b5QlUOpm5AK+IpHRLokNB8ZZ9t92pRzb+WmhwKJlwBU2rF+7sQM
EdfIVhmu7RHtkcP2VrMHOpa4KcngSjfxETNCY3vkZvjZAnrGAekLjglNHvUdb9UwzekmopVraydG
Y4/sPebp1jIwgN44AZmwtGnu2zbnyeVJN2qfxk71KSCo/JKE5yL5nbs1cOEHcBMqb5YiRWuuwzN1
vYXCbZ5jNGasp4+J5XcfwCUcHTjQIiJgstmQ+GVLxV2lNdXn/eOZSJUlm3AxhR7bROxbXEOUt4pQ
H6cUmaI9pVOF7qKCfJHS4ncR8bWhNz96x/qKK6DtDl1412l253Us9PW9MrVQGT8exJ7dxCVGAK89
HTg8ngoK1feJxabEO2nIqxWRZNmqUgmO9jvW8ER8Ot4RTk4pkSfNbbQByePEpkcKD7DAJsdqxgFd
fUMqKzKSSl3GnzsQVUdIq5TQE1NPFD4Ec2AaWDUabDTJdys+wytt1spFnl+R7rFQPRE5a9JRIyZA
Mjy6GVEBpbS1rujtLEf3S6fGFcByfyrA4d2DM95qkwpPMNG9AdKDBBA2h6D8LJlgEt1wrQkqGjJB
jP24LUaBxzmCh9b39dJOEFPAKelT7TQ81DD9lUUWdz7EVZ9ewbbMA0kI7GbWiEdBda5tbmPNFaTi
K01d+cnSCaR3JYB+tNuxLBui0hQwMN+B9vfnH7dYxVPr8DBlBarJEQYyHoxZtI3xxXfZCqLaEZ02
MnPW5sv8MkcuIiA+CR4ld+G7OQ18KUzpLJVWPEvyY4dAlhu/Hwbq/qShi3m98n7SxLKeqg5I0q4J
DmOBX3g78hQ7qLASP5NQQc3JQx4baay2683755RtcwsJiU9X/lVVY87rHzErI/IlFtLIelfZVH3k
HHq/JXIm7f9zDze7YX0lRBYBz3dwkFasNODGpp3H932VbDnrhqIRaxAKyHst76twDzANiXvafSSj
0+eu9x31tA8EHL2ie918VQ5qsPq0kjPiznbmadQjY0KXhSmcWvlKilIY+qH9vmyNjmIjponspIOt
KFWJ8dOeY9L0Zrelk3eJCKMkod5pB03zzQTdSVsb0vdVemTYSrMAKeqvvzAXLehXAr4H0XMOZZvk
nhtEktPUyrWBPs3kZZjlbI0t45wwKOARXJ7rntACfjT8ZXBHUeidLMRgbbkUxw1fiq6YjjqaKE/g
XxYDk2nMTe34MUKrP6qd1zU77/Ve2zvTeierWmQ/bKT1Hxs76/j7pgXKFfYO94jXOZsRNziPMjpX
/5FI3y7VFo5fZlTAlqrRtn6hKPEK/M8Fq3i8xxRYy5w7GHiNjVhGvqdNi9lp+R7Irdwmrj7l5m7z
pn/3jzYxQFiUkvzMsmYOi4zYLvm4NFcTkzsVxy5K8X9iY0aC8ZeeTZ6m/6peTypCYChSJsUEHzm0
AOYQ7r9bji2UxSOyZKclT76biKuIMxnKz20cvwJSge1yuN5dolfbk4xWNpRSkxiwbH5Him3SU0TE
6+4kaFqNObd36GuJZLM7jTj6Lobo4iF9aXFLue8g5TA6/4qiUp6ebBnSjMkcju4UxAxY3k8o/4s4
OCu1mkxsiWZQ54St5wsRgjj6EMXtJvhIQJ3h1B5KthQmoi7ol6UrfBijGLjA8ZpY0SO5W8jUc1Fp
7uGv8BeFTkgxrTSMBo9+uLDiw4uyQ/cmwh1uhpuKvUqcgO1zCltfjEmjMm4F1Syf0Rb99rgjmuSW
Ca7x5l/hu/EAU84bo7WiCkq8A7CaxZy1KIWCex05M9Ok15zHPf1ij4pKnUNiK10oKtV+o/GwqbzI
dbhLfp19ZDKR2ptWS8Y/tFxhTffdJWA2qRQEYVkTAqc9p8d/nNDRCHI9eSY1UqjcIIFzNmC0kt4k
eu8lzkLS6VbWrF4aYxJaivfnD0eb72ZMNTl5vCJKtSy4v0o5UX2F4fbw7TWC+KAkP79L55JCkixT
T0RjTyo8qx3oDODvK21oxda55oI2DZqk57tZHexqWWECQ084tUEL/wKpx6IaFpei6CukofBCxXTm
Xa9cWbI6fW9Nnp2SY66C52XDWA9zdL5W2b99M5Y86xVDbUB4G5E7Ib/bS65JXS4GOBZ1z9+Th6wx
wX3uJO0t97748BeEP/8qbr2IPo2pkyjJ1f8yC+jzVIVg9fpKngvJ6SjHLV33cFFwo9Xxqx/yudYp
WrCsxi7HsZUsnQW1Ox6BVzcWAofHFcRuej66AG08YW+TRzkhQo34zM4s7nDBULsA0eveMCvfGQ9A
ZngvDD9sVjo0uuWc2N7q1r08jQpnWGMJk5YWeDOjaxvGKgbk5SLN6oWfiv/7m6Z6f2Zn1Fmr6XfB
njz+yknrQIan5X+6a2xa5hK/3cmtF6aGD7/hct59FTD5uVhZ6skYQ3eQ1jTb8PPe1y0d/ipM4N3Y
JDWnV7VUGK5cmar7HJMrG7jDWZcEKShV8NhSQ7OsjE4jiUrfJ1sq9WvvI3B19JD3mmFF3rzXJLzk
/gIKpcLlVcz6eTBPvfqDu8ZYII+vXnhGPu9tHUvpNsrUeZtBXd2WZgd50ee3cRjGw1AUFgnQwq3g
7Vz8O6I/QlHjJ883qC4P3Vbpoqja9YJOFtgyejACC5D4aXjVX6fmBGxCZ6yXv9bzf8Otylq3aDBc
IGtoarx7nQjIsQrpFYk7gp+SyQR/oB54P6PAVDIlFbilM4hqSXW6XVqVYqpdgDK+yCUPvXL5FCt6
/jCWZajs2LpUGqJSbTxm7n5wS/TatCFtHfVz/vK3TaBAUycWLgfn9xEb+4gZYoQkQjGEH7Q+SGIj
kPi8HRienQUyXUU4lNnZHR7sgI1abGTZaMCVP25of3JgmQUePrt/0behmKnhe16KD0KWUD1WK1Ve
fzpkLiiHVTQd1do2LMM5aQsdS7vxAYzganhAAgsI7SpAkO1ornHI80ZXzWlsgE9u+STS7xCDnhw3
yPmjTPnKJNXL2MlKyFSijtxv4qXHSUdOCd+a8xT7iF5rGuqTO6RKn8JoIGB7WO4T+VwOXvjd5zkX
jbcoAuWcuP1cqmewV5iZMePRtVQG9waYvEoF6KFIYeTxyPtcBZwGOc41pUgh/u2+r9635MDNyogj
FFWiqfktNKP4HXy87sZ8gw7JKUmPaUBwq0ZLrJciBN/vvND2yjnmxznUaDUHFiag9X/gEditc3Se
VSSdE2irtKvYr+wILmyM0x+T/CNjJ+UGXyO7EUA37YV3phcycEM1qNsjtI1Lfie7yDdvQ471QFK6
x51E5/eYllfnIJfy0WpTY+hgdAXRTtcUjLvbuUzeLo3uocDA8jAq65L7kXctWewmAfPIO8rX5u2h
MiZHWgZf8hzorLb35ZbaDbAis5sO9EOuNrG2po+ulBH0dhmFoSeMTrI7QP2kmjfOiN8/r4A15fU8
FKArSIA/Ta6uGXo9nvIjY9RJnoFJ1+LIZNJitXyeoEhVbdbMkdJ31ckqMYB8u5TfJhjnz99SdE9a
rd3wDDycenvG34dHY2wOq2OgC/sBlO7Allv4fnSTke7CIhlVkeN9s8cqoxrYR5T+nsoKhw2ikZQF
yDfv527YN/ldGs6rS+BgvOK7T1xl50ajHt6MuCSUlb8FiHXSalyZSjlTWNGOLtN86K9Zbrm69dFa
Ag8FRg/NipeH8Jp14T1h6DsQd0c8wK2nkM/0JM9dbAT5mX3y5hoEzj/G+l18WEiiS44lCb6fqaVi
GN4AI+0ND4vkXqjTo6MIE+9ZrCOunow4To2Sb+ymFFTDZdkOknHItahaX3kH92CKrYOmN3v1S9u6
DvlaIjdeK6SjAuDr4l2gL+575XCueWoWGvx5FMj63UhwT0bcCXqw6shxgHcn1sf/VlWIzkDY5VnP
cf3UqQTFLhxqmFl6eNhbnbGlXrQayXwdkZWejRwOVlzeOYQywdn0MvWKdnbeOg4rMVdb7wNC1FWI
navDhXmmVWDx/V7cRUs7EDuWyKN0kCMkbhlJFO8+UAgnCJg2PNQsDWIWVTVeLu68Omqo8lrcrLZu
X1F9zN9JfL2iZEp6HwG5f8F4nL+Mh9SiWV8TnCom28KeTzVLYEUq20kQyQuOPJ4Th1mKknYx+4if
J5JqQJbu0ujJ0R7M98cSM9JG/hwxNhB8P8gHVweR3+OIg1qD+5iWXMoID97hdLdyP5UEsN1TqGXy
Tdod3YwCvw9LVj0kX47iRtf37W5v9qzuGHrgCKX4UHv7KzSPGq9Y1DHB8WzXWzuu38MrP0MPD2Bk
82ZQq1u20rnvMTFs7diqp/n6blVuhHn1Zo+YgNcgRrgwvP/tnUJu+9Ho9WmPI+hRPwJR6Sasax2n
iYPaABxkkywlpzR6sivPlxQTOgFwpaFlCqT2d7rSnP6eaIoiou10KS+JxVBy0A/B0pMNCCzUWtuw
L/mJEVbiAJLvFeE+h0mlMBDVz4bM50aT3AZg+RNJkWW+H2LWh49X3ULM15Cfnyn8dslk7VWRHC/r
2wMdL8rYhsqDP474CJ4FZ4nEz6lzGpVUF3GcEkaQKhWAy053ahRGgNczTgk2u7rQ9BV+b2StpGWK
jiWcNV/6ktjU4s4vnMTvZw26Uz8qRq4yJXPCmnECVuQwjvyNgS9y6FIjPeqeKGXbK1Uk1kFf9cFT
hSkrvP1oBg9lKvv0UqZiG0EhPXW9O3xxoV8VXQHOck5aBXzwULE0ex0FahHf0Z9ibNpDJbq+Qgwn
zNMoo5r1X3vvjpo5c3/Td2IN4RgiAMlzCmEo+ZMcjLtar85AEvD/nEVWCJVucU76sFr7MdV7DY4B
fHzRl85Ma/hwvdJ+qGXH7JD9ICEr1Shc//uy6OMk8NRmQrVzhCxbf4sBPCLjeIiL6xpIGXVGYJJX
TPXM67/+IAzyOzKKAJ5TPUxRi3D+IyFww7PYJV9lnvJsiDkXODt7b1c94IVdPNVxOnbEx3DmXipH
e4J6+k4X1YUOltGkdP03xpI0eM9nYjbELfI4JzOMlFiA3U5oB0vumje8G8oq0kH/5OW7Dkoptfmy
gGw7PHNAZGLT2/ZsuAQmDWzjQnnhi2BgPURhAoOhfb8kqpgRy7WCPiNiCoeTHcya2XiqKKjxRhQ1
YiVb/UG8FOCBRZsb2R/cf0EejkUqHJMdt/0bwxaQhK+VKK67vIrzeQOMiMHxVCsjgVt6MZp4W0fD
EsEwoORbuz4amMl+cpTZ+uaCV4RxAoBuzrQP+7HM8PdiOpuOQB8QkEdkBZD2neBrKfw9dkPyC2KK
W/FqIopMTSMqPlm3lUrb/OjYaW8eCaiAbp9TeBTvGHm0h5eeFt1vy9skruxDZ1mxRLm8U1/I5KHZ
ABhQlf/aLGdZshJRiBhW3wqop94pJtYTkQb5nTOS+j0+Pl5/02fbtkBS3YHguh0CuTQewgK97R0R
V7RckxCtrUP/R4jcyIK0NZ2gZuk8g+s0AN90gAdG/EvU5D49yI+Vi2moH5gDt1XbvdamcQ9J2qCW
Mac/b46TcqfHhH9FnN13iE1o6iIABNdMq17XaRj3wp+pdMRBM+3FJF7zqGprsa071IHKPjr3hwuP
QTpLeNKIzsKxv1KH8gyINXmJLvPC1NgQj8gtaUO4hoj7RBOQYfqh4/LgYHV2DFDTJGFoBuvnnC1i
vTgbed98xzxvjsf5KizhbhYB6JTzPMJQW9qNkGItrGH6jOfzhBRRcapJyk8Vfzov78WVKXA4+lwu
qSBR4fKBVIXPwW01Cov93ggH3JPEQDx1HNpd4Uz0kDaIfC34Cldv69+fBFtAavOwgJ2RpnSzFqjm
syaZHIvPx+d3/dCl8UryYc76NgdkPMnAIclRZwoXI8Bh2wCaedqTvt81KpPH5+g8ofpGD44PHElF
TPDZT7xkq8YesmMjwXjOleLJ+0FJpRLq+Cu1QAwMJmZq16ZAjlxtzcYT2tZqekpDKt0yI13/3fVD
b0JDYabDnvzl5B9bVk3+lPxuJXm7UL9MA7xJubjqI6QnzdsJLYb5hvQ9rbAk6SjOf0xG1yC6NERe
cm1JlrC4U6cUaiO4rR3uXkcGtcV+GJBraJzQS5KCrJsxkyHUBnrJ+7ZGEVx2XZuuAtgObm1yfkx3
8h2+GIJWpEppVHEfAh228EM4nly3CucJ3aJBK9tKydbmzihSf3C5C77dOc1p8H5GBTR0JA6fwF8Y
u3/bY59lOydofsF6sosLE31fBOX7804tWjUleMZ/Tj2MWfSyLak1Vn5i6MP3lD6tf/BDgZMt3AIl
KqNhITtnU1IbgROKxWk1Rijeuq2Nneozu8z3wEacl0Yw+AdHNU1JkmhgEleHX0/sS9Yc+0mhVD8R
nm8rZWlNLm5I3cWB+n0loahOzhF2yuId2YuLYsifGnEgIEOljXlz2jaGLQnz75oyU/CmD4ia3kmv
UM5gx+Wf4o3FZz1SUiKn94ojXFSOuV7fRtKBL/esXVRxagMhuykPHkpHLSGhcnLlwGz0MUXbq9Yk
DsgISMrzRkzgBfUafQAKa95UkrmMmUDcI0PMBb+VeO6z5V539PaJFCvqKXmJF13wbYet/CTmCqzx
ApovrCWuRH05f+VWKLvJ5LQLkMJiBjAY3aAfNadrDWfZPipqgfa5s6lVvDV7Cv20Ew1BkdDjteUa
qW1AQ3iM0kgzUc6nNxnJ5+7/4qZfU6Z7k10HdWYdtQnn1fCUxdTNItIIgaqovd0bRcoutc7ME6k3
eEwUlrGs7tClzPMidy8H2c5qaNq6KJVJD8Pk6EY3ZsBky74leVDpo3qi9S5qYUTEN02rF/v1y4Yo
lSvv9UvqkZcc3ab3rRb90cblH0fiWvjXX0HlAVil8nO0D+2isf6tnuy/+F5ZgO8IO88hjNUW6uCj
OnLHESsAYsZ9kkiZAEz/vE++FeRjr7m6jh2x+HvcdWbRjTTxjOKor2wfT0Hs8+51I0hIJgNRqp0v
shIkerIJJS6cbC77oQ8jrcujJzqYyfy8qT7wcDpUU77l1Kxq3YYMNtXjsuP8j3GZwbNJpYfBB6aG
6DIwgWSjDQOa+LLAtL4ivcxHZAIlcMxBaUQmrwqj7mo+ylbd0gD2DhC0tMLPsH/+8Upjvw8Jisms
Utyg0F9ZTImsnBkf/zXIlAaX6Eif9BRz31fojpMAu4PttjhJbl+FeLR6LSxvo3inODO35MM7O3a1
woSuQiw6dt9n/6P2/kqgGpnkRhnQZicKldckZuSDx56GyWUXjRGdeOtOZkdIx10UgAOttUfWViJo
I4eZbRW0bGcCxXtQ2J+NxCDciqVWHrZzDSLQfhvktE4zt1MM8fqZyXlfd4jBl/BjUh72IyHcXD8n
1qQVi5wHNlBNE1koCgAZD4LOJUeACmHRgde6Wnt8B/qnl84bZXoJP3BZkIhGevxQqSU+YPoW0FG8
YzfU8hYKjHnq4nL4U/+ouWd7CzVljHnCZ7BkztAzsMgPGLGZM0LvTfRyrp3kRAYewW7QSEMXmN/8
YqyFNuTfpFXnz6GNdJFCx/a00FEuj2zjp+qXJ06U07mAaueKv/1Vxp4OkRPD2O/t8n5jiMvb3lvF
dtUJnUHZx8b9ERD3fJIf3SKhv1xucd8WgXCGJwmfSqIoFL06A8wl+thg+hQKvOug+wlsWlarJx0Y
fv32uQH/AtKuC/lXdEMhdNbyv3l2vS31/P7+g+hIyN4sDPcg0yjgGWt+Xlzb3Dg1MB+k8xf1hj/T
BH7SfMuT7oz2BFegJ09Ky6GHQ6IjjZLrGlA6z1z/iFaf4hpSNjOOtWcwnnXaM2N3MtGMQQjGuK8f
K4um6/i+QmtgfhEpA9z3U+/1l7Y3G4rawrVRrAliZkvwB2ekmQ9/EAejBl7UfVhzT+zki32SqzZ2
MkCKsHPT5CZ2X4dhPhJtG0S2Ty3RpusprLTZly1FL5Lr/yStCO60JrKlqfbuo288CdPuKO3bb6AB
hJhax8FlBw5Dc90Lg3vbtpz365eNdADszwy56Np7vV6qQTcfsXZJ434ahyJfwcMPIWiv0pzbM71b
WOPhhUqOUyutlt4I+ziZCAKy7idFHlJQg6z9SOFYmdZlI6nZh+yJH1FuErRG7vSF8p/kebEapQYl
+FMZCcSF9EGel0wm/CrsYiR+qyzUBoZGCAY1N3t14G278zlf9EfPrZHkrXwa7PnsvP9AWBvr7m1a
Qqor6cycUVd2RLLTwVJ6ezIrsRC4f0OnvH1i2NsifOv5mM1J1kLEEuV5R0ZIxajlyA7/oETD59NX
FwsOiXXfwhUhQ6gB76DqYw1qJ/NSPi3ZJQoAH+obye63U4sPebRtyoXb44NCRJs/Fi+rlt45KEVw
fI9EczCojNKAscnh43yw6uqO/vumczB00PTmR9C2J+fW+sPrlFM7xOeu7mnho6QiEoDRRPbxxPkh
tS6NCaGpnC8HdVBfbTqw8rs26Zkh/dZWttrk4MHqs+6TIxn+gPixybfybBlf5QiaKbffvSR5hBvh
TTqJGLrrWPxJz0lfLLxlJjd0i0cQReSh/QH6CIpscEwzK1dI32VIpgq8tiqvyIyphgXK80BxGN8Q
sOwHlJOvACzTt/Mt9GS1YPi+vnA3Q1Wft9QWpHI5DwE8wV4dh0rk0SAZYCAvja8EcR74lq2d10/B
jAfbhyFYPOzapLaLe9NmysPrMp5XklRfMwzVO4j0c3aPmFTLRYIN3Vcko6Q9Lvbk6zm8RcDlKww+
uKhYlERnIgbcGY79S4puTSuNht+Svehu/kn+5LRvjvD5uDH1o2Wsf+6sHoK/uqf4iajvmTkhEnxR
R84iUoBc7DX2udYwIRMJfYzgbOXQSJB6RHCvl8U0xcDBc9hqZoicwBV0G643oP47TaPmMxB56pTF
lCIfYwecw5kpIKk03iQnJHHLIPUXftrS3+zNrXxYWk+qEREVhLshHf5mFDGa1EICFW41bzwFNptF
FGxZA3CkYDuw+YV5QaHvXU1xjK9UIEq3U7S+uC9+nKyQJQCy1wty7s3BLov14ChtQUN42phUBIrm
yV0E6gSNzn8aaCJMX2JoOmWX9CZRsFf/vs/IeGeo8F2SPDct39EcJutxpF7/LJus0LQjAMKpaJqg
OU1D6znpwb+U811O4YkhPQxT4p9cJFuRbka2UvVvexAB4AQRcEGLA03Vo6LOTEMRvfrZzewbp0Vc
R7gznIeSU4iRaSndz3TuLaGhxQzOpraUAqPMJoKGFEi93Hypoo/w2D7xUi8o1+nHyLAFKtPxmvCX
yBR0k9V2AGkgeHx7rWNXI92hWlTYY8joei5N4wLdFLbQn92GmL/OsEkzYAEqAZZFjSFFfGsjT2FR
SFDjlO7ccq959nJ+vBaL2Z/lVKYCQ3kyqwB6nhClL50DHSgnw8i2j7lP9PklH74xnMKsgyrQXMnZ
b0OOZkPS4RdHnH8ZUgpIapUIlC9eevTjSwRtgQFFveeDlsrQwa26PmiI9eI6ZQCWaPauUf29+VTx
YX/BUa1xVty/knpgXLpsRjY4OsFP1d2SvbU41L1Gq7a4QepM+BGdJMDy45jmdHUHeXNHYdgSDRC4
ciFweYeXG9YWJGV/I/PRdogdlcSe+WJ5h1JlefYLrjwG4DuUB5enyBoGAI8PndwXxp4djdkwqkad
ju1WYIsqBw23iCtmnHCWU79Z3azpIqG6Rm9NHAcPfo6xZBQhSxjpxwfaBP0om1F7bAJbGJzl9+Dt
yfW+JlSroHlmT3x6MdBtz/O3gPzcHb7EmycmZh3rAIcXdD7UITv331mARBU1sGRopZIUwxGbrBTU
JGshLRLh6SNT/tSIyThWeiuAHjTPSd3NQKLTWotMcTYrjd2oZs7l6hFAgwobYxqiKRj6hHety0tL
FPLLAMYrXW0S6SORUpE+REkzBNMuB/FZS3y+ddgcifZieyYDPp37kGsKs8zB7gE6M2ZUSsNq/IgU
U0HzVBiLzd5yMBF3yy2fFqQBfGyVyNtbtYfH4mdIeHd6ScL+btLPMOI+7wid+Q4OgRuquSt3tqdC
dNH61dOj4+ZB/xGQeOLGUKxuC/mmLbSCvFVmWPC8ExVmVbIKaYiKqy8Jkjisv0S0OrmA+pf3dNj+
hSxCmW77G0UcrguzA6aRgtTTCaCDUlrr+RA3vMnlsB6pTNIHBXs+7C7UZ2i6sxyqfQSMsVwdBLzz
7NOu32lbYGtD/66ZjyhEIRmMrJAnUdYpUKkK/56n+hNV9qfe2gsBZB2f8To5Luv5RIgNppME7b7c
K9j4GqyHfQV8nFbzIfIZeUrPDn3ug1dvsnyru8l2dUeDCUxnhfdV/TdT91jiHTIX/2P44NboTflo
JbPFyXS+Gc7KjBpOPJSYRI7D2Og9pcUJNcSdrzYfoe7hOqZN5+WEk1tgSvFHj9sFC8ikQB2EFQ1A
Adw31rTqw+TWx0hVDwkdP0+3Pyasebiwj4swx4jwOUtAr+MTtU7HIDeg0CpPAu6uBJwf6WzsTgl8
51UeD9fKFsq1G31UM2dpoiKbF0xBps8XlFDAzkAlGEbu7GPogFz8XOFHlwuTTS00UASkOhxzBXQ+
WXI7qGu5a6c+GmCWSq1Sy9kUEl9U9kqzjklfznzfgKV/Htq/+lr9qVnPEjQWne2nnd2E8SrnE5Kl
NSHiLtiGKb/GuApHoUEQMUWxqNcCEXkaFidWfkPtE4XK7/dQhhHOVV2ThzdYDDFIFpi6vCTMLeuh
TfsG+kc2WvchQeirYBVkRxHnNirsrTBdqzSOm3GLjNyInZQSNAWw1wURtdJLgkdFd57L3JuwK+0q
SeZj+AwfbelS71Lnmjk5qM6HsJq9VFWdvG5aXAuCASZ+fBvuRT6uwpjKMx7sSir1ERnErpKUMeCR
geNPtdw294GY0JKUHQWZ5Lw8O2H3KP2ZsMgCg2ANwzjzmW+Rwb1GeqYMbsgzblszN46V67JW/dN4
ArrEfOy6DwO4UbH/x+TtAh0l+pL6bnOAFeTF6E2p1MFeJi7336c0reZDPVOq2Q20N8bsRdv3wa1W
fTsUAx56M9Y7QE0tBXz+hEPpW9ccj9u+Jo3o67cuFX/g8IfKZITQfjJHNd5A4lGqzohFwdMYpOub
G7jAep73P6ZCX9xfRzPl4Lcf3v8PH+OCLnPDv2Rg0GddhSB0NtbwKpvDYjoCyqbAY1q6NC9oHzdw
HYwUvB4LmJLD8m+mhD0MZlT34g8Mt60HKzRnyAQrgstkr++Xy9qXVBjI/dggTY4sjtoj+Daa5cKQ
t+CfdBN5vj0Yc395B67/i2beXHesDnMHdL9ZOv16YfPPuDHY1YWmQhMNGn1FMU68GdcggBiuJmc9
7NLQwVYQh1YL+Lg7sYhCDzz/RkrCW5b17XyXWOyazz6nZnzYPfzEYXLA/EdryLZpCV95aOS5ya+U
18b5y+U7rMlqQHB8Z/JudO6ahv+E+8pS3YuCAErOWFgdJ0OV555lo2PgMl7pNfGQ272P9kPe7QD1
hi1/1lbRv+5eEodgVoas1q38eh44nWWDMROI+wU1/iQjTEUsUfFJb+CLO8ChBtIJdedLFfwGMt1h
ITGn/s9AmLOihpVcF/1MjKOud9d6QPDMLWG/NytfJ2tlmhxTMDRKOWqUsjYHF9FJ9A7gYW86kWRD
ICFXp37dipPHgCPvL98NnuXlg+ETtonF+dOhN2oMqvubjN8BCntIm65RrCGpzays4ihiulaO1pBc
u8cvdAOdI6GfVoN67ODs3LnHNd8YWeIISB+jacteTQ2B+XKjuJSBbu+UadkXPxubda/P8fijfDZI
xISP7+ptowYJBGGnOGXEh7SZg7+AEltUycMvHDDq5qS62mF93lZaZ/eXtQawWOczQce9HFtAIPcw
kXL0EcWwU00i3HN2CCyW1D15PRh7UmbUt9Ybny+pqqbQsYT8z8Chjwtj5DczNlB0KFuvnuAF30Ez
rAfanrZOg+phjPbkTsgeVUstWZ+3zRPxiqt+lzxTN55PZnKxXtZp2LjcPJVIvpOwUFI7qsQsiXza
kCNFI9NjxWDEFEHzA+d0BtUNkACfMRlWxIlqRTULm99F4Qx2ooxmgXDRWW235ACm3ILddzWPD37v
/9KTgR6LG6OXXnXHbMOxYmyGfhqHY2QAoUz/3OxtExWNaXfjel8kURbtfYQARaySP7mfYaGoNILl
Do9bZEnpJeNraUYrricyH/SE+wIwzr8xbzuoA8hcrjKrkoDN7qgTwnURR6qp6gmD50oGTHOTGJI2
Are1BWQZj9Bpxiakn1+ZbZE6dMZZnDu3bd3OtvK6ISENomWqbQmyKst3NvNvxG1hb0ptp29emnuw
iEPbTfoNOCIiV0Cle/KoF7XVLkoyz0Tu/ZhBQUjLmdWXR1iTqQ0WFOwbo0GYSR9AlUY49wW8pCpN
r83izL3qmPiLWag+4lYxWymHewuhW8urk288JZeDQd+hPUCsk2nRfetrGqy+u+j2dwrZreHJOUYu
pOqf0pNYFsJ0lpXwYaJDSv7x7a1tAR0UmrX4zMAa4JM1AT0RRh9h8SvXZXb1tf6yXrlaQy4T6yoR
gm5ptvC+MaRjU9rc1IxPV3KrM8XF9ExDVCqymFmmWOj8MdqDYnysfkxUVaNSiyuBfE4768S/fM/b
4ylvINTMh0CuyUkMa9zUWJvxWEewdaWmrXe/OHnZgNGEpiGTP8NSKUeNiVRo1SDgGi0TcI60bCu0
0FKCDQcURBA7yOIndd6Kua0ThBgGe6Caxjvr3pEJNubkGfoR7encqa3aqvD6VXGRRsN5WISSUTk0
Ky0QUdnhgbqdshZTc/kzmIfy4v9HnBaa0zqcQxHIr7AG0u5NvAsJKx1bipmaJPXw6NoLr5nDLoq7
GMWAiYMEwPQ06tiALQtro29ntjIldEJIysgPFmMIflNoTPjwnznwl2qI1hBMWuVserl5o6vxYei/
gnn17dSqduVV1ds2xDgTC7jGGxelGfKpAYiqJuVuUZCS23TYa5LGeIcsFqN9Z+MYAav+Q9J9ZdUh
Vju/M+hmtLsQnSrw/fPj7nBnePlc4/Tum5bRcpYCeacnqtS5BoV7bVrxm8W8fx60gZ8PkVFsqEEF
0PxpF6oGkba23hMsh/VIBTv3//VQ4z8LwIeKj7vxAwugDCOHXSge/8WOFi8Ypetrg2NrRfa3YXBd
M+DBkmpXTZGu0Y0lEH/l7E70fwtmotxjFvFbfL8o8k9F+sjtaQou4+XB3c5WzVQ0oE7bEeBoY5Rq
YVN622LTbTIZZmI6T2gwnnF1aV3zxwv0FkSd5L7HeLYEfkmM5EeNOr2P2pXIYRrVnuZOy3JFM8TF
2NuKC7mcynbZ8dh3vcrbtV+KlY9uHGtYmkZ6tJVtUc4VkCIqgWYBO/EMqGyiChnoChRL4OOqqjis
021HzAm4d3FsG3XZ/z9MoJxQVLlp3zb21SgnYpOh2mug7zsww6N2LzAwwFdSUBqwjEA1uIzHWz6q
tWMyx5vQ+IJWitgBr/P2wd/NnvqPmC9MAsGqaX/oJrr6eD591DsnKRaI4oNfXp5rzruLkIifVG0G
aDcoKHO4tIqaoSCgDKf71duLjPDfkfhpDgKBpATBNB3xpiIcr1M111VYFsIN9HbeQDHIIBxgvF2j
S60L4cB58Vfg6X1oO77yALyBjrked5b0qrKOfXGjC7AZYue+HWEa1Dp10io/CDhNLJ6i0xdcElkB
OFgBvJQp2Hx8C0x9FbM1qYcqFfubp/bPN8T/QHjspsuXIxRjKfGouUNfDqdDGYJkFazopqoFLBSA
vuuEIXOSda6sElaiWJVB67LYHV+le3oXZzO9gJ+ENsP6rGZX1Qn4R0Ix+gmbGpGwxgNCZ6XjnR/L
VBZCfc4BeermrCE44oeHFvc0IR5SWYjMWk7qUb1vwLwF8htM85LX3BXIJU5TkRdRrilk4JaHs8Gz
b1FU53+LNlJPP8C9IMoIQUcm20zufAhAO6dTDsyrYo8gEkbjBZFWElxPZj3ms4HNjbpwi7aZlViR
jeqaIrN+44IGvZcCocZHV708PgE4u3cvYXPhV5VOxW7k5Oqt7ZrTcOtpHqECD+Wblk4XpQ2Ok97P
JLsTXqmp4E5VuLBAGTfxSC74/MmCYQjW9F1UvZ/XWpZvGfdVAzA7Ac2HSvDzaZNzOw9YLT4zfUwc
3D8z5dQutD0A2D9lI48GLXaS8HlK2N1woAS3gJTep4k6CSj0477JLiuhLeynAWAf3Vqq/ZzOPcF0
qPmBWAOwdU8bHl8pWlkNo4yzGxh/nnHzBLgN4kGl8DM+VgvoOZyyTDZh+PHASMfKs/TcGzO+M96l
0bH+Kq4Nx3KJRiaIXTrLdNw0HC9LSAQ2CTE9Z1qqdGwC1eEkdXtcXOheF6zBxfVwO+JmUOpy3t1i
x8wtCGPORaSqBE7waAQGZ9x8Q22BSm/eE0GZuBi5QpA8DdzQxVyiAIMMHArkygVVeYEdxuTWpeqP
B9z4PIrttafQh3JBQ+CObPAzx9Vj83zXqh6kHAqZ3iZoXsQsV2ySox+Tqm4yyjc7mD/JEwa2o4oI
MujIbuoM9tcYhOqcaFrrlHR0K/svRSrJCTo/EfXNFA0BHSTb1jlKJBNYG1rdypSEs1nB3Ruswjt9
TyejCGrVS1W17fa630D/nHNN2B4eSBXyVcu/TUtpFGA4IjiLTMPWPBwLfE0Eyj+Ym43P1dYJ6QuC
0XWUlwyzLeVdV6ZShCS3wklQFgr+MQYhmg+2rb1oxVECB/WEUl09iG6Xo0ZoHvg2T1AAgTkYj1Zq
8skAaHu+u3TmiM0ZFsDXwuWZMn1yc09vtgpoeXNF2PuZyoCcWzlrhWy4mIp1W7QrCEAKbar+72gV
xamMptOYHclH40RriCj4e5Qa3y3fyFZrB64tlk2uOASKiKgJJJoDNZihkLhIQYzJYpAK2MN6hXee
ZSGyhMwzsrASyeYscVY5qCsM0lj9oVNridVCOc7/v1k/ziljoQ/VUIyU2JKERR9rL9mfN2OHBuD0
+cRsaK4md2/QIHIssC24DoiOZnmzTHOo25Hkt3nzAB4I+90L2OFX6gCBiCTDKuBi9G8+q6fWHPOW
YXMufoJ0HEmZ/oTn7UQCaDpaTQCE6qLITQS/maTwS0N/0QBSHVpGBH2PTbxPfGYsj6xPstIQQ4Ro
iQFILqTAOz2vbTtNqXdDlEibnCtEsytBqJBEfZx+6COoNaMCWDVV0+J6rQKNQr+fF+456ebKYlTO
Ufz2+tfzAdBowd1be5Gmpk42vfA8hySZUoHjIERoNmiCRLCj91HQv0X/Mg3k0dcPTAvl5jBqjUAk
1HBrN6pPISrrlA9cBp3Cosxucl0vJlUxTfJBcKAKy7Ha6yloJBgNaT3jwZwwKJyE3Ufby4yvi2+V
ZCasfk2JUP3QuiqIG5N3wcSiQzKLhsvh0vrJY+vyDgb3rKiDUFCpvBnx4DxglJljGJ5RFM6mtU/x
7x0SWfCHrI9TH1ggjLdWDA/lH5s7CpwOsyXVeD9V817UNUrQO/PJVv7NJJSBfBf18vvLUprfkH5+
UIfH221dK1eWYscXP4fcdtszyQK/ZE7MiEE3ho90Ye1GQhO1Wy+5WN5IWnvaEVYUK3+d8ugN+VTW
BobsvUasQsUKgBibGi9Qix31Q3jgpfz5TcnsxfIxr4AmIuN/89DGPGVQba325MNKu/QdwqBYgUNg
WvVwzW8Y3OnRli5WpRwpE2aYCGDRI90qedxw5hl+Qon5q2LwvfWITQagQgVVYNMNtOBKOmEbbpVh
nPkUb0zxRVsYQ8C7mYo3ICoDYUjUOjVJt4XaZegzRokdkp2Hi1listbANURBI1Drzyuun95bIR/x
Xdv5Yo9Zj5r0woAVU6lSQ7yzisByHdVsoO/yFYaaS5KeYxMTPbKZM82ybqUDOW7YBwiMxxEYs+9S
B00YQ66M+xwBDTq/5rIlQZvHEiznQKkep5/cklUruPUVqph+RAbPHLHycr+HAukaWk64IQzA4pZy
8MR+POJIXmorHOjrYtSxwtQbMXo+Q176ErDc3Y95hIJnKA9tbNEicux9kvJEUho4MNKkjTTqNINF
qp0nCYCOVE1SSsln2izlefvnAUaw74yVoByatH9PWOaxFFu2dRBOwmrtbjKiMw1CGZWrxrkl+OnN
cpEyu676mCwitEmyhBmCm8b4bsFJvh/kI9eTY/bxol3f5Y4tRw3ecLbU1gb3NV4ST1A0mZ1jCcPe
C52o6q6noMzB9hQfJH0DMuhdjQm2lYz3Vfz1/Cz4qTaYj3DpgYAWqk3knWarx3uMD1Sgjlr09vNq
uVcRcpFpW/O3HZnRDAV5NHVb4yONGJ/3QGRd/kRFEefQxFS4iEpIfwI/NUbqUmt5VzRwDLePajEd
DFXxIbAbAFd3FvM0dq/+SGGTzRqQsHqo7S373m1oZ+0C0lTkspdzqod3HCmmMNiVl1FOWEye900O
/EdPC1TfxU2D8NzAHCjKiV/GtJ9eiroaQKM8AdBuk49p0T/EHlOAPfJ3x9ygoALkS+q5kYFtXm1v
QdFMmcQ3Z/KsbbQCB0SeIf16Be86HCRkEPPXOTAqH8zWboi6nDSi83g3FA2SFalhNjtlItAF0QpI
Rbk4SrQZUEPhWh6t6R/WcAe7ekwIdWpSgnrH6LGzOeMZZ1v+fKp1cqdZw18cEAQBTZwBMlOf9sLw
Q0FSBxvhs8qh9X0j65QfVEhi4EtozCbzqYg4fGpkoCnqv7ux6A5H9Il0WLg9kRYHPtM0ERWzpBV6
MBnIsNwYtj+MSF8HU4HuxWvcqzH7J9xXc6taUfTHLl2VmS36gVLj7z9FqjliMP4YiKAebLhYAOeM
efFwbHk5Z1XC8qdIeoRMdhdLHEC902dpOgfarkbD0LCAiQ54C202Vj1M/VThCSG+q5oYfNdvOvE0
nogs9/uQfg5DabpPMLZ88o+7L+JWsHoa/jOkl7KiY5mg1oUPmyIQf1iTjclqQEOo+LQjsu52zUuK
ywMwb5XxI0mvIadM+UXUrlprFWmIZ2FttpUTSad74Ex4unESbxAs4HYJTWACLJ29GYNiu4vSdiYm
lNlPc8bUYKoWvgJEAJqnuJ5OtBu9ML4SFfIHsh3Hhqp8lUbD/kDvgH1a1xFRW+GKxMrbc2lur+tZ
2P83/OSWaRgnOqE8zApt5xh+mV55fJnw55bDO+RH4j6+/hbztWJxUzaFqAObYC73AF/tfO6ZUL4u
+xAL4ico90tMVzKtJdrPamnX+50bw1OPHOtUYmmjRTovVytLfHIyf04Z4QS8omajEpak2mZrQyTX
JvNc4omtPZFynfcFP7EZ0a7zmPs5ffuOghF1n6gjE/JV6h+mZ2gEJgNTVGXDlwrCYwreyXouiSdS
6qPyT1OFg2iJvmSbRCpj/uFrcoJGx0ehpFOf86ZavxJegs9jB7M13ZMwzFyC2guYqlDL3dwoyCoI
LUUKt+AQ8pSiGSdyfkZoBhqhZ6qYe46S7GDRuBUG72sqWDHg7PIE1NUX1efIOJnqEaD76rDtgF2b
PGjSHECHlCLJAzWU3kg1SHlwjNtyJkh1A3pz/TFyIaPKBCFrp5OzTaHG6ND3bPmWVPYIRWbWx1dU
UmLi7EYWYeT6ROKCSU4bMgjp69fbxxw9cgh0I4F6hsAURbaWfPDKLH1tuExriHa1HCJNg4yNg8C3
X2rCQUANRzKN3Xm8QDeYlQBfcNrG4CrIF6asg5u5KXCT9wOcbEKScxLed9ppEIelE7dxTUA/Sdi6
1qPjrS9LJlbhhTAmZzN+OygSGlEQhDDaPAva55Jy+ymopzwhpn27SzveWAMujST+pYBft3uR54c7
ogFonYSsWUvSkPaJXoWVb4Iz0wj/pXCcPElc8toRz4BrDc1Ur2zk6qF5RzhtIrPD9qgZyjrCN/oj
7HC2Lmd4NLdA58pAuchX312uBV2R+wGXRwXHMiJdPDIY/Jsog1GgajmrrxscRnPVl1vnLIlB0O53
CqQcVi/sYkxaL3u+TkI0VK89Ialr+i8LLhVNA8/MAMiYz+mTkakTOIcPS8hW+b4gt+r/qaE2MimA
HpON/m1muyAzO1iK94oQ0iHgriNjB6+mbIQgJ+mDwA70KZHdfFZMf/uoFncRXsPvGkbqIgkc6SgO
pXfu9TebpV48ZnAPVOnkETCpVsfWxoSgWJ5h2bMTugUIccDcccqjS7MXnYwXd0XonRbaccOaGTYZ
05GTkwrsMt/3p7pqe0G+4iRBOShBNVZcqepLhMEjRBhFhbyo4vpqpfYqmJUsslzLQAUe94DhXuBV
QaczvbivvrIuoEXs3p9Yx4IQNPcAZD0IQEcD5NUqsqFT+1yttqmE7XrFp1t7WYbkBXNKuKo8R6DG
36bn4m6AyHd6zI1usujQx3hRewpYf+hGt5tRlkQnqxQKNZrsJE5g10yewh5TqtgQ1zlvcRJfmQTY
29+JSm9TIXyn0Jkz7y3lpIvJSLOFav+S4lJq22gzK3adak+Bg2ye64tlCgNdLN5iqSjEhk/3Zm4g
xZc/CgoGaQ+ZzighkcA89a/zirzgLNZbFu2anHkp6xgaI6+neJotx4OzfOW5kqiuHxaHFopPg+zv
tZhdG+5x8z1n/p0fhHJI71FnEsrsPAfOw3HJ8Ag6cnHcYgad7X/h7IEoOVpp7gMFGqP0kfl6RYOJ
NXCkmCI13Jr7tkBx3SYE7VwNlRJf6rYsLuUn/f/fGpIz9aJ2bDAFoZ/kT5Hw9RV8CzT6gcoWAdD9
Mnka8UjD6lpP8rfWkPq565GgjSfVqLCkQKhmRyJab8+43VYpXPT0c9C0vsVXqBvrb88Vp+cZL+J/
jLc4eezlbPC4/BNWfmgYV6/6DaQyzG1aL0VrV9bPHxCYB/nPH+gngd7/atCuv3FsV2FWTJRHGZgS
tFL5KAWQnaG46D3DSpo+FcqrBm3y+//DzAZ6tfqY/QGNFeoXGA24Rk+OD5fFHC4BDTDnqqpDdLmU
/4QekvGa3m8LDd6eECZpHQAzr/DJWIuhyEyy/GWIZdxA67dPNg4Xrw9QFm+KLRTDWP8oD0Tj6kAK
xr0/oQzK0v6g3at6aF0O2X2lRlb5kcy0mwDIt6Ojk8nBEMzjlNLzn26lVoMigHd7TbhtcqTTf0Qy
CQ6BMPLvbqkn3n11UmXAJcWPO01penzAK2zc3ZjS2i6gROUwIFJ8YG9LMYKTC9DXgmVWuzxeglqd
JkbKP5KkOGTOTR1dqNpHKpyoDqePo85QMuRWkVYTXw2trXcXzVXsqTj0Z8crSnAkk8STCsTUQgwr
8ca4QDcsEBRMG/M0nnNVKIcl/EXA84yAiboCxK6pO0KKAwhGciwK4nnUiXtmfzqQwRxQfyR5+hNK
2mNsIrkDESJPTAt/+e1LpHiTZwxcSbi0njLLOfBdfUvNND35shY3LLhuX38htosG37lNy7UKWHJp
yvnC3+VfQ4zmbQo+dgoGdyNurwx2JjEvkt5N6jaVj1Xvtx7hnqEpZXCGvWD+zjKJVN/dtd/QfVZQ
VJbRStx+JnpWC3iQiInvOlRwJPZ9KxX/jYP73n4U+P+nJmorPPkys+P5JD+g1KZEHEX+RPgBc9Tm
GvaYEG19s+5pBEDtybglMaGNwv60+il1A5BUJum61Y4/IjokZ6xVRiwtaUvWp1uMvFW/QfpMzlo0
2tY+3q0iWUDAqax6f9GkO8zSYWnnUVdh39zsNWmwxgN/oBpF/KUdwZUBrqtcWMfsqANzaefx7spR
eo2A5rwSggiMATY7ogTbWdc3hXAPubnJM33ZedZGRFQUbFBENuty7m1+mvoG9mx2FSdNke+1IWUQ
8nufEh7Y28l2kbAQUG2jiDHsXwon40SVYXEbxgWGtTAKpfxjleoixwx7nWtPAT9k9EHJ6PBrm2m5
IlS2Q+hGXvtk7tkatDEAqrF7nE99XX2AN2LD9TUFEwpV+adkStBGQl6IaZbAPBFHEsdZELdBERfi
JEPLx28BnEmyNtMcs+SSaeVZeWXWnZ+2LCTfxRRpyiZudMgvEs6v5skyp8a2fwvzPCTDw0i2QZQU
K4lcDHzT5067vKw/NE0++1wJzk9CufotWKQehhFsVnRK23jQN+7FdccYAkobco6C5C9vaIUpQPSG
lHEEzTfvtzRtHt7tzgCExBRfbNRbi18dB4mVt2gkVkCCF9lg/CYMvY+bxyjle9PoMCQuI2y8pqls
lMbmRs4LSHftZ6WjB/IQ90TidLR1GF8/D7uP6h+XNe5auOkAHdlngF/CHMA+sr7a2q4KlDk1Etvs
wi2BLi/0p6lWjkndmyeVwybPWHZD9KaFkKvYruq1thUIPNOoREdtddzdwgHA2eetRITqt2TYuZW7
MYKDwAO2oNNqp8p3C/N0Aakntaqd1STUTT/dukla+w8pO7Qry1KUcXSmtf39CDZ5jOoy6jLjhcC8
kwhW8L0ZjD8QBUzEsIqdm62AE/+FsVvMt2jTBXNwp9fYOZNYvKAUO431xgipgboCuT0hi71LD9w5
EUh7ynuZpOruOMjIhA2PfhIkJPJgrXiCpdhLoYhUS3fZIEN3aQTb5h0NZ+iXNS2ERry6nGMK7oie
s0/k9qfaixECcM2Tah0FZviXcVLsYDURAIM75ZQh2C9BgIOBmxh8VoB1a7UmKCR5sfOsZSBMB+2k
A6RzP7/U7JravBb+6M14L9JhC1GKikSlH+Dni3oVY06Z9XisIzpzn2riMN4It14Lp3gjExrzNTqG
fRutyk14kZyJS68iEx3DCbFLIKYD1z35uei3KOVlBR/EpldvT40p6IUxkNnYQaCG+CnkcT/HdcV0
UeRXyRdlAeVK0SWxjYKgf0TE/mR7YUbjjvuv3VjPtUgwauys8NxTzc+vBlNwp5/qvzwWl5LeglV8
jZpRX2qVygfQpitj6b3hqgSJGF0hImLIsNHjFxPOMEu9JWkQ3P+XIHM9ZC7w/8OGVEFgdXxgs55G
3HDc7LkrXk9/jO0YB2zlFfLkZFL7JZ56+fMSlLvTCiAUPK/njoPjfsvV8yCFV7OAow/D+2RbMWd7
fF+iGzV7rDtPsSq4JgN4L/RQ5R3oVUaIB0iARFFwaK8FHyg9D6J1hPRlOto9fmE8TdbSNKTm1kbI
yBCd4TPB52sQTJwUgqu/7DKkdgU+gkr7G5ce/ee3eC1fyyt59XtqDTLtwsCMA6N5F+DiS+wT0X9i
Oi8+BICYsICPKFJz3/0Ca99yoUlGnXYKhC3TI/4vQCesSDCdHJz+R+l4BEDh+ASZ4eA8zd+QucsF
OkilCEqmUOm+Q/ZpT/g4bcuzD4+m/H19OM7gTm3Oixl4LRyfOXga+pHM9p9UGMSwg5mHJPYdsEVP
/J0uwS+xG3mmt9m7u/NPOAbXgGwvCf5IkOan5XfrbiV+yRj4LFZyr28phik9Wu1A2KqUJro71CH9
oS9OzfeGx13M4gZT7oM3/95a7suvwA3pq/zHkRq9ySCsdlF1fe++dHJ/J9Y+DPwZxVTa3VPtk1WZ
lFYgB52lL4ApYBcOkqL2p1KFYP6I8Mhu4nNvvmMExg2PXU0+6QOxnbs2mjC4uw6OirmtZLzFuG6q
LVn5aQcnou7MIHYICsw63PswAlYO3dzT4xQQ0jM4A18WfQ5KhWg/17zrxtLMGYzKhh1lLwi7kDbN
H6BrXmR4wFMf1M8cXr/mR+Oix7MByg5l3wt885zWCGkb8hYVNUzofpVEOOw3tLfSLN21tfU2++Ae
pzr6sx9r+WN4Rx1qOEsUXMrjXh48fk5HNPwMM4r+kANfwMaC+dHNIb7TLoRneNSNxVZxgrM1hmq0
Dl7ds9HBwoXRPWqnpIWIVYNmqsU84ribMFEdUKZ4mGjDaV784kE5ML6yE0Zad5ul9hoMSLFbmcTR
RcLBQzkkCbA5Z/Pbuezc1CxojJbmk4oVMWIP0nSAO9o25PEYvN9qcXboYO2CQYmofwZ5E3YGhMYo
oQEoUeEIVu/z0OH8x5dlSrsUCTFnimlzjqIXyyLI/hgZrHP7ZPBCI+PICWIlINQcDw4faQl6aIEG
TFT+ZGFtWXnrS1OYRS0qpzKe4APzcnzPyPnt5Q1HHTLaUZvAWReMWa0+1oUvBPYpL3McooM2PFaW
SqhlS4Nc9+SwRjMOe28WqXtHJwhHkW+Dpy3AL0eC22d783v+66GyaypD5ztd+C/LEP+nd81yblU7
iZ1eD6g2wA3MhMlFqbR6aqG5MfMMJ0yBmxz/lyHMTj2PHpey1gxUINto5GBElt0OO5snefaYvmEB
AhqQn35smgVKa/H2QqnLxWhNx5SUvf2LobCwZMhBmWfShJzEO+ko0Vt9naqx93IQoHbDmRJplL8o
F3VxISMjb/mZUwaaiRF9G3s/8FU26pc7varbgdnKRGnoD1jbQKp09nzL3djXJTNyJwLyXf6RoqCA
/zlLnvMn4urOtEegDh4zAt70pauOorTFQouo9nlROF8z20GoSTokyg/VPS17b5iyytqfnO0bdvJS
eR39YIo3MsNG/6FkXBpDIctzTHQW6tJFjrbqxIjzd25/urnF4pgZfHi/lJK+nuCt8On7j5U/177f
ynNbWQ76+x1fEEhfkrX21FMZYVM69cAZpxNkxAByjgSsaADXL12T3HNuZm3mVPDz91hT26dOb53s
kBRaBMqWncaXl6PHz9ILIJFCQICW639Q/lG7QCUEQ3SE04J4RnPdi3UpTp1GKz5dC6g6n8NdLrzH
hznjbuOIcSQsKsxK5jGGd7+ffI4q7A9ln9f5oYr65P4gucjZGbuzP1f6WX/lsT0AwowmWjAQoiUa
ckA94+UlqMplIMmEISK412/TvlHsovrN4yHMB2+IVDKp8MFpESUPJ1gHlgW0v22bQ1u2Ug4VKEq0
LKKtCe4Nif0yB1XIjisMSVQwRGVc9lkMfM9ezL8hcwOuIsDMVD8TRW36bHo3syKpL+424U+ml9cr
XOBilt1N4ovUmqqFEq16IUYfvS3eJbMg4jQ3Mu33g5QrVYxQD3LnPb+CF+oGF7jPsmliSLjMZ4fu
Aj4rRfT8X1+Pkdik3DaM6uqAFUaze9OpQldw2qjVluxT55Og0YhKieX8B28v9L7rpb6M23Yb79ud
7UPKeb6npkUlHPNvMvVHKat0jQ3VjfBE+FKb7Hbs7/oQTBgN1CrF/OGWqVrOkZDUCZjZCznV056N
lJrQjoFXMbz3rgSJxFoOivLSaWKmH63vn7TrhwYvByyb6cpaflbs+hrd6eG8bJCUUo079p0D/jFR
NgFn1VJNG7GPJGxJsugMwWLoD5tUfjEfytV8yoE78LjTM9+RA4m71mt66+UTTuStshItRH4n6yrr
hRRosT15HHqISC7Aq3ODd2/zmoF5bzsTcK9YSWY+IxuhZUllI28O3KIGctiktU7G9Y8hoMEjpJ+K
KQZqqo4E0AKV29MXlNYKDGRd1EsusiPlHvMdY83v2ArFRPH5G1r+aPfN3czK2TX84ZwwHHVuNDm1
2kRI1Syquv6ZsZ8pj/cueXvramQ0m04vWLIKhacgGfDUKhtvHu7H7VPsRfe+drVEBpuWur/g0nLf
UABAdCzJkQtCQSpcMXnbMg+qKWkK8YRy4UAfAgQkWFy6X9G4hKSlIGXU4PjzI8QvvwOlJ4bKy/HJ
WCyHd/Wsy/HlUjrKyjziVlVFhD96t5HVtC47xEjTqdp0chrvvYBd2tAnZ8jjAlMncG6l7bWtRod1
bcf9GKz4D/kNYlrjzWXQpF82BuO3BGdbdoO/nbrrNplFwB+HP6l6EwIwiDK0cDRO3xQqOsbOZoyD
YA+d+kLcp7buA7y+1Mb5ae2DLPvRsV4RwRjLvPC5wXJQCnoyIELd1cihIqFJjgjA3yLBboqyfM0P
hcuLkMYH+4I656mtCoCYj7dzUOuVm+ObXbBYSg1dlUKNtLN9xIYI7Dx5BBKip9mWNRBRNk7GqXTq
FvPuvAYXk0NBQge0xHGq2AVZxlU/sb0PHkX+jt+cW5IhLsN9YBV0ffojUl6myPycMEfzg5W2V97h
3P+/mbDsZfovfF4D8wRtQOxvkTDDP2yvuYu7EeGNPtDBEsDnjZNKf+gLgx73EdkvA2F0LhA5q1Ov
1d2+7kRI1zIWGT5RV2I48IWIZ9AkNvJOJpHhBPVWCiE8L0ptaxC71n65c3UTJd9yobwK0RoLjOE8
9b0CJZc2rtu/d7z6PmhdICEv3hKyRIPIK+Gk6RwCmQcwhruwm0Y4DfTR2yvaDDWtBnMBFtRRVVuI
+Sdik9V25PcMENxUkMswD29Qm8vfKiuXUs/VqR76b4k1EpCoyNSIAJydlWHTbMJrUIbZJ9/m1VDC
ybw+V4H7v8+2N9xdAeLDHd6bC+vnIu4E4C1x11HT7P0lTRhWftnhqqwPIMRvpr4k45TjlyzN23//
dgiVek7NMU3/ER5elzojcR7wFClD3uSA1E1ied7pudtdwLzwXPj6mUir4m9prneHNFcbpTR3MZWD
+FfWDx9/NzS2XrNpm5LSivrFwfZLmf1W1yyAhrKpqEJRvGu53K0ONfChHB4of1YB4KnHp9E/9GxP
epAhd52Q8fIloPyEjn642itNKMG1ypGbqZ6lAfDW53zWrzBQkRK0jmsvcYgImuQStHsAHaR2sXZ7
EthK/2MF82HNZPo2k/JpYD/5ORw23/EN1Q9v1RK8bc+cyQlqUvfjfvgy6w12RpC7XoKTiYjTK8mk
EP/hvVbLHBdQmWjLgehkoPavDTq7PDcXSAzTVwzDyG9CoRFRxKxoML3TU6aJYBFTTmsNA9OuXIrM
0b65f2I8Pskfg1nBiwRhNlgp/0fmamx5wHPUA9cR84vCKePN8YYrVa7e1wO3iyN8xqIQlyfUXZkV
7WxUbjZFrVL9unxVyhecih47T9oibkDnO/lFlKSFcO8+j9Yh35s9B2Cv6z9ymptssOkYqQZ46v/L
E8d4cXux8sDyVHkFUhJ+PtLOrE3LJJFAyakAVAW7OSFA+6XZ7ZeEXpYvO7rWYkjHfVbbazNRKGf2
q5hccxX5qzmPhJvju3SF00SOfY+luJlqw7GOdk01Cis2VjHhCwVHRFNClskJe7SMyExqKUYnLG+c
Lg/6+T/yGKjS5lJj5afE+pUunsPZtwiZf8q7JG3ARtsZVES80tHFBB9ZFkkYy/uwlTygoRRI7jl4
d1k3WTKTroxvLpBGrSxCOyyxAzUcDL1UOh7qzw5qdhhGS+rMFJc+EKQmd0Sux+mm2DufW/hbEbCn
UfDwIz3+RILrO+7yfHGCzmeYMfRO2UlepwVhbzRBXkrygw2sEFSMa0KZWvdSwtpv6WwrqsO57msY
HHhKcaowLQZW0OVgyAN/CPPL4jLz3kSjB4mxTe9Fm2PB2vqRcSMWnJfL71bDcp1v90aK3edQlYc5
f3BAgotizFHf3CfyxnHhx3vyI5gN+C/ZuWduv9V5RvPuUleTtbx/+ASWR0iDyUWsd5Cx6il9GolJ
1sNakDc3pqQ1f8mBL9069sK/POj90dA7aOc7J7xHl3yuF9UBBsoKWJCKpOWI9jpGn1FxpELe//+5
eYwIViuLdTa2Z62ycQsca9KdIoYVEEV3BetnV0wFF7c9D2X58Etdta1FTxyuozXSJ6nBVpDnD0C3
717YaX8pzuqUow4vR5UFHqdMIVWCPgTFRMJb3fXa6uHMeW+J2vEM3tfBdTsCsIfqUfzrPgxD2wd0
twtzT80pm6adeV3fx77LNJOpnsss2BENV2jfILQ3SZxkyy2ln5EYHqlDIyvGm+yKY97esYZrKP5o
gJg73IodBXgf6H90yjhSaMYoQobAcJy6bYAloqWICVQP/ldWfD9445JPGGNi+dcGHc71l3iqYPFY
f+tQyNWv5kPZBbAyCZKKSBfvZN0sdd/IQy1ciMCGSpALVjOoZd5i13WU8voSq1H0Ja1gHaeG++5F
hYZNcQ8Cpbs7zYcPfCkrEDwCNqDNx7UsMV4v31toiCdTMmcRjSTkv+rWdgsa9e83i2r+igPL+vMO
6p7qyBEI8neUav6Sg105AfsKe6ni0iIfkmNFM25EJFHIzo7d5fV8TGoSRgq9kRKKpPq6gOs/oN9j
UNQxfedeSwNrPSuihrdGkmPgVacHA7rfPwhwywEDwYRw95jat1u5KbjSfpPwD4Mav3DzTd9w1rZ3
hFHV14Ppzqjx/gKgzdNI8TIs/nopnIqLpYBb14ahxc1oKv/bUKj6mix4Ec9m2gx+lso1qhBLGVJl
lXc1osScy4QTxaSD3uwEdHbWcd0s6LJSOe5trMPorelprGNn24sYQi4dqiQ41sxatyzduHLGKf5z
khu3ufIIVJ0nkJrc1jp+sUM1HXveCafEslfnFuVYuY/HWOSLWJ1vpi+mc9Ha5ctqgZ/XPTur0rH9
Epc5QvGLaGX8JArOAMktaapjYQCRnUqhoEEgBLV0IupXGNPZXXgMAMrVBa1TpaW5at7pCy6UOCFh
gKvxUrEnzV1D1F8sIMD1+GBBcN1TL1UKQTE3s2OdYVFSHz5jTlp0AWIS6JoxGLtLmgCSDOFdqgfh
yBSSNy+dDWt9EuP/BkHd4MWzan1/AeU4I8/lCv49O98Ml5EaYuch7vQmr4wGXunkEumaNIerlg+m
pxfGw704/TYVHx64bOmpASRMB0g8pC56tjIDvKONOEet7W+8TsW59yRjVmmvjCi78Nm/1dRSe0OZ
WG/VDHm+gO7EJYqAtsEVxDrLDZRPwPbxMgC/uhB/mUjjdzFOoFDOoREJS+M4DpPDXdLvHFhPffdR
g5jHoClUByV4g8QBo901FBCO+KG32JO5Si/TKYtg5LmjZeALkkPL0NwnGmfMZ4qPc+1xA3su4Omt
5Nmxz3EXz8yyBUz7O78bJlWAsNqpUacAIGV8ZGe7KqTTbsusAyPG3mn/tFL3fZACKhyGz3JYHXs7
nHfpDH0AsUcPhp4HZqEoAFz67mtIOzmbrirSnRO208ozLdgSmR7I+CDMZt3n16YtrvTO/sG4FSnQ
2ftsivRBWLXo/iWWA1JeIT0+Cqi/tMyybkyjo5qUEkJmKzz5QDfm0jnDrrAZkDgGYlOvaAl5x9sy
XDEF//vN5gFg5evGKk/bnGoBU+XeXxhXtNwTioMtO4ji8qklbDlSeX9DPBWZmOkqgN7ZS56L4tXw
9YuNH9GKwxuSKPQkET8OqZPdYu7bkric0dxLU4xWd7sxT3XpJk5apmHJHySFLkAykmGEJLmDBuZ8
Yrx/C9Ttn/EF9oI+tDUmCdCpzAJCYmHXIssUYFlJ0bYmugeogB7pmXryrOLBAgVHmp5p0uUdYdzZ
to+Ryf8DOD83aUc7qLymEIBdH1WUO7+SemROBndfmSYJ2ZpdAiCUaZHrKdqfUo32UX+cYz3qX8IP
xpVuO+vp2OZ8p5w+pidu2zjGcv5szHeLa9mQSgor9dcPnWQE66B2+tDUnp8Ol8JESd399aKw3ahm
fC+HK1vA4YSikq255Hw6qgWBJw281goND3zEhwzOS48thKjEuDIyK8VMp2VaAFq7DyIfvC0jWXou
PdOYNP8SbElq/P5upmv2Y3rj2MsjEY28voZX1e2l3DSMXHOxZ5mwU6l6UFUlxCnAHZ4pGMsEIoKC
DwkMq9u7mlRj46lxmjDFRn8kP1nhnbWLKRKeQBjSx9spsJNV+/9m0F3t1Jb2xjzh9RDsijJOS0WT
Snm4IGqyAtRZp2eY1XY4uyNtvH2L61TMSXUiuKVVDxbc2IIvUk8/wZXHjJPkcGLbfbUjkPO/gcNU
s/CvP9F/hDWwVnTi5xcAQ7kV0NvspNWR42yFrqAoMs2QM9RFYtOypBz0LQk+Ca35/RyxmJjqkcN1
KrKUiVCLRn6fUapkbplyF0vxGCzw99QVmov9CMlrTskRuqSk76GgHmQF5V7Lb5qiuJZNEzWlcsp/
LFe+oZ+5BuanafdcEfyHZw5z9oEqYA1LD4AdIySXW/6jWYYUfnY6KeDewgWN2ezbNS3HtyJB8teR
uTWbs0s77XrTuoFrmZpolIv3LWQRfmuZqxdwgH+GF08SEltgMaQ2LwqovrigDow/mtNOc1yWW0NM
Cyy8tkSFkyQY4C5oQk/OgXYXodxHD0N6OHq7l6Seg3XhzKOsn2/0DBlFWdUV8NUGDbBB+A/W4Lv7
Otzux5wgVXao/wnL5Tv+lZ+HPweoxHaEAzN/7KMvnOpCh2l52DRX2m/ZhN6kX0hyZeSr40Ue+ipq
lTdaVx463hk4emW3nTYCzNXDgZCbec2i2AYr7kzeFJKXbLXlUfqeV+rKf15o1ppYpqJSXhsRW8dG
9UickNyi+Yyy4eDSz3rDGQVkdKrmBetiQmkH4SyT6Pk6MQTFrGnnY9cd+H7BcZcJ/btp5XctUToX
I/g/Lg7epQPoIAkJNuw6fBN42D/iUgQ4qqFtLhHqow9AbbIP1mvaK80aSnnHOomfMgebzwkd5Scs
f+lnhJKh2Uok3SleVmfLCwsWBch3KYnSf5tEkI788qryUGcFpLE7LKIYn7uur9msJa9tcHTMTUXZ
zUEtryo8AtH1qNakEc3iRvMfQs1A0MNBs9s74gmXhv0e8B691LY9kefCN9CYqsoxGxHOsKXFQqxh
TLFqLc86diEhV4wom3Y73nOtDBMNGqvV7NTb/87M3SkfaTliuS6Ls+zVQp9SYmN65i7sXOnRzdpo
T5Q7zdBhPjfuw22OUxyBpJapdQsmulw39EW+V+Y78qQWjZ781SdNNE/wo/Sl0Xng+bajAINVdYTy
f2d0RrM4mc5bkaUMCNDaTu0mYByQBHFDq+hOn6w6X+Ib1jTEq9O8FkH8Lq1Xd5HKdYuOf37k2GzH
oLOBXdQv0HsaMHll/P6Ux4kJYh5kxyRefHG/BRYYHYf5urbM+nDFxmUp7kmXmd2zox+fe/jQ/dKb
MRgVsT+TjL2qbK6Z00+vq+MIYd8utiVtSB1zcCkSWrnxRZpkgAZ8SZBIO8Ox1ijRAzCmVroxHwvw
gh1n/2y8NTAJJFuO409g7Xc6ihOGFZ80x6bNccH8ucQZYD/Fu2A16ObpUcbTgBwAlnZ8xKiFOn+o
pflvcC14OQQdTFV+x5rFTak2USSG6MrBB1UpapE/txS34MIz/cTcr+EhaK68ArJdZgP9jOHyUCoX
YMGbk3jFDYivvtEgqKyp9CYpG57j/Z5B/f1pRpftq+OPmwwER5V4sPJ4zAKmKoDw5D8CSmUW11RT
l/dCdZ+6+iESarMl/rTQGc2nDq2OCyLFMMED3dSkeXi1ooEKWzTANHFP7YN27R0MnOClpoBNqLy3
iqPdNNeUyIa5G1NBKbIJOENlAk2PnL+lCGn6VTIFYzhCFFVP1xqm0N/H1s6KN8OMtoiBcmURX7V2
aO9zgezMXHAQhHy6INmmITLl8fzT0vgqzVqqAU4pIK6fHyWywfSwVmCGG9fFC2Eb7u+oEsp/abr8
+vgYri3u7mGgPe1U/Nrc3SGKwqvSlOVFUQnhiE1pIied8XJKq5dZw4AL4yAo4pduxW4tQzTbyrQy
1wt/MSUvCOWKg2LsvX/oWwSnmMjlktxYsbTjOA8kxjtqHiLt1IFVmlCynS4WzT5Wo3YX7mhKazxY
ilq/W3SEe2YHBzmR6fjNr6swDa/ypKCgFqpm/rwHb0zao4eCwr67NsVj2m0DtK8GmIcKFKZfUydm
7Nyt8CZD+EvOLfw+gZbH0km8qwjyqR/oEqKDPlXLJ2FyQ7QsOs+kDAb1eeA1lL2MHMrxowhjiQ5u
+0e7cETfyxwaNxxPpgNB3qPnN3m6KGEmc7+uHTjkjl1NIj5+5tlUA2dStrgbkzO9HmLaYtGsx4Vi
VdHIf58sZlWVqxgtoUTI9qPsgJ89edijZlHhIaOB5dxS+lwMDk1k4gfh8fNHmiJiJDrvTgjeHkxn
Q6AqelN5staqmt3vc1xbJtnIsa9ZvU1fPBcwqANlj8zmUZQamk+JUbFKX7KUVeBcxe8hup6GAdD7
HzDQBwsuByBvZ43jNhARDYQ1mBEs9vKv0VnmPxiz7ljXVBbxZnK5ZYGRixzYm6WMyKGX7JAv0cJk
uv6Y8IQiUMJs4w18V2SZfDv4vS6Q7u4iy8IIUKY+SoZDO/2x35fs2wdDlvqz1Um8xi3g5A9G1Ppk
uEAKeJAM7qxRbFrrDSBpb6wTsqmV91n+zsCGXCZDtt5ELLEPn3+dRz3TO6EqOtiDbqO8yTeI/NWP
Kdz9GDfEbcWEui4n7jqv5XoT5/EO5ydDtccraMGr6YGte083A7zY3xZ49+aT02+Fj+3bYVevK0ca
VJC4Ligbfv28fAN8pg+VHDtAT1G286aomLyvmfwdXPZkbU2HmHfVNn9U3ELXObvguqXDCHhn+KfR
arg/f9HlyiNJCqIbE/EUOSU4OFtS83qbopP6n6MNl87A62yEZAkLBg+JK2gjZGhVriZQ2niErNJ+
zWxi8CI4qgaKb5Rx1nHSd6atURrIARte4kVF3qWVt9XeOIugdi6xx322VzgQtOBUCDhegmEha04+
DnEweKqzvVP5OsVYFhoh7NGq7krd25+4vHH9+e/8XGQu7oqUjLB28jZFrFzcD4BEPpihkaPvE/hk
OrN05+1UdvbfVNZ/i23CgW9hEDG4C/qhKycUPOXRGNky8Gh24H89+Y0/T0FLTxre8zHxeOmHjMxW
va8GL+mEezm58iyLLD/tDlVmkIdKzPBg7KsaG4I+u8efWgW/2yDD31Yde1EKrpPETn+xKK7u2kZq
tYca2XZXKHNUXo67dGHmy8u2LWO114Vhrs7mBBuKye4ICav4V2Oi/gAhD/NZdf5ofXMXy0kn6fSS
ePD2pGY+Tf9Jwo3Qrv6od0GJe4Y7HAmyu9pqgoq4VRUYvuUphwcc2CJd3Ps0U4DNnqg63/36lmwd
NS4R8S6ffxDvW+XusijA6NkPZsS+5VllZwljK3Xq1S6ztb1bs2tNTRe2pecIkQZlH3Vb1aSG5hj5
M+574p2JADAWb7oUuG3VvTArc4YFVJFsN9tTOvdS/U3R2eldL7ymnGy5yfJVc2k/76V9ZaBpdT9T
o+RJ8f1jX4Xinjjx4npHvMAXGXiSsYB4vopaZ3iRIcUbMlOgedBnFJAeCcea1QkiXN45iR6NLGR3
r9+kav6EeDtPXdC7lNEy81W+Xrtf30NoPiRnJ4y3/op7ul9VdG1noR7NVdTaE67nH+1aOr53A7tG
2pcjzThEwVffhwB2seCCSAVLlVIcZt62qzR2c/giv0ePE/hHsv5qgEB9S7FXvxJcOzUmqldMjl+P
OxiQTo73PFYvV5V7Le3SkagnFDSXYz9ci0jOppbph+WcvD8KoFnCAl6QLtIJK/YYm6d/olVGiyR+
cWjsND+/mMez8uSsuii9MBhOAinhtdpto0OwwigcGs/Mycmtp3Sq0U+EmzH9O2mcGVp3hjzd0xYg
SM1l1JGNxgKkeN8urxvTb505Hs9zr36m9cdI5RTXcBAZn3H+bUJRa8yzfFVKjRIomjm/pP0Z+Iyn
rRkBLfnS4UYcSPIjR8yyxUV5EbG5UPf7lGaa7y4sdaqFHQcEuLy8+XMg9IT4FThtqPTJUn7Hx4+m
dCbSv/JDOlGOyc+yrQFqprwYmUyapRujIfQmvbNUARVBNDeEu2pmg7bU2qsESgfvRC2xBGmVyyXg
hdzuCYjEoIw1qPN3FH+oY838C5QjHMkq6z3FIj5LzofbU7wFIisFPYZHl9/FQnUHQ7NT5GE6NR3z
GgyDQwT6/m/BNS/Pn+BQ75NxuCy5AP/UYd+QZFjEcYRFmdWXw2+js+WCsLCA773hGrjvitMIJe3m
F8QDOmUyPA6UdSgxCpl3CpsZqsClGWLyuSPDYAVpKoYx76TbqOw9XUJaElFgd91LaUQ8TIRq706b
x+caS8Ns/WpK0ABklo223Tb1xZGOCH1FGvzMe4ZHQ03KdbKzClJeDeVvtVf2Mk/DzBrRRMmUavA/
p8LQ/knGModni7F5i59Ki6UUIvDYqHqyteBqnXDmmNbw5/iXs4fspbM/GpzeICsU6Evs2xS7cANF
BoaH1YKPET9ixTPnaoaKWLxO8uHmd4yYY3qKquCTx4gWAv2qD1wyAIHGOvZY8tDe+lkCbrGUdlqP
YrfHt6c43kcMM6wVC0VXH3rsMytaN35hNrn9GvKpgb+o4HhO1kWzWzQBLV7RY1vIVCNz7BANPR5p
iIzHDNJa8CQ4i8UUFm8GOEns3iTCRmzH0S50LZnCeOr7XcTi1wu+4kBnQg4m8mVdLhrYKCgSlKy/
DSF2phByAl/uwURzkHlTN99JSfHrY96FOkILNY8k7+Z0KrGoEtdCPBmAJFvJjAiHkefYB7UXpNyE
DioK3szJO3JKawsPa1ULvkkrXSK1cLlhsnm2ix0aLenmglwBFPCojFssGvLdYt8xdjKkIzzpsIzI
Ag2s/nO+lvPYIJ+FJtw0v151ZcV+j5FjOurA3cqeVwQGBaizTB0detGKurZEK93ylUBpfQJm4aHt
V4G63NioK4bmRHRr4bXDGu7tBpFoQ3HEMrZzdWbnDR6Wr593HyiHHKatv1Rf3+4/HNRdB34XNrTK
KNw9tb2d67ogSOorKSy+5ejzQCo/qJmo+AkJQENCMOWPp6FGims9J/nI/Qv53GHEQZiTpxn2ICEy
VhYqLUqz07WG9DD5EDyZSZhdntkJOUB3i4T9XenRpI4rcCb0QH9FfcgdGIbHW0ugfZopKECH0BC2
YSOPwKEWfOLi9JDM6pggE9hkuPo9WNjjRlRS57MbgmdglNR7u/gYQw9QzMaQrdvPRK+aAsNFX7JC
IVacnKKKl/ObJJSokto1OOSloAZb45BRqKSjtYbHUxUjfp/bo9/HtdfQ48UYi8VTqRVJwWr8MPcK
ANOveBPzbawy87v7sp7snco8BIZWzwCKgYKzHNeIvo0fH/CGJaLxs+9c6BGAlFcpi0VhP7FqZV7C
R8BCK0eOmuzreiqNgYesKsHiBr7igCU0Ot6A0XPu8FEw+/4I+S62YnyvykbVmwtmFgeqU31jX4LQ
BOQjni3dQZiLW+d2HNHsCAlmCK5M8LgfKeE+e0ILL5AvAXwvRRUNrIW230M4L5QnPGKNPGUFnaFn
1cKki9Gg8Hj/ro0GFm/+knMIWyiPg2J6t/VfRlivVNn0p5AEwy39y/XE1S01BGz6g+hHDVWsFj+h
ZrcCvHVxUvWp/HqJBOZxacvOBE/1jGnqTZTvpZyEiDr0kM6xlCRBNiQFXnbsNPm1zJttXkcbZgRE
y78uWbT53juQPO437/+00HluVJC0AbvuCIT+ZBVC+5ikY/Yv3+Wpm3u1PLFvK/TI8BnUoOf6BLC0
3vOg7A9E3xsndaj2HlwI9Fg3O3C0kxYmlIFH+zBmOkrWNf6NrljA3fJQG98/ZR3CBXOMRtYz4jt8
kpv/DIvfCgbc4Zx3G65U3cHkbCV6XWLxz4JfYKP3MNRMzkOeApLYYMSiiHaXu+guOdXq2iQVPLx3
igkf6kKD2tdOgeHVtymUJB+XDP4F/MMEgZs4JyQtcGj+qNz2R4bA5RNh/AdqJ8LogMzSNbSHSfYy
5RbiDJrN7M9bGDfxJuuXJEcjNJ4v3XWItYMt3JruXXyEgkfLDzn9jaJZH1CwyMjFxcDzAt3RbQIe
UQQY1T6hdxOLaDRdPou99BCZ5KtCnaUDkvSKFJml1uJzw8wj2iDAn2DG78c1uvCj1+5ejYALT9og
v/7feYOXVVuAsktUTN9OwSuhVSvmx5wdTuIhDSqqcjJc5gCVJeKUV3FJ07r0L6JFqLQ6DjXyqLSJ
XJfrRSRddrnJmhog4XA+BaFC5jAH3ULxi8sAkzMxSBUv9i+O3zznx+B+Oexv1epxEfPVcv3+JRrF
w/D4sOWdrIUofVGEoh57UCVb6g6rWsu2lOgBq/TDipU9XplIQ6gBi2JXBdKzGZWrh9IPJdMMXpLA
bub55Y1wTbhDUhu93VS3vCg02xpEvFYThWRDqV6fbD8kOYWuGCAtspdak6LUDyhHpfixVhHZeDDM
4m2mwznz6+NsFVjuJq8OelLZtmGgtozxcaFvhDd7NhsBAAvp5pG+6nP7tqUx4h4tIyjcxB/PQvYG
ybBmo1o7u8DiNGBLMT5ytSAwWVKdLIFCMc7u2vfF+GZSAUSYLu/mSsrrqzAtChDCoUnJJfEEnJsa
YCPbsr+Td97KjlfBRMhos6pTFKV5CRJO1ioXbKeJx+Wp5fH6LWo9gfwpHElmkOMmoaGKsnyVX9d9
Ml2edycwYFrERlygab4ZeJF64rQ9esEbDceZqY9tltZ2va7FM+rda0aiHzgb8VFThAUUL4GGYzxO
RhgYyFpJLndRtbdUj9d18hmO9PO//d7iz7ikbVzlg4XyWb28yn5SsnobD8KcoXPGedU3Ov1HQr89
juegfHs8+e61q/+RQcHFzQRs+eLouYsuIIYLreTgbzvSTPPx5AfTKGT8PgPg32ZAVmr3qihYyqiI
fUOk5rNwiHEGugczf9Ka65A0PR87TdhSJ+MBryDiFOMYTMbRLhYTYh17jfJtApUEkvV4r6Vj4m4V
E4dn1npJ7O4GbqTREYxtdT4QLmNSreg1Jppf9l4W+628v8PB/Lheakex1YZy16YjxiP5DkGyaaLd
iSO7+7eENZSSLdYt6YT5Eg6y+Anlw6scAGYsx60CvlNTz8mevf8GvmgnxHd54RqYLfxQxyfIHRAd
jo0pXqpEp7d61TbmeKIZ6gsJJDwXoVoiB0aE2mssAyQmzfZ39Lr1CckT4Qwe7VNnamtKLu20dysg
QC/8r6KuWi0OsYOJuY94mtYE0SKmwZS5sExJS5ByH9T/1cNOB+Q/mQa7uDCHx63BmtgSHRcZoqFz
Grmx3pAmOQp5ohZkj+NMMd5q1UNXd2RMhCnOhQhFbUjscuri+EKDZyxmfX0kmKJrP733ElDE7/d/
prJZvYUAAdJ3wo9lllNSvIr5g/RU22qSquEY/YltScVeZZdMGaZrRm4zXRbLUoi36jgwQNreog4U
jBvhX+cEFmQE2xsIe96oI5TPQ9x3oSNtyS+tcAlR8esMbRcA5l9hmKdXLExesIYewPuug16ut93O
JIfISvvk8Pf8X3ND8ksl67CkFf1WX/3wLi/y7IGiQs9UHBr/gRHzIa6aBDq3v28hCm0VpZQtkjeX
NAU/4EEW62KSALo59tVR774P1rVKhLZHWzqUrt17ReD0+pyRgfYVgWPPKw70cmsaUC6MiI96fdoa
ARuExuDmd8fOGaxVEAhkbi/QaY9999DAI7fpPsc1qMdbGTuHRU46zNEZwrtX6ht2362Jf0xktYoM
spKgljbWWJz0XYG5stSNlFn4jze5dYCQdZo/+C6zMuXte9klEbhxJ3tQJzqoiX23z1bR+yctukXx
eu3eqoPGyHXMEYzAKO26sAoLGuEice+PuojrzICsAmX2XErJkJbYCQ4J8Vz+pp18wI8jTXVZ17Ni
h2tYYDmz8gcG9b+VUaJqpIumLinvHl8lx39hPUrQejvfplt5zNrQvIBfGedCDV5hzdaT7M567RlD
lpIqGcXiZc/ZaRzdJCKoymYMa9c2RnlQF6Lq0TcEGj1IBdh32F5D8+tURK5+Vi6scwKyEguHr9b+
KvS6NFpHO8KhjLnPnnE+rxDzmXnNmZ2JSVknXczb58wYIMCj4KcRDToqkLFRbmRry/8yppTj44Ig
lr6WxPvuWSsza3Q+2kSkbnyokrJUjMyYLzlOkpYbgXGaoRcb9qY8E71mXZJNho8EpUWgZQO0hRjd
9uhbjk9ArsOttI+yrumW00Mip5KCHU80av4Es9eLvg5EUkVp8D9JUA7pC7pRRYKedempA8ETHyfq
akEDrKtMk8js/0SKfz2/HfLKLKOT1lVr7+VbReQjZdS69Osl87Luo6DO8KgZ8HLKdVEEUOJrEIv5
itn4rpwjyDs96lQlQSvI3GEisimFZm29npXyeAQLYWoc0uiht1jf8q378T0caHLpoPb6YddKQHH8
YSOomwDLiqbZKMNX4aMWXaWM7Ris2NeQOCiEVJyER6rOq1wLsiz1H2Xc7XZoWYKLM8R1d8qRAXrq
2qfULPDX1bWZQ0lIi+vFcRI55clDva5TigQwYvJ7XR3KSLluw6gv+jElV2a7ajc+xAbD9Kyr5udd
rOOb7gvgRjeSgtjwPi6v+zrLppu3JIrwGRWuIWUgiNaKecxvn5NAMvtfese85Zuh/XnyUWBzkYv1
EAehLJZptnpy7xD0GEBtnqzhC5vLnzyfdXM8WRcAOWpQQMXkrF9gjrpQWH+P827zs2dTYNWmEYdc
7lQ09M5iGGaBq60MrhgUl0GLqWQ8JG4KkSUVUNUCeVTN/jr5L1Smad7ID8eFnzlVLCY2JOh+lWM5
nbBzxrR7aiIIeJCfno/hGKNw/+axIMuYD6Dud1WyzB8/txLRz9Uj2dCx0mUlft/t5SI4Q0m1J8W3
hESdc9Bb5PugkFx417wDRLqQxzoXWE17dTwfIQ5eEdHiz7MBflyCECLXhmiHdUZcPaGyNFNYuLhk
3zXgbX0bM4ps95OuCftijs8OR8OVk8izppmvMSZu3OYUTEC+tvWqNer34kJutahaoLxuqgrAWDJf
oCKEen1ZtsUSqktwflpncs4k/R9gwTi6ExRiFhsKNIogQZahcl4hezDKXOXJfIMUE67Kqod12dpk
eyHBivhD/RK8re27ll0p+vVMtXDYuw16NLgJAi8EfNS/OlSHOYFZAbb7qNRswHO4qibgNPiVjsxk
j/AGMLfthyELw8xoodncWxRbzAiecpOk9AWJJKDo6Z+YgVG44HewFAiVw7tdhAuEi6t2q9DVZ64x
gQOWsKJ8war2txkvzeXft37zAt3PfiGIeKvD3okqidBieF1/BVf6NU83bjV95d151MzgFqo0uhJh
7TKv0aREtfxiVIpUFK3gUhq70zCa7ULyyVskIJr6fNnOSZ5xLeMEC1GFFwGOuwMAa23AtTG/7ytj
Nr8E5I7XG+F6wGkOwQZdNAMRokxGp22iDcdyMbHpOyolJvN3rlsR9Wp+k4szKOZOvkDfIHqqITbH
S62XpULrgoaRI8UewYM7Lo47jD2zDhyAeUMc7/715WEHD5Gabk2PeKA2y04AmOp1c6Dv5vPyA/S1
okuxFKkp913coDVDw8BRCQ6YI6EmyBKD5lN5oYOT+S/fp+W/5dh3pdlapmRdUr+2a7qMQ1zJr1D9
ZvkuisTxkroc24VoqLtoi6Emdcg6f+LhnmMdALEZ7g145MyuCZfF3qeoATmEOoH4mbeQOAzbFSvu
qJ6raqSBncMQABaRKRAqRehHzvPFnqIMeAacpwjuBmetKhwyQvoQo5q9Mk7HcgSK5ZQ5X9yxTHkR
x9PLGHrT6xVkOm8ILe6cCA+7TRtZqA1PyL5zdVZDVHpAHoqb4B2ouOvaPtPjkWoAi629pGSV+VXe
HTcdhCacAiItkuJ7BQeGFkCo76AODbNcBaNMBJCUMBvUyjyZf9yc0+nucbrGf9DZHmEWNvzNJXKV
8E5uZ6jNfpWz/AmKwC85DMOJ8jXCf9sYKxFVl60SZL59XgeABj2ECZiu9EPJOUKh0T9jmeiaw4V/
7XIEk34fBwEeCA7LfL6Vdj5hf3oa2q1083jV+9llENr4VpT4iPZ6xlgkxWL+tIeTB2FZdskZRZaF
0ZJUIN5/ro0c1ltFSldd2nEaabMXKFiVnoXaNNilVJXktDHIHyflJKVxwVleY7rIVKtDpOOq+M32
S2zCHH6BnARm2YmB/DXMPL0ILmNpyhhef0XA/CrQ9CE5h882KbhlYF8M55O6X2NwRe7rX3+cDwRH
dPdH8iTeE/X1DpRcFwNFxDA9psBKFkP4AY0Gd4i5WM18Dn1JYSUrmZY1fLPS34DbwYhUUC/T8U0A
WSwTzsZSCnnAbWe4Nv52mZTJ9CMJtb4T1dpD9Q7whqCxlWmZCNBzJsPKa+/E76WsQNxxA3XWviwI
oz2k4sqpWF3GhTmZDcVTWXuxvFzaFdliIalnLE1Z8TIGRryUD2SoZhTL9mrB8uK7gR+NLdCGPQzl
dOz9ZR5gJ5hvb3M+hbJ9UIQqByHTTNdA0NplsZx99zvS1OY3XD18ZQHRlrR1AwVmfdMu7ghHwIdm
sUadaiCdwKhLL9ZN2SGuPzEi28DM7WejZ0QugHrNnimk8xQ2jL1YgBHd8mTYEXlV9iVq+MqCVYFg
i8v+8iYk1fFSVxl1Hp5H9q9fkW1ICt5/b8EV8CVbpSsaB5wm2/q0AczX7BscCFxQ4x/Id0A4iYPy
OEwdEndoZ/Jgt5846L8aNYxAvvJhfQCHi7yXvNoDfpc0ctUGCyY8lvZ6hsOl+PovnCeJaDjVwTrc
lFASSI+tComftDChDG8LZIcuBh/jCB1/vp7bbOyQvOXpJh1H9nYIN2qKLTlRQrJ/cz9VDBjh5g7l
MG6nif/OcUwvlUPx3NCYRpiQ7LDvXXljMMkkjszSvNmEFHEfXs2TIJSLjidi1p/OGR2XfLw9ovFT
0GtagGycjpGkzOig0vTXzbn5QYl7KL1wexsUPKkryKoo8aywo88l631WVAIaxeYqsUQfRNPl1LOM
ZAPHBYCpDm1i5lNDaCb2PPxqwq6Wa+HEe/FeIZd4f7QvKyM9t6KrTVJmagmi0HdwaxZb3mWfMFIE
adcrzBlELbjb/3pp4x1a7yNGpdkLA5qYrkujTlpMUkl+YkQ01narxCCqWaVP9U+bhJwTWRIwe42b
0wm+G2tDW7vWLmZforpCs5TvctgL7IUfVMIPKT/7Sz65sZxrq+LdnpgUr6QfyV07coWHhsSBTMux
r/DszJunThnPPwYWLZFlGpqR8Ur4Yy+7U3nFrHssm7EoDGqfeV2+ehAcFliNZiqPSLYdsD9lzziG
yIFcqVKKUh1JNF3gh59Dro8Qma04z9k1ckhZfLYmzSOGjevuxMGTqic0+2FYpaK6y/MC3idVsWmU
+uzg73WATnVbj+vZKKBFLR0rkMF99VNelZtqNW9pRxircfp7DML+9xhQJPW+La28gH5U4u8+ufOy
8ad1rauPA8hIY0hIKbrhlzE7py/tJ9P3EL0hlra/Gn30t/MP0SaB/6+4pkhd7HDNOjPm5ffxNDk6
/Dt4UhYSVIvgpoXRkSB3Yl0ktdplzbdqo1ucscAuUhP74qlZZcUrGBcz3E2gCrBEp/GkWZFrl1et
G3jcVabqXb4QEnTWCXODaE1IPRv6IqwumXacV9xX1QfXbv5HcaTCwqm6wDhxKSacSZ+j5er3JvYI
VVNN/L8QI855Gn8/D1uVDcLLOJfqMYzXPbhNR12beT80iKiugcqCjH9yFYTMvEjrDCPCSRTWmE2W
o0qXx6mRb5BFHZAxCZ/0oXiNZ020Bjf2LtF5JdLR169tmcHJCULtMSDP8Qp5AAH1Ghb1/v6h+t4i
yf1eT8wgW9HpTtu/6C+fZBxWG2iaEqwxgfFAWpzsLDCQRBQPbjfCOGabwU1sBW57S8zDNdT4s7g4
w4DauWNm3TU66VLT+oOjqRfCGiEofpI3uIIzemIWrSH9nSm9kvSRD2E9CxVxnsybGfcooSpXxwfP
9b6sCUy72lXktjbS/F9XRhv2vIHb5OW6duzgNQHVmcj2adaTceqULM+6DnCwU4pRSjtQgCCFTURI
5H/z52aGCmQ7WYBUDVwLJM5lMvAxACrrnFqJvTkxd083OgUHlnyVI/AZCsdsmsMWLB40EUrdexIl
WRTnUJauI0VhUomKvH4kyg5Z2sFv5uAty+pwgGq1FTr+epaOQwDSzXWTm5VTAKqPVhcobVs1O8mb
DoqpLArJ61D/UqOSJPC+0gvV8Te+Z0QikXUdyxeiubQLsapDkO9T+eLXJRU/8PeardbGHqd4MCje
Uw3BGxmsysPL4+4UR9XoEiHjWtegDyFNiMnsWrxiaNbTcNDF/mN/1dhQggLJI4VuKyv2J3TvlspB
mEi+lvJ5ZCHnAfVFOiMIZL7D0iej0ZseoMEbP17STqLCQH64S00c+GCzEheSHOrDa9/82yDlR/Tt
U9GNvpCkS1HzMvtQFWMwAX0moOYKrCNyGSwf5/lCB3faVITFZsfX9VJoOc1o/xQaZSK35qjQ3es0
iJ+3/KjoURdeDY7chvrNO8c3OkTdhLXlXJQU04NISx7KJUmoF+36Z1L5LUJT3VoYgyaunbaovWNu
cjmn12Vi63YxB8dNKJSQY7HsMzZk9x9TX2vu1RwOCC72F2AX1h4BiG8d/6Q21J5W0QvbOYIEsTsD
nW69c/GpXsQVQYHIM8cj2kOPJGEbGi9f/gBlpZfaiRLHNdBscyKebPcfrrNRzu6ytZRCBFLvwJlV
N92g5rwH7r38KuIszkJn+hiBQ9ybGJz+aNou2mTKs+sprcTVF1vjUW0hrST2nlr8ssAzr/W4XmUo
CeF1Af441VRQwxq7JyZ++s2UmVmMzzXECeGzTQ40odJ4Tpi18M5fG+Tdoat7J8x60ZJ/FuMXyhLY
4/CkXK8KPFhWGGiPcLK+fqrnrjYSrMw+uxJKafXGdYOvkxGTkHRdk3Ntdj9yHkIMQMX8oUPaJXo1
CeAigJSFjlc05DrEUH+qEHl91MWucF2XUzbh+QbD/JxuMyhFLqOIg7qa5+jL84ojRlqx7FW/9Dwv
QaOOWtS8gwqXPlctJknbclsiSv6wueovn/la2WRT5qgvkt2JXJCQRowILt1OUjUF6mY6RIUAWnX7
7wMEghy/WsllBDk9cR7QKuR5lO1YMr9/wo2ebbnKKJpjk4VT7LBEkaS9ZbJuvzJAz26MkpQ7Or3X
syD1Wi20MUo5JBaAnzkcn6LdsqAXb1Fh7YU28Fv+XqsRW/T9WNXgsSlCVSMa0tmtnibkSmLJ6kLN
M4JB5M8DFv1dJzKFkupNgGdq6roSS+46eJ4sENiOSYbTDGwd6V/cdurf6mLXxJwMfCt+QEaKSu9l
/1V48gNaSyQIoe0OITTbfzgXkAhfRnccSINLhrQFIbczk/UIZp1+B/9tEh2to4CP+0KhubdCt8FY
sfPHwaB9ac5wk4jBvzqkz3MFmjpvpQZ4pBumaSYsy0B8hLSttbD3qDtHetjrv/o7NcEzGxqK/NGj
ZDJDJYpjhfhyMUyHo9a+b+5DK/QQbulHz4NtV26AkZemkLq7DOng+5Wmy1WNEF6i7B8lOo3L4iEc
k6+vw3pz5C/Wt9hYn1EOJkgP4ilZ38ZoqzxdmcdRrAPeqt8RBnq6SP3WgzI3vmgehT16cCL7P28w
WmowckwCuYOdHJ/m+j2bTg4xTej15UXQYv3jhZ+ACURaROrdghaFlSOV/zglg4AfxrkqKIIgJ+Wl
pCymFBCV4C29iRN4+fgufhP1YjD2cikaYtlCd633JoLD14eUya6FL6DGf43MXgyAh37m7bRXbpTr
G2dsgkHJwlyKQCezqAD/W6DtOuSwfk6Ix6m/UNbJCz8zyCP7LklxAvbTWvSqGfj3c6gDlkW6IUT/
sMxIlK94qVTp909WAag52nXaiurt3NF0QptRkwObXRhUxfirjfbgKnSH4fBeSPDJvdtywMDUGgtx
gpaJGhp3D/fPUVjlP1XhY89MKEwgQILgIXdxb1eAApEjlE9eY4j+j++ETGOWFVny4zis8wiKqSza
ZEaE21Qa7Kc1x6hF9r17gCB4LoxQ6qH7LCAkSYhDljeSWBU8BuDPSDjj37l18aaOWwB9YAfU83pR
XMycjuoLmYwg29rjpqY3idcamw0N8yCbzpaKy3kSBEGKaC4mau0+m8jjFvN6sFAwEHP4Ixt2FrZR
AtZ60yjZ3j985AbYMjGWzD40IQYNSujJBadGJ24u6VzUkKlcIVTmSU9AqJPlGYBoKW/ceqquN0j+
P+XKeDwnObAl+Eiv1Ku0GdjdSonjEstL1k8Zu4BQhtfaiLeGI7cbj+yTgHjZHfNH+LiEX8tvgo3H
UcynsPdI0QjbJVbK/tGYaAuDZ7gnDWvqg82PuFQxMJqhpYC1qnVMVa784CBr1izgjEyDkHmQbPnW
udq7x8frenXHPSMpI2IM+ye7iFZmrYh2x9s/yMy7B4tXaUXEjcz5dPU+Au/KDKUyM3qpVGmAMeky
OBQBuuR9JmQ5uRb24E9f2t82lAa8PCzwo1nx9MV+0qMRt3Znd0p7FnUQ6J92ok1LYtS9++KUfcgJ
5wlclgVBwr0TUZGK58PjPkxrPPF2O2ziEiq8KH0X6O9+H9mPNzGdGlb9YVIk7eZclIwpmP3nWZBl
WXYTVJdxLZERG/VsQAZKUVRPW99HrLLXYa/vOlnbThxuM80AtUC3vVRxsYNGGX4RuZlYYvOB082H
zc7QD69CP/vV/D15Fg38mj2HzMyfCP00R8yZ3o2EaUMMdmza5T+VG210EnRY53fDX3lv3vjfommP
t1O3SxnOiou3oHYocjBSvm5vik62ISpRx+Czaix53HMPErzjAT/REX8ATdRsL4n+/k0/uXQfIOVr
dC6edcCGOoS93Xz5Kj5e90PHDOwMBa488hHcwQzRcyCVIbF6ZeaV54+mR2lJKhVzW6+7ctISwWsf
5TddbAI4DuEDMPknPuWKL8b0jVBFRRZpmDJYzg5Z4j3KyZ40JYKpa93StxpU5udyrsMSDabtpD+f
SDT+lCqaE4LrP0riztgcM6P/1GFzhueXl51RpC6Ab06J6AkTyHEr4UbJRN6oHgN+ll/r81Jbf9a3
MSpBEZPIXiYOX3ETBoJsDFSUrI7o5PWbq8I/c4hDYrrpUF6Ap1fqLmYzYFIVThyOGErvYYyFz44q
kBeCsBjL2PWjaTYCHuUsxGwWXNbJMduhKx51zFmFfTQynj61tV7BYWbtSBn9U0Rw6lcxFbtlaoiz
aOLX6vJX3/v1nI9y2FhFs3yXX6LeODuDWN+BCtONVO39llrawU0V8YFJXKnWY/ZC2Prrec12tU/v
spf3tmF5XYdb7DdkBH4arX9j8hyNhBWHuCysgjDDToOqo6yJLqXd6mXtLkZJo+BVYMOuBNO4Q17Y
hyWIx/ONPiMSNmxmV106BPtZa6oW4h/fec9hFZO5m4J8gXhRRDgRvck8Ia0BkUN7RPkBpaug0BbK
yKn7UZpn4RKrJsMeM8B1V8igGCsqmDwE4LTOYEgoH5jYgaib78ds2t8fkUBbsgb1OCtujoy2ulq+
o55E8GIRekyHKSMtkB+ON/6mikyCahUiq0aG/43kDZF0i8Q54Yk5ctG/i7ZhpCOS60mOjYRrCUW3
tVA2cnqtxd3cWbR7eEFfHB4oKDkj7FXA/GkmMB7VCng1nP6DJR8yhFlbs+sIfw76T0AZyPEM4MC7
9mxe72mp7IvPeLABQwBikwIhqJ6g59CLqV5Yqf3IWawVX6/NEOdb7cYlD4uAXVL2TQncQh2rO04W
c8iQpFWP7UlazkBl1PrXYfrISpkF7fZv6FGWy64aCnfX+yCyh/KZGFxDY5ZRoWgweCRt5xGgDlyK
APSwQJXOcOyt+CV032oSITp8e6nXSF9tWmh27WoilVRysu2HTBoZyDf+H3QVXNDadB0CF+Y7Z218
DlYxr6RBqSt12jBUlByS2p70otVyTieCOwYxIzf0tmF7bN8GH9vvt/EVrx0lZPu3c8LKW8rCr539
gitz/+m6eQ+2mVEtNWGs9PzVrFg3/1p4KSXdkDfYrY1bfrkIQbNua4biG2LtsmoO8tqLxDpa/c62
x5+i3ct+3vH0V3DFEu+uDFW6wuRXYKlh/fmJ/a0gJbqTqMJ6TX0vGGAEW5+JbrLJoiT0+xpLlfIc
J27GHFjEFWp70FZ0EX/AGaaulYJc0BAcGgV0L6D2GtDo682lMUxhWN3ukG/NxdqFDwt7TkMSc4A5
xwesW7ACd9O2GJ1jAQir4U8mnxbp36gz6ODzStiJa0pZl1UxO8HCLplKXImWJuBFv7jzAxEgSOtH
aJV23hlgmGLhM4gz+S0qrrFnLPEvDg8QKFuZSLBOU1xXdJ2NM46bye71APZSY7TQA0AbCHEllT3M
sbvw2jTHC9mO1y/wy2wrjE/SEmJcp3o9urka+K3EzcEdT660or84gX3Ec/2BY67T2oxWjesGSW2P
37so/Mf7JU+SAVqakIw2xrZyFlO0xUunviTJDjBgKjT24EC8dkEZ//Dzn6WWKeCuDlwdgbAPTjC1
W1Co4725Sq8NrB60fRUGCtRzNn8UO204B/5wgojQ2/+EPtEWvVOlnOJkkTt90AjOUPaVIRc57J1Z
YRucMglxWEftH+xy57aWofRVQE9oKlDjTDd6Q+AIETdtuHpZRcIa9vbez67iC6rdWpw/RnKzU1+d
0qcGmc+85BT1AZ6qOtbilr87J+9z8gCjZlOEIVSElbLDf1EjMa9zZbJFsa1Sf2DmCRhO3pmUgrkH
rDEm5SHz3FiXjUyZKlSi48m0F16wNS5RhpnkvhIV8MktwKhN11le+osBn6YdJUDwIQ4DS3GhSxV8
CXbGhWx8daVLe/xa0JY2rsMTEOuo88btNkgYC6JWjX0dfO2zr56YAWC/ZHTOP3tNyzsmNbaJODnw
oNe2cNbbJkOux4PFe8aKihBsqgwn8JOGggJVW7dswuKCUsgfGJt0jMBu1ERq7Pv4zW4j+i5IqVwL
353JT9+Z8EYGRb1pxsqprvvnQ8nUF+PjcJQ+qH1RyJzs2kc0lc48MBY27bXBvMqxlw1viXK2FAwi
JcivlS5c2xlKvgewa7Q8T/xNPOsYiVc/tMkxSrpcrjsFp3ft8t8pIN+l+Vhz73QdXS6/LihRHvx3
2NFcMYx+j8dY0xmYmr6WpwRuS161DpaPNfRM8VlZLNqX7U64Eq6QphcKMsF+7LTujxRVXnG8pmNO
QJx2pJzLxVa/l9g4jBO/AtJBRJpwbPgLlHCX7erKo+Z6Bsi9D5hlQ+ZgO5PTdY8NvaImrzZgxXM5
gVbqcvwpMp7EHYPHy0uXVbQs7gS4mZXZLmaa2xbsYL0XLdQ2+uOFz6FIb7a6zCrjJyQBt+s0tIYf
ZzcAexIIfhMtZXlx5r0I8qEwQ3zEV3/3MDmOCJdRgGnm3oiZ2MRPpRJIfDul3+U+mlPhmYsaMb1N
qFWCjGVqTolkKxel/TK2NfL3Csi6Ghj7lHgRmzYnKUQz0AN74pwtZ9cGFV5OUcUqqq7zQFqKT4xL
yv3fiHrkLohK5xJHG5OHELx35YR2VjoA2vzUxmXEshBHZDApahTghUGuJL0UBV8iBHrA6fBlG8Wf
XIbsGqz81yh7QEFLKXp41BL1NwW3PkUqgJRWCJwJM7E5vIRB8lh4qK7C2eUjeCGCfAI1a75ORyso
tTj3aPLwfO+du+OIhEreS23cUcESu9PUHHvNYMJ2tMF59QBfTG95T1z01HOh9Ks6d5TPQTIeyN5y
eeVyH7u/vevNEaxRB/Zv1jmPyQVjObHvr6d/8bmVPVQ/HtMJ0li6SYrGptiDNDs9g8DCVD+xkiTw
2M76/g1BAxQdgMPeP9srGiDPx5jnNKMJKIPuRB9uEAhthb4UkbFRJGK7WxYOY/xFbUtrMpqCu5ob
T1bkT3x3kFeuy98YCw0thBwbiPQInqgakBA57K4InjlG4xzI1I7tCyR9t7cUOyChNL51wMIaZ5LR
AmA/hSrl2RfLt0RKraMU/WXrmMdTjQQXASgs3peGmkB/8cTaunRQwk95sVAqkBzry3/ahozRW9kz
Now6jf4+VoebDsD+7tu1dmZIsC/6d02GMyhJFTVUM0dyuV8fAc2CvcpJ7ycNva2R4N55Sy7Hqx8j
+RQSWI3dxktBvrMYfBH2rS6dA84ow7DfxDEtLfnuhLTQPDPzWZZ4AkXoP6c2zBPLG7UushT8GJ7k
+k8h8VSrOx+ZEpNRPeFWYWtEYSviBajreuY6QfsWHgUQfw0VKLRRM0f+r7o2Xy5QKauqnO5LpQAg
b8o0bRrkMQgPFDH973q5PEqMrB2YjNjn3g3xqa0L/4CDfpG+WPbMs8MALlmbzQiqj61EQzcx6n2H
g3vvubcrtvpjv/KTmkFTL+eAdU1r/O7mp6J9T/3ZdGsIA4vdqKPOkpKx79of0IhVJWa937jPwCeK
QhL4sYPlodGKhqKqFt/r4DB7HXTdH6Qyw1gqYZznzXMg5n5tAwrp6vnmWy9VfEv8tAx/WlvxGlZR
T4ay6DNuow2gr6izbg2T5pmQAanR62ThwSpCpJkyhxrNQ7xzX4bKPdWAJUMyj/DYL3OBAbdL0/Lv
K95w9ckrOB8dchKGpvb8HD+eB/1vl+WSdpdqfPYHd2WlzNRxbjurEfofjtdTersKmMbHAmB4c7bM
jx0Fsgmj1Bk1hZ6dS9H53V3q2dXP+9ToCTc0cpXqh27Dww75P5NEfbnh66YHS8Mlfd+JLrSvrsAP
iNW6WGGjMdA5LYAFF5t/u3uQduO3KbBElFZ5ioy2FvyZKG74t400bYU1OUJjLfB8oV+sqi19Xb4T
mZYcl95MTbk6d5CbF5EZx0q16fn+g6/oyab0cj4+njH+1bjXM/YblCxXoFhjkDH2GOqAKKLP5ozC
ym5r4aXtafhpjKAnaIgWVw/h28fddFmtN65aeZvhVCfQ4uPvRYmwVmYj7FKt9eOXVO681sD2TYu6
yrH9AvZuqJhVCc4UWBQvnmfC+DXU7WvlD0xJHkY7+0U95COrV+oyvyUgrOuYAdcHjnoGKmAPhWzU
7gz3Rw4LhpcOypMqvne83WtlPYlSl/TNH6uOkN9tHvb9SPtq8B0sVS607a9f0EYxrah980xD+WjD
ntURp4RWgDlyGhcsAEr+GjXNk8Y/pG9sXWhzf4haVtRz6cj+8F2gMH7m4tyQZ1d+Z3G70gsIBMuW
EoJ19MQaU9BJTkCKxsbB5cOIQ3yIYynJyQKpbIXVng1+ZvyNSoknjYzBzDu12wtsYzuA0W8tZYh9
NE2Lxsvc+7t1C2ALM/fJ4sPF774dIbKoQAS6XR0wYnFuJyd5hG7gpHIl4m9v2Yx/nE9UCVokSpOr
y/Ypji4X6S6LyRoLi+sT3LnMleqOPvsbOrKtcBLdnpEcqEp0JmFLKlMXLegaWCHuFvFvZRt8YXA3
g/LZ3ZAXogEDKeePRwacWuoeefpb4YBbeqGCeC/JhwkTYSUCc4P7fjm+joKRdqIp7rrQ7+JnMK4g
Bx0CpbbmqNKgDpAWnGZvq3LXlvDYMiJWNhA7G5jnRMJbYXj10xJJaWVEu9+nF+2vlQJClciWdD/n
EHIN3wQc/blHhoZLI5WOi85vM4/U8mqttqHMktJgtibWF9fempNRf5eRqjNxSkqTFM2hfztmcR/d
/WaILNeZdRXGvB2gLov9vY0IW6PJ1PnGDRqDbotBCb7C8cwyYb8KK/ckDsBpavZOEm7lGRhaoPx0
RRN2fSToY28YuRoThynzr9NgzrIZ5WJSb1NAZtljfYiMnwddGDFWS5DpOdsgU/peHBla628QjjhP
fcZjqszQECg2o3YhlhJ1tJgnmbZBvbjLZGrJLBueJTqqoItv0QgfaMmxRsrZH8CGXBy61//1g/X7
JZ/IArknRTDPxD+VboprI0naznCMnWtpBjMmKwTUoHeSHxi1pDQFcowl1c7q1/ruoATxo4BbI8xr
cXM+B821HGMqKlSKrqLy2Wwu6Z4Uo35IxY2noZQSvITmWc6wvzsOh1k1y4TvQ/87f0olW7ZSx75U
4hPBd/+9MEl05Pu7FnaMdfxjz/02kp0Wo4XQuRMQXmthkgONVqGb8Yg4JEHefg7whgJrTKWzSI+K
skw/fMWlj66KXJjqgCJZkgJOH00UOCHIEc+IfNEsYiCITrZrRz/StvF4DdyQ5LCG+uG0nLi/7EfC
Rd/meo+v4kEaGT4NpEzeMFAiU0TEo2j3+mWsutOKCJj9twpVVv4CGh0P7nnQTeEdShRp8Qbi7CVd
WkVbIGwC/YCX8YpsfVk3n0216MYSbYoGH+UfnoSEnXj1fAXjxe37K1rbum8qgN0X3/RRQbGY1lmF
1joIsDS6CdD/jUhmX+qvmCXxn8MWZQrDxyvu3RCwNpFhPeqYggf3gyBHODwl3ZVZSw1zOwCj3bBu
mcgbVARm506qS8kZkyRPKZIMVJaaS495OiGpGl2NP2vwZlK/Dsk6ejvPSVR/BmKWUce/F3ytBRgJ
V3CRbS6J2xKzmbPXqAHXz/eNfOqUetDSq0O5xBgT8TIW55QSc3kFJU/j3ZK0Ct7jzVy2x4aJalcU
lE84OPVIIljzb5NlctG00NcHbPEhSGXecRfvwMShcEpxzX5W7tkcQXSt+OQ+HjxDfER2JpIv+0lQ
uaXNrObURxtHwFfCUN+SvgbBXXJC9HzPf/vnZuQDTLQ3ssODI8AmqjEe3Fhs2rdIVQfeOSBIEJ3J
SvwFBy/2tMmAm6rz9NXXArB72DgiftbSSenjKzFr3SQKkRZv/DEqXBhUPQLfHIxsYwwAGIKDln01
SEHlBUbSUNY2JbMtIWHP6N900QNvToLzAU7f6KX/Y05okoWxHnxmCxjJTK7oC3dkVTZGjWHSXpf3
GM7MxAYxPH6qp0zf0xr/OzBnoD5gStcVKluT/ld2Np/QJm9Q7EEDhnoj5ye0r4VU8gjaEVJ2YILs
CvaNUJX2VDY2v2sK6O/eyWIS8MHrfJ8cUURCTQIegRnUirRCMbO7rxGLYQHUxSEz0jf9kSdigk/9
b2w1e+u6Ww39Rr2L0tuSeaXBIQuBRriOYVsI/EcY7JMc6uRl/xCia802RZOkrR4Q1xEc6Y4duto+
dj1iEm2ho/L4L0TyIW8zmW7oAQ1aamNPeL6akL9nClv9sbZNmXE23Irqjg+N8HrvO7fUsqzbUhLi
V9B24PencZbwX5Gegz1pYJ8EkAtjUOgJdCQgRWoSy9jKUuqyxQcPXdB1sntvGLP3tF7Z7c/NPJzy
zzzxm7Y/m7B/ik17bBh/+viSWcU+B2gM0YjIM3cYvrMex3SjihYmLBcR0NgdSSHp0ZYyexGOOvis
qnwE5oYuh4FQTlpM7L+5WS7kjJDkJdvLb4B9pIYcTdisScTY2HnuekoPXb59b5Hek0llz8lSrR3d
gssQPT/1TISGfNEbr4HuMoXubTv+BVZnSjqte18DUrVw14rA/dN65MBqXe1KcR8BYHxnQ4o2Eeb4
Y3M5kyC8im/l1OAi7MH/3q6BRP2tx1fY8TVSXDH5Pas43Wo+W9gL82l6LJ6MrNwKiowJUr1AUsB0
JE4y0nsCRfAmB9LFXWOQEKSCgH0trUZNg22Zdapn6m2KSaxcCTfQLc7MTj98/nCkLutxpcpEsDGb
Q/fZRYdiFiAtgeG4HlAZnwpPTN5SmVSfh9j2d1fkzFeqgZCQsxE8kEXSeS/CQorhOozdEDVd7z65
LPCg2d8EXpfMaHGqBiSIc+8enq1kS2iP/Q5eGkmqtPn0CknZwbwVExYQstiAY0Mu/ggHVYpmYt2Q
HB9qbAac6L+TsSV+i6Tf/2ffZpHUhhPPdRzKkhazgoRigqETZgkVECuvyWm1SyO51H2QGBSfmz6J
KsYDbHz4BmB+rvw8W8tu353MCaLJLITXUyS1EQijmE8KO004w8VUdAANY5AOAzPiEQEY34BoajeP
OZO1+A/XC9jdp72SsY8rtQYG3qHsyL8mpORp0EGpUvaR6FGNMxwbPJwXYD1gZvinTdOTstWs7diW
I5GT3JoJ2PyEClz4bdUI6XK6Vouoxg2SY1Z94Tz7UK34I8wH6jT0a7hZaBwwGUFpxiwAAfeC5Par
qS/EFDvJ2WZx9ZgZpwdIa/u1OZOItoSQbb6tzCVs25b1+FEje6UlyQUxFjt4oxbp6WObUnYKzPvR
laVnrY5Cohdd7r/IrZQltUFYwbYJihDWYNJc44lp7i7/k7lHymClutnSHZK8/OaCF0EkM3oszoPS
e1oHUHFi/KaAene39u6o6mgP+u76n/9SrMvWpiDZAgqyP3QL6EQn8B3Mf99x9VHaoLbRVLWrA3TC
uRsBST3M6cwXyw0gJe2Ax1xi8LaExSKi1ZCNHcedmDgkCL5lZqhCMKbCjlhfgKztymLEhy74t/aL
Dgv67HjUd+OIVO3RbUyuPoWaHLLH0ez+BnZr7DVx2Miezm9Yidgdz9iyJQXaeo6JEwJmqu6ds4OW
2KFSQ/KbGSRq6kIcyhAFrb8hzQNdsmRMxwVsjPPkkyCDmiLOCeSARLHh8B1zNfTbKvlzjjW1kPH6
9LXdeT8nxIU8E8OMfxQfXrocfgXlsTeHmTSk1tV/741E//g2+FdeYP6vZOKwLdSLESo6CkD81qS5
mTzCx/X5LA7odhzuTopiJ4lslY2n1GMXrjOjgIvduyf8XGlHZwRpHwAe0Aim6VYjYmyL3R8mttrk
0IU4K6xMXt+cmWn0luZQ6CDLtyRW9IKTV8h/QIPqaARPm6xGdYkr9tUdrr05KbQt7I4X0f9Y0vKF
IDIWm6wwSuctWV9R0tZ4p5a93y1Z913cRgftSOtI/yzkW8bE9kBwIDZzF1nW/vGNnXICQ2FR85Ow
elXullprVhNmqEnFrY7QjxG/0eH8aV0pr8Kge0y8KT9IboEXP/HODpbObeqAg18Gwf3J891D/K7S
p+5pFakrqVKxwSRTnCzYqXnVQgpBXqOH6qRazKNhHtLVuC2aJ66GdHmj21kJ5vc8WO1acdLW0NbF
k6QjhE6cIgekK0oDO0NQ1TC8Gncj+dEtaFbntCTjJ13A09b+yZ1ga1sqzxmHlxta1TT0J7MwgyH3
Y/Asv0cFuuSEP0za8E4vS8K3Nn2S4h46/R4kBK0FAjM+/xJivCpecvwPr8yBJ9xV6ETon3SrK1cK
K6wFE4T5x0GkpwvnlWD6kR8K0zAABLOCLgHutpqk9ghheqeRh+0fzCyR5z/Y+ajLor9DL9GBOmRT
09W+Ss33NX1NGmmDHjkpzsy41n+RAH6IKWkhCNroeJYMPUW9DjT0M2UtEC8FposWYqQFgmtqFtam
2Qy5CRi6Dy02yEgXddWgiqjisOmmPQyP8blrc90bLJGslPfL2LUOnWzjvpOOfVDFUDZBbxFmuw7D
21Y0wBONYLr1tAanmGvN+2Rucxza6U++rHao+99RynfbddMfQfmgBvyqAmPVX9gcnqDnLYMdnGb9
YO/OpAMCFkwF5fYA10bhDzKLkw++gwQD6rSpHBuQoL0PorcnAOArNUcPRt1DAvp6TavUMjN+gLx7
zWja709F9yFivSOdsHL1yn1fcGaWa32FTGGkic3U1cGkk07kL+dRnvxfzUeAs9HgGRkwAeolPoxG
AIYccYWiOxuPTGWr445ICOY7vxP8EZlfoqS5J9QjgNklFw9embiyHOQ0u5CWzUQSAI3K7d5bF6g8
WT3/qhFUU2GR3Hr38jPGUAzAATW+0IvuHmWlogUKdXsBsaFOcyhdFlTzGuAVossur4N3mSF+v6BH
WNm44HAbKa68uiuHwlnGPoXbUcP/FCva+/S2+eBmuAiDac9RGZHarsneXcY4hH4AV3UfRE/VX7QK
UAZbz9eo3LCgI9OZVj6KBv+5PO/G9mRhHG96lxnnDg4GN1OXSz1B46A1GDqAP5fpnbSsecZgeQ72
oSaVKV8yXY3Fg8FNJU44m6Ev3YjKBTb/tIFR2Wlm82AVIUDgmgyX+nc+wl1P/55+T4lS5vgwPq66
IgNWpQdctAbN0FcyBJhcN5Hsd93RskltvenG8VQtp+TFCqB0dlsiwbkzA9Rgs5Qr1oQeztrP0S60
3an7oCQ0fET/K6/7JcQyJpU7BCiuo7idn4pPh6c65Ac/GjdeyrH7OeRkVnyFlZL8RaSN/OWjO7H3
b0Gbv5STgI09owbjGk+tBpweDKwbRwbe9jDHlI9YUhro6u2r5u4mEl1na/0Kj7hRk6AryzJ3voc0
lLO/SPExmGhV3x98c0Ss6eRTjTcj4+yKYQh041kLGVKc5awiCrjtP1ZD1FrUTM6PSVAGTRp32DmM
p1HeSOcQnPaf86A5/z43Cu1P2yYKoT7ZaOxpdhi2lzXg96oUAvfU97PqrqnRqA3qsHO5tlaEahwX
pK0vrpRp2c7rZ+tswUCrnRY2pjuoTG5mEQI18gaU3hOQk5JwAKXi79qTBzCRizwC2g45lqaDyJcX
XQUxmZJZ2LshdHMvu7tgIDdgDeZHmWGh3qmh8Wi177nGJu0M0SWWYBoEgBbtFcvxcCXJLlbp7yzq
0I6b5PlKO9Dq0KSXixatwujGUUzMA6mqF5Le7UNuqK7mxFvd+ETGHVzW5U5QAxjUrIAnCt1zjEhM
CL+pDyccm4jnHh+32Kb9ebDdgDAq9t3ECdeOQeTdk45Yq+M0hN3vXxpOYdLEBwoELIfLuNBmlMRt
FKjxcniHnB+jaW9O52RRgEJjanLnMAAKHgfxzC/OeSUyPf60oS71B83wQXQrG5JWgQpOk1Oz9SHQ
gre66k2xJP0E8qqt8VIPoABfOx/9D/cwQRsIFpJlWXXl706+twMTwhyyJ5U2Ibz2TcTS74g1R+r0
TizBZcEgAq73QeMPYVr3RPQ9IM2mp34gQfxs6AITrmKZUJCu6eQeMlgCE9cjdGoLDKfyVxbNx4bY
q8JZBDjm6kNAgixOL2kdmE6SG5UzDW2SAO6+KcMW03H5ga6u9EarETO0pQtYOnrVDHVIF33mfUVi
DAGw00cNoBmirFufaV3CVAHHcmtg673LlcRYXI0ZJOHTpkaeEXC/NnjVddGqlkxdiZi6XUcqT5U5
V98gmvwCzWUAVwAVes8mn/FRh/L21fduNTWFRRbPeZIx8wKI3AZ3tqeBqlUjDSd7PRUGTOunDBjS
yD3hKbya+YotE5ONSbbVtkOIMnfUjB1ju7HXBM7M+zFzQ1wdEBffKq87bTziT8N7qQA/xTIV/fpz
oawG4igomXSQXmAzubRBi0fHWsQN1T8sseQi0eSDHblPXEfsMa6TnkmDMIboyrPWjPBmtL+VJaDL
8NE7ojoUFnpIYjFR2ampjgaeIpQP2GfGZogqyKyQC/or5SRtg/mpVgYAj685zOzZW7A8+1vk0tjc
xIL5i1s7gpXtpSlYbQkie+/aBblx1xkwUaK3LgrCb+c+ZwHus0vGB2876EjVrjypz+a6cUjR6jcI
EDoyHPPJ2q0pK8d+RoNDC0hnythTNXQZjfJ8Efg2pSgmbGnHKkhmTnodnZ3LLkKv87aPBDUuCTFt
TvcE/y0M1UNhPXIvuKgcQdu87UUoQyrHHkKfh4cBih+iyQwjwryoshyD1rpqS/QI9NVc5lIronY4
o3Dtt//Ht+PYSse1EeIt757On44vbs8Gm2GXgXYUnt6lIIiIil6HQrtM9HnhfPXPk9T//zRqVAQz
xOrTou7jcxw75RWu/h0gbZZ8BZ2JozPK7EuVsnYU1l2WKhthr45SMe1OBsvr68YXMb3gwXmReg2J
aZtroGsT/ZRZQlZGdGTbShLipHqhfv38XjYBzaiqVuP3IqN8Rb92SICyVbZ1dqAzXH9uefRx25j+
F85/MMLFhrmO0dW0+yvuFs0rhryYOyZvjWKnai2sVNpSYhTr2ARn+xgQqDCgPFS24TDoSLzup4rD
yol9uOABA0yhg2Z0XmnURoD8/gKCoV6ddP8KSP74+J1LgErDcdIn9/ZEdVTv+N3lUEgU/haLOfZN
ghllp/Dhjg/FnNzc/mOYKcXRfxSY7SzUjOs/Vd1mPz0VlNxLzk6YOiOwLnV0uuq7R7iURzk+JKkF
76x4xeWv40amU1o69ydS7mkERIbpEUm66tEMgGB5XO8uF6sqqZqmGoIHpYXiRwgiZIaUVwn/PFSR
dvdE9NFkRWY1ub98Ls7OhpcviJwA5NdO82tpo+A1kV1cb0UXsZ4Q2dFLQGwNYXW9ZhL2Opewe4LL
6awwcJGHZWk847/nrquXxdd9ZZ2r//nZZkOtfgH84/ZnlU8Wl8UDRrunk9RVQM5mg4iZrO3EeyH5
8kDNInovwTPTVLt8+HjiiNVybbrxwgwOZPOLh3DAWQPDczJEvVDapfLJhpBZtmteot+5fxrkDwRI
JVq+jCXEHInyUWx7CvxniVybLQF602o/gAgH4PSFRNUpCOM1etYE13ySoDL86T/haKMYwizfFbXO
SZEJQHRbUmAPJGcEzSER0GQYmfNunx3awpTIHMRh3bndckCGTnaFWoZm+BbCIDJFpyhuWCa8Vlq5
3qS8KTFURePAng0tXgMui6lCVXXsfBaJEChoXY6QejasHym+HAbcqEdP+42d8dxH/07M0z/qZ/91
b4yYIDJYVTwqhgpeGoOP3mhuExp4Gh4GwZoxtrPaftnMauZireOBpsOc/xxi4GWJ16YMJ5TKMjyG
0alBlFo0jkyBroTjjnFLvW/UgIB0Xy978Te5oUF64/QFX5h0p2Uw0wh5qPm6AoZ4Zk8pT3+yk8pH
lOE7V4Wsvp21Tit9qa2mE1UN54juJHCANf8Q2RzIqNQHWTioT5MH8hgJOutO9+asnbjKqog62TuR
HrN+n5wyAKKCcbvcpQIQl/Zrv+pJ71+wjPn/Zr8r/aEq88PKdEw6/JVaVdfrC426GOvw6WGwC3pA
6j0MrwRyD85USMOJQFHn7w8ZPNunmUL4mtKTscg4tv1TTlmVTk5eQkPhAAVu0KHR99Z/X6NJmt0+
AyWs933etzeWRPONwvB4DGByluojGK20ik5/2k8q04GXUmc5VyBy3A9QxsBbmsY/ygqgXF6ooQMU
eEWYA7LzjksL32dGsP2sOOlpMyQkA5x1jdO6T8XZEiKWJTNPJy8mhddTNRC0R5pjY9KwyJL/4cUZ
NO1mwCK+qePzjyc3h91IOlWPoCLgkrbQkgsW6utwvEGzDnO8EeK4CxEs68wvZfm4Z3uOwatKsPEC
k4egY9exVWA6M8Al5DAOhhLCSdMWLLkIqEpKlfWrkWj+34g3shcOjIVNx+Ym/ho7bRE1NswhdoP/
eTVuqSUOC2eFooX0krLWdvC+6tnhGcY+3Vq+JW9E1BoeIok/9kPaZnJDV2L3qDERbRt/A85CbebZ
idRQXwF4nvbzbewp7xiy32twX91AtAsSLCm1Wr9iiDqOGw5vHLtoSIV20oxVE7NEDgs+/V1PIfUX
glk0oTBtLfeIehKsYg9J0ZIV0S5estLYh3/f4Uu6kIDlWKlRbZizSA4poCjjQMNB0sD0thn35NZG
8ZygjWZwMO4sZ2ATYjZziGTZFVPbnp6B6qQQ9A3qPmYEs5UwZWD2Rv3NUmkjB2qwJ2hjLXwPaxle
w069DOKZMWC9AKWQFAe46XzGMn+BCVsSjO22+VvySNjQS4VQ743e01mlRY9P6dh88wJydJhFCNKE
6h0lzky1G+hKW0GtcnRigfYyQk+M0ucavAF1JO9XEvmR/j+UjCqfd7d0OfcbgdlNwS0L0BnlTiin
ZDtesS9H8C6pnzzQEs6kNHUJ5k2In6KDvxND3A2z0cPeZ2eib69kIYXtc/VbrXUp7iqrwAGhjfZ3
kvdaweo5iqsMytRGfOEByHsM/ICeHawOC+ZdfbU4UK0+dMSTvvyBMJgzmaGxTsw5v4+OPWBVS3HT
fqH1P7+BOydyEsw/krDLdhq76acHNEv2ZlW9ZH9He0wjD5cMex3C9Qs9qwhutId6f5HoxNnX5b82
/FSyQg/gtf2Q7ErKnpor2W4KwNi6gUSZhE81rEqDvaiKEUP1XDhJG6EoG4v9gvQmvLQA0Ndv9OBe
DqaIqhTCjCKiSJokkPhpulJ43qzyF7ChENEtS1k3Thx2FnXItY6tIfsVhwDqDajPKfyS+a4FxXMa
uuZpcaAZ5jxJjlx1Sak6YlWMFxGX+Kr52MzsASYDQhph+RiZjKzyOlq8aS+dZMRiBiHhiFdKCTFs
6mJHpwtR7gp0pJqUD3eU6HP1rJLZ3L1uDgsmsRJAFygeWfT6skF1yJ/uclLYBWa6Ydp/psHCbUbw
+Q3Kz5ZxK2bd/XhJClRo4ARiT5ns/u901RKu3PAzo0G2jfAf1Fk4I6yw67OdKHhmYjm67/UNKNAI
N/X7/ianYciA3ydaKOuVjjbK7Cbv3Xs7LpeS3kPFEkOYd4HISow/NMWq0tjM2JfM80c8l4w97W+x
dEiKIdcu5+rNey8x9jSxb3BCLuzcl+TaHjm/QM0igUuEppKVt/UwL00DMgVJZlJG8vik6nq4af3q
RT5I/NFKX64ZiHSvZWg7+wWvEWJ9RRKSN7KJ/NqoKo2i8kcPoNby+lubGI0M5SpKxSDAr8sV/lgn
Z21FBHlIE0nhCdrAIZNjT8/8CnEB2/FEfoGvnY11IJ5IWFb05Aq2PqYe1vkAMGS947hXKEm8hUmP
nZv74KgRjWjc2T6NPmpYZm0GgWzKHgjqcZ7ltlPXdpWezg/WkK813M4+gVFixYP/bq6qHu7cm8Sb
+4fnlQaiz+zSIFA73WNYLl3x1pWjbN7M0UW95izwhdiCkR+/bkS/hkstLjiaRyBl09w+aGNzfv9E
tIqJzxFzXtQHSnhq6r0evY+p68bNAwyGTO7hJcA5ukt5j43CpDtkxNNfUtuy1dt6iUYabPp+wx+5
SfcVWcHbEOps59fh5OJxpmF5/J7ZwfTAb72BbBemyCt+mkiVVwvM/4/LWSzROiKpN5TahN+SiPu8
Ecf5uX2nsU05F4XLWI36+P4OrijjgsJHuFpun2KhIfBq0gqu6MQ8Ndt5HK6J/iQ0x3k22rTixGyV
ES1FsCVFNX8iLJbNXZpLqdbk/ydxdx1ME+8yW7QtUFqLPbYADEob+kPccKMoCyIV6uha37l8VlwD
9yWG9o7shvdh4GMxSiVwYEdwTJ6MhXy5+Q5ykoM54QqNPKqHcoNxAp8eRMvseG2lHCAuxfPHJ07X
KZfL6YP1mB22BR364baicDRLhZIeL4wczhLrQdyy28m2RFZIw1sns0vS7Opwdb3oWKX8/7w7pQqt
f0X0exi+6ZXAJYpJ0v7w1QACAWZ2HmPe3IHEDcyn6RAO8SI5WupV3GKRzKnH/hXrzV1GI8hanD7v
rWkM9zRtX/HqSW9VTkcIPbIHwDltcED9K6sVfIj0qT+3u30qRclSBJA04sFRAWcLVVQAqc8rGBGx
cN8qNSOc7IMH0ZgD9IK+C5pQuM1Ab2OCJ3APuCgLKjIGW7JNxLZ0SsYJtYGZ0vYS9NcnMmRhmY8u
E4BDG3HTqHLKIOwBvyOSueHNO2ktFIoReLoe6K5IZPpsUtwJZ2Jp1GBSkBBWdDcodnLL2D0WNBtP
wOBBn9C4jlRDcgz6R9XqApj9ABS9ber3dfyOY6qyqIyfgaGSh+NB4MMOGyyISR42+0mzkUxOYIh8
3z3sZqqxPYpSnD4lt9CK5W06UOGwoz8iO8493DfWik8xLJKGGpeXRMjY17rbvc9OWBqVXnV+rJ05
XCqTu9KEoLjpmIE9qsWs2FXACh1NnVATtEt9fmVstnrUEX+evDDsdLpDpwuSQtAAwNr9cwhgLTXp
DAbPXN8oZnd701yqSpM1wPv1+46t+BDqwhHFoMgEw9aW2wAr12WJrvzWSt08P2ZTl0eADoOgXuD4
D4L6rZw0mq/02PRWf3HjDrifHyjNwbfFZQnE4JGt1A5ZjTLzMuTnH8gKP0y58Q66laxtWFyK+Z4J
9ZzWMGS0QQYQGFptGVcMvYJHpvfOqGmaVBbxqHvlICvhwm2z8WuJf+1pksU1ulJSDRE9wGXj96Cz
aCNDyXD5MQwW9oR5dnG1fm+ybtSPn1ZFI6ee0xKBrp/clGsFzIlPQ1Fb/ZpT+Hyi1+EWu0OVHW0e
yJHloV6pG5L0gWDBFLAi7LQwmFUhBrcHcSAvWN3gG4JHhlN74FpnHelQuVKl+hNvo0cYvBQ9RG2z
Ht8+jiljHnQ7iobDTJGK/yhTS1EPuUr5IWAx+OHHFhOCwLHgKxKGJEgvDKB6Lp9bgp1yBzF55Z6o
7nt/Zi7ZucgC8F5OUksRS49XW65f8yp1zBOEgsOPEnJS/51eurAIVf+qNXco0RXK0YlckIvjQWOE
S8EM2vnTFB896u5mTsh64cfiVCqefOmzhcti76/rkjBVgdhKNxq3TcFiLs/pEmZGXs2lY6n3nMYs
bf4Vuibm/CG4zzajC24iv4porlH6KZR0HOm4IwYZRu1vCDoFKeyxenDYEY28UCgmKzuvGaRNT0O2
h/7cWg1mHulf3GDRy6+NbFlqDRpkYPDEGsUxZJnXkTNxH+0ezRxKOakOBfBsGrcKTrK/5v0uk02s
gPPwbYBueUzGy0s/hf8rsc3p881iHko7v7jpkmdo2+aUtpZqEjionSitK7MhpDJ9jnO3BYLTdWV9
s4dY91wYnRjetUdx1Vblo1agLH4XXBJHwx8I0Vi51u11YipCtSejvdLifOzJ0YmCV2gGMXksWC/l
AHawUEMPBZKmUjelRwC0wpmIwjVbvyXx5yZQV5c67Qcm5tDEuczAUW5KO2A02x6cZEbJCmSZUCkv
NBc+0OT/EWrn/1boD0nRY3iUHiq/BTPou3lzcCUsTVOLpVLY3XzoeB6Q4qPnMc7OmGjVgjWHXtOS
q3aJ9s+7tpGN/pf1a2G0dj10khLpxafsteOQfxHSjVsFJySiHhvtYadnGgy3R5CqBt/U0cMeGrFb
8v1e+2kOPDO6yRA3c52ezDodAhLixEXZ8lqMOhciIgTqVgTIns1PyPSbVaH5vtPawZG34UoLkJTj
EKdpNPjEEZQsbE5C1PIfwzlty0LaxKxy502O8QykfwLxsufqZJs/bChEfKBdyfllH1JSJI+ciKqg
QaJ1J1rmqjH3+G4xWJ26x82drUBh/0U9GkkU5t4I0GsYNipyyIMnoQE8qxuECE2Ear08yPAe9gxm
PbzdScjCYYVqsiHUyufHf0qsuQI8T1KHDlJigZD8ci1VTy5idrJUmI61OcJWBZ0eP13Lhdn0UjQh
U0h9rPEJItfwwodqmpXICRyTLQzr5E9clVhkEhbvhShZ03DkwK3rop1rVL7e0yDUxmaCx6azqbjx
HD5dnw3+rfivIZk9dhaAGAlc3Cj5nzdf2EvcsN0ZU1CaltRMYyZbN4/zCVkqBkwvOwzaD7/lS/mO
rRK91ZSDSdB0kA4IU4ks3wluznh6b6fomeEWojSbJ1D6Ih+jJkJ4JIPQrBm0+GltOtDqRMLiU3u7
N4wW1vOE/wB3FEKIPUZFeGNX23AOxV6M/zkrZXaT/O9gY7WVtmhJVZov/4pASsxt4pCKex8jOiF9
6AbROJfmPGEWtGOqhnoso6ECiMNx6OBEqNA9qNwSRVeX728diOqlZbLLffp5ZhWV9SeNFbMg3aGH
qBi4s8y/9LvDxeHer+Nlg4ABQBksy4qeZgdCkGp6jbHHLZlBsY77RA4HyTpomA0jMB8+UwRNGYDn
KoonxXrGVV6COdUpRDZA4/nwM7BqC+t6NJzWm9TwL2kCTLVW3zMAlCcu56znyF1Ww2w4y34oSedA
vp0JrNmQ9H2oTj+DEO/E+HaVGnoTGMsBhdeG749sXRU6HYAcdZGCz4yvRhNHK6fRWEHoan7C2fG7
eH5HaONGHy0ynSyFYgU4WQt8R5AecAR3DXx/9mpiKe/qvdGiTorblES/dzHjS9XBQWK7LfjVWqFc
sfk27P4fLC2pbcLpfOmPryXec1Y2NXeoINr/KshVbmZqicrKdZhI1rdbc2COtjKyBNbHDGvZUfaG
jlJ1mUy/B5MV2UzpKcZKiowzmR732Tvn19+z0fiwG/LyeEVoexINRMt/j469BACxhC30koRYmmZG
Gu4CspcZzp8JZsQ4+oWpvR/F9beg9vmeGcSZHpJyFTHhDMwdyvLtEkBmiAUTp5+nxfy2iRA1FCKh
0ZDAXEjIazhVVMJZ5aDk0XYzD4KGT8tpUxCk5bNGI+TfmKMECfsclXD00TvLEuJcJ5GXVrMVPQf6
pStNqzrWAG5ithHxz5bkLHcZwsuMKvFiDP6CEX2++piJ8Z+IQOZVP2JIjKeTmQt4arSBV00ppRDh
XOwz7Y2MdJHx9YluKCU2o2WTfh++0asvC9tdL0RiunXMkSKXcY4VXPmHiLQBfeQ+c44J6Rsrx18L
en67wAHgkBZTiyNRmgUKlskIy1/pBnnqedDc9wpnYQn6/9vckP0hXWsmMJ92DOcstH+4izky8tZN
wLlTxxWVTI+Q6B5TlLUPl13bNj4KVGXMvDEPzkqb/2JpXYnvwxPIVpGtHbp6LbyQZbfzsvnV3ydh
BBmboSvcjEnZVKEdRe2KvHhk/s9voJFJyzO5PSj6V/+LBJwhxt2LtaNtMJ84wPOouQjalHR7T9YS
TNDSc2ALNf/kTtWgn6XBvczrarsD6B/LLuWe/+4UegTNrjdhTiiXKxHXOPaydlH92VCoAfRErsmu
T+KYWBqZRChm1vG/40tTKnQ8LYyEPvFOfGOueJFuu/JQ+HHkdMxlvcEwep//AaC60+9EM0IjOz6e
KwIs91weM25loGOSlwH8bfsSm+s+/F8u1jeuwzEacltOLMPvGZAGU9pw3iKtoneNzn4Oshst0sBa
zFkzPY+FP7U/IfEvuq86hG4NKdhxG5FkpF5dbfDSRHHaBq/RYPbSk56WW8m3LyGJWuaYyt8zDlC1
r4Tj/hPDjrbsIBb9ip78Qrh5jLR18tyJjdo6A32pXHXIbv/3L/vQZgpOtze9FYH52UKvenRiV9Q4
n3OCDyqrlekWtXni17lj7/jHAAv8v3ixcho8yQg0xyh3fPIpLkbXeaXFftFm+CRqEO3jlYY5ih1b
kyAyIUDJTTW/gyP8jX5g1acG19HzhM4R/F6FJ9dcXSFBg4+d7DlSpXzQXQyisMaCS83dPgIgx/ej
mliVtRs2mh0P2LU/UOlcTCawturjiFLONJISeZvFo5rFyhqSTU9+Wgrtp+BKMUl5//6N2QOnt5DY
2nkk9icQ0XrieigYteqlvPmbakVNkQe3og++Z2oxQXugx22mvk9x2ntQjrH3Swx4hcQileziJT0b
1wzqULTTHjBiiFkHZDDlb2ZXTF9GzyRUfrj10F3lzGoteB+ErPffggN3TxHxMKGZtNUrBgqUecAl
7n8XOI3OradWDFfjlLse5MH4uWT2+fngjBHe6VQcab/6Y3BcVb4k1VC0dTO6aDlJQSmXoZ7+30T+
h5EsRDbsp91PXEii3hFp7WAH4MRzTi62vQvPAgeQPwg3x0ihav4aLM8mSt6pOPp/C4OFoEFOP5gr
oLiERs20mSrCTWHNUUP53c1WKQ4MOCWP3uLlqv98kz6XTeojHG3+m3ahQssYf4kVN0JIEah7AFqf
51ZGucMqXm006bzamSGw6+P8MNgDcxXYcbOoa65Hc21i4ZSkZmH/o09O3csYRWyD/QddW4WOwPoY
li9/MWnOxHX0Hv8zyhLjeBMlzKLZD/XC205hyaf6Smk5AZuOquesWEjTLl7iNzOtj2EicY+M9PQ+
Sz9yM/03qolwQH3mLl3Dcqz0eo4h7TThhTbo00Mnnxo4ypjXfmiir60sMlfnUGTg/KXOJ30cUEHA
7junwI5ShMXSsIsy1vlEoshLpCarEqlF1TKBCIgjtMJzS+SqdaK4JeG1pbt1IHFuEr9m7rXFTnwq
5okB4Ig7j5PpXjHNlNmdR/eByf4kMSZN2AT9T8osttGIlSfYTD/YjC5PMxS2fXP7CxrP3Mh0VXuu
r3TZilEOR4yY7jBOAuVuqU/02GAqccd7gNWUSQCuD4tIe6chldyrIVJ0Fy89nG87cHFpwRL4/baU
nW2YP86ac7AEiu2Rom+ismxFh5i14WTxn0TYPqwLdA2z46VD0ba893v0jQRjS80sORpOgj0RzKh+
btE4fYh8t6Lsri/QVOX/xLv4Wva0tg8N7kM1t4kkKDMD4NgNJfnokD81K0xNzyIDzi6HzI9rGJDS
SjWlxGZnLZygC2kfNKO1UPSOPleQDGuEN8TP6pvMSc0YJpn4XvCRwnVN8XbfyvDGPDGyD3n5l57p
y2MlVRLjp0HGN1/tbakbCThV7Wr/fhwrbKVDDoPxeElgIp6E91WXwKw1fv5g7DJep0l8lukH+SMy
xNn6OT1HajEIFO5LqjLf1oery0xGqLU51l0ALKoXoe+cjXeEFrXBeE8U4VljLh3kcCkYhNlHeMkR
AvKeaEm+JJq4wc11PFg8iQln+pgmmrAeqXF3gnsH3mM1QCLRMlNAB9/djKJgEb8mVctg+0I6oSDc
5MvGOQdq26HkSGZL73hWmm+aciir/FC1nw7K+RJxbdhiLjJT3X/cWupOEepJeN/R/o0nI1+oZE92
3Un7wlHSySCxSJAnuRhyS5Itab0ERu/z9+dEqkAHNGX4yN/JgJxP6M5oXyOYprAWmi0sR494vc0k
TESUB3ZCusifQ3uEg3pm1KSbNpM2wASpLWCa/w8rntPkZQUh+mp6xgSWWSxnZOBowaN8E5OxpsJW
6PK5zh+xEk0Vus8+KmX2m9a3/S4rdivJsnr8X/MXd6MVsksMqJW5Fz2N5hOEGQdSvXOJiOltf1px
yNfLAcjxNXEu8OJNugqO9WmU9FZjB/fpPQdVz+crVsRkXMppqn4z7Y/159VeHSp2Z7aohlY3PEw2
6YtlcSsO7VEiL7n3wp0Guj8uCYDEJ8cSdmbIkIDVeNw3YVAbJIHyCPwA9hxfKRdolPctdTQv2TO5
6+kPUkMlnsW0no3/vti29mLCfyj0IJYKLBO4A66uXjNkapinaA5hdmhgsOQfMHevE9pGUPqCjOj3
Qok5LD3Q7M6b1O6J8HXXKEQ1eLMribkZ95A5NU0aZ3BsOdcSU9ye1abLLAUQNfQPx/KusEkO3MUI
2XJaSVZ3FGRv0l+ijE1L1KPuX/vB5QD2aPq6P4WnhrphN3OGX0T+biWKNV8MXh35LxUcbAQrW8TF
wYBxVfcxUKxjwYNGGUXu+fNO5tNvslFJzBBBpssDgKis8addpNzpo9j+wuXotdDdiR6gjLMQquAf
56HZVvYn6Xucmp/zfATCHXhAk0FsC+exbZYPMq/Pnnh3ovzvn0QJ8W2AEr+QCjCd9zLP4q07R/fD
5NG4umzAK6etxKaH7ZSiuXlYeJGMUya7N+P1jCtINizeYlf7iOZQKR3TFp+BaQuw/+FmcGiv8eQG
XpixBncINXPfCKuJ8ZwapopBe19zZ2zglqljm8aHFvN1NhASHKUwwqhtBrULsj9vAUMqQJwoAVL7
guAWdvGqTJ0sIYGyYNufFeRlTs4hAqW1D/Ycm7pFbL8bnJPFAYfQv4+a5F5PN2t/zXuJuq2HaSNo
+72wA8z2fsVqJgu0Mn+nMraOsEN4WxiXqb9YftwlW3hsQpPSz/uulRSHuhqaThfyvsQ3Ak0VNy3g
pYcrzYsSJR/9/1fMEax3/m7rXMabrIeBEz9ja8rIgFmXx4JRmSWXinGid//7uxSQNaSDxcHsCgcl
6aNnWsydimf8NlIE3r2uNQOJbF1BT5/lvKiv5DXe5Sggti3q7TahPkN1RjC9FbhkQxvIGWDtgTBh
Mt8EWn3+Q7JwmczbSzuFZj5o3Np2wOAwAKKqWvH+EwxxU/17ArC+KPkIvSzOMkpR7+0Za2YSjIP2
ay7pQ0Qs/J3w/KjKklOLl/YBUGf/JXDGQ7QZml/T2Q7Asi4tYxeQEupCb4zWh0ezoOJyCJRoiAAU
QqhXbP0iE3ojhVFdo4KBh0kHVecw+ynJD1YawjFaW9TqNz6YZo1uHy3Zc4ryTfF4L/OkhmPSRaZ4
UUZ3dJ5ENi2BOrtyxFxBW6Or/G3FNhQoxPOUq+v7Ergg88Ng9sM0PIyQcxwbWGMTqReGgfn4Kj5I
1p8m3SnSaqJsrtwkzVy8u8MFbOXWAAh3UcaIN+Vs1zJbUIOAucdHk3DLpe3k0JOOJiOlDFIwkR6K
tGK1LwMKQitn8gIYqav5bes+yTgBIwF1FTvBW540CEeQ4NebpY34wgxWGNQeWt1/RBvrddYRpI61
2uZCn/j5cBleqQafRnaCgepQpIKg91rp7AMtGKHS/Dtt0jMxda2NL+03kUOrNY1dDsIRqH/0/SxK
OJYKz7iUO1Vz1ZZq6mueRk4XPVaOsJyaPL76JHd2w0pzjyn9G29mhj6iaB5Hr5WXUt58Fod5UA1t
2FVBoMfaWhjxGjWW0LeYix26uOLCp3zX0R5gj6fvS/Cv87e25bQ8OYMHMDn8TDJtPDRer5sSe6zn
90FSKKDmVYpSJE/Ku2aCFD758dt9GIRbdMXketPOxDsAm42l5Aa9dTaIxwqOwVfixckSDiqd9pOP
gp5UDnyf7ndWizkhFwFBGCioqhzd4k+eHy0hyGpbcXcz7u808KZiHVEWtOSw+n5rcYqYLxl7rjpa
9h6lbl6TiV5Is531HfNFi01m6c+5dzBwPxIj+fxpyUrxXjYLFJ6Npg1J9QWzE1XNd8RRQ8K7wews
7Y+cKg4AEc1dC8lLGeR0xwLi6xeNk2rxcEkSYFsMxZqIYNYBO3audqSVzSrJMTZ3uhpqI+1eEsxJ
aQ15ECTjabbBC2qz3Ro1K+YsclgWE9OL/DLfMGvasGDOGhRmE5lzjctKNqrriY24KA61c+ZaNU7s
yJ+PyH3GgKslOjtGlAr1wIvWog98hf+7Bl6t8jzcrcPLCWUqGvwQ6hU1is8AOnHQHq5rzC1tZE4s
oR0nSppy8K2YzeCsWHggcbqgTKWL5exDfwWGr/YZgfrGPecVeE2rNplb4mNFgFprlX2jhxB+LNU/
7XHqppzXzhpV+V7BBMvqg/L9ou0sizzSI3e7a8Xdo+QIkGGOBrK/4rJclGToOgg/uS68dWyrdxPJ
Et99xzpg9aWgDNwi/F0OQgAR2lSjpy3doSlJ5Vt1mtk7mwXw0K8vuJu2sIQeZE7pnxwbQCgpIzfl
OJVrRlSvn4XaXVg0ChGwW/Qq06xHU0bw9CnRVEEbMuvcJ2CkfHoCj1dMl2q5KVW0rlN+lnBjOX0w
sg4y0N75xMzfUw7ZB4Zlq/yDXFIh5x2Pka2zZDduG9K1KjofOyeP2JmWZYBq4gUkaG1OHsWDlYUh
CM+vh9UDfKRsWskqfWSo8qAhDNQu/LCABTWGkQ3GORt6KGE+MKs6dB4KUnEyGl+b6/V0D8K6Bg13
Fb+EfgPcsojqrWTeZ0BDpzbhaOiZTKGV2X75+08WX6pIo9RIt4U+mNshtoOPE3S0r0/JrTGRAcaJ
Jw8O4udg7heBZ+UUlZBpsd+ctuOSAfxdbZ4596CBbYbo1/xYShVnyDPbbdSoyXOMNLX0yhRuF/yQ
rgwQ4+iexmrS2cXH+wUkhlX+70rBHSnFlMlHXz+iFXD/y6nXkbHpfm0nmp3u5m+QWwK0b0pCFjk2
LWYJz3bgsUQDdmf5/lKhcahmlZQEFeWOgiFxxcWPr6n/cCEohMj/eXl6TmUyHkEYBRTVx400bmkj
qif6HKKefElA1NWZvNqafsCc1UGfX8afBmBAa7FFpcNsRwsrdVP8r2jhVSBrapRAfEmP6BWSwiU+
YpbjWCG9B9rQLMdSdfoyH+SF+N5mIR717djwVUWIYVIGb4vyahvaNQJOcqD1vuCJXcsj5gabkb3s
jpuRiyk5ZFK9ywTQuU12DCGh0v+BVOgMBklNdm8SACn9zXAha7TIU35zQvkGoqYphM91EOHu+fO/
upDHD9kqIHxZa81mqI5Z0TNifWA8UYRPOVA2jkg1bNKaJnAsE66txMWcusWW4jzm+A+si1nGQGfB
ymz2tofeBuarLwf2qNf1+4ysITePzGHxyGsuyT+cihTZCoOWrjItPBuPSqY8rZDHDQFhJ0uDnV3+
ZAWyxj8RQD7OtQ4OpFMAO9pRBsbLUZqnDytXdwV7EbttFXt+ZFadxIxWPSeIVMOYhNoeSnx5DczJ
S8Yy6cRrozt3U4lkyVHdhIG3y1Mt9J0ilXbEoIHHJ9YQhpOYjfQRtZpZFtHlIKv1TSwqvTzauN+b
N9+jV+bMThkJN0Zh9SuJ+7Cj7KI15GBfZvubQ672jIb0G2+LxOc/U0ORxLlXhxmcMqHQbY/R92sD
SuXjqMZ4rGlzKdOo8/VetOQDF6aQU2vBbcuf2QAAW8vxjOPGEBPz5Bbu4EIoUovNCl//ewHTro8E
xqCabl0RzaUiIoBBdIPhQwV8eVHw3XEkWQwigDVSL/oFkWDl7L1YYuU4HrZbbEQ1qk9aLqMxloUq
64s3Iw3aSNM18i39RJUh2V/htdIdHPjydzOttHV7maqkaj/S9r+SBnFZLZHK8vVrN7Einjfn7G0j
fBrPTMR1lKJbyi+396srJu0eOelcWo2GLd9sCzsSUFaXWi1xCOeUrdhRXy0hQY2bmjRSdaVNtcZy
e4TJTy70eIyLY9c6QnEcTt0S2s0l050ezJW3IETRpGc9i3sXAXrc3ZRl+sKfXAu8GsiVmkYFAhj6
wSsz7Flg38zRp1SIc156zFF6fXq4v45jzzsAMxiW8VL63vaxHAZDW0z+pRBrFwfgU8pLsgS78BFP
uPZrKwJRCBFByUq9TLRA/x3Dnu3oyrWtaVn4T4YVme/kPkT1axvUyBNlYAkC82Cc41JkNk+1kS9Q
eBBkmCnQCeTQeJuHYVf87m2v3mQq5mDxTpndcDBJp0iy2XNRshhkCmhjqcwx6R2235VtaqxfgGma
iGmgmIgiJ82KHFyBjOTfx8mVoqVPMPpq/q6e0a6/5oI9ceRKTrVOtkOrBWoVMUvDZyxN5W8FuJdt
4ReUMZLSgHmjM0XLGI+mtj2t1Lepo71866dcgD/4zSw2yWQtmk7XpE77jmaTCZ7k8WVvH8Fj51HI
trBPvjc2GPzWfrnbTlVvekGq6h4MszuSE4UavRY81lrMGfBOCgzFeKM7RScmdP+4efjtTJTQJ7CL
w4+I4TIkyVkl56GKZIPyvBFaRjFeV6oLqXpMxbou2z1BZ41863E/7F0gMd6VgGZdB9I6O9wECloW
SgIt3xQ4+L+2OrcXzoUdV3YiBkrZ7UfkocZqDJVkGamvaXNon2Rj+XSXj8lmi/UQ4VbwbJ5h3RHA
7WXi7rxHXOPe2ZSNdvuXAvI/5MrYktZTolkGWitZJ7rKxfVL/uuNfqFjwg7OUL+zKdlAUfaWQsOZ
IZ3KSSRofolqD5ZPPWYKr4RzPPc0dzQXXE5qqVmWZ7rZkV9ddYjbWacS1FN9gq0F4ywI6oWFAqBI
Hrrtzx/jdDYwBQCMRIhRkQtBPICTv1pSFqgNwjIhzqw3bBTzzrX8fcf+k0Z590VR3bwPDzLowGgH
78x/eVCyzpZ66qFUrgC8rjrYhskspTXlwNE6CtSAOqf1uasbmCzvaxMpshyKCEf4kKg+vOr0OzKi
OfWTR6Xymgf0sZgoAhUrF48hnVHdbr8BOXsR2OMnTMXtEOtmk97Ewx0A49qFfPyCni4aYZDsf58/
x9YzskCZRPGUGRa3ticKqlSi9ujtmtFRYagsuMM2QVZJR/VT3Tkdyg4wzdA2sDoWLm6cKo/q/Z3H
18d5SZwr5/KJ+arqweHNhqqXdA8T3uHkJDZnuCFXdAuRItblmzgu4BOj14efadRahSRH3k8pF0Ra
uTxPUycFpe7vNDN0ZFvyl3baeXqoaWrxg+DErbAaulU5O/KjQgSH2R4g9PWqYTcfflsD5Z2paFbu
p4O7LlK/BRVlJlbfBuxcoBf9FM1UZdDZLs0HK6I76spuYW+XGa84FcxB6D6CV1k5UGFHxVPepJ2n
Cia7TYQEm6CEC9TKGL75PwrLfb/SfdtEJZkSth1cmRqsWJC6hK/HtVICHxfgM4MLTH9DeOU8y6Lx
p6+s2V5h8pD3t2ZvwxqPnl2DmVaKJrhufJInDigMmydnghJfweALO8XXJEjDuwxjmsXqNekLGti/
hrr+rqTBF7tBRuaf0atP10ir1ilM8Dq2UxM/Bxj7hf5Gqu0FAklvff6E5djyaRydqoin99XwjPG1
3rPUE1ntVeg3fah8YFwFKzsQ4EAy9h3PwPOvNvd+7o01S3Fs4Gm6h27d+mLOgKv8e68X4doJPGca
YDGxFmDskRl4czo1TCJ3d8mcepgdIJhFcWJiQ9oEIzmP0Ifb1MAQX7DNsRublca81OPqus21WgZy
WxlmfcW3BycV0EcyPAYC4VCEMlhEo3vNMxK4oMqZECIUvfpoOulMRRIuB4AKPbg6PMijmEoK+fZp
FVgD5MjqS2w07dnVm6BQwbR6E+Cg8B7rIiLjvYmenPZ1D0B4TzGQoYqWMpL7WrfnQ/aQOKFvCcVd
G7d/9JEk07ZUpIIri4Si5f4Ok96Z8nl5tQj/EiPeWM7lStJQ/+7pZvAyjqjlKCJ7JqfcafJ6FYjD
dH29+1VPOiM3bKcVvZ5KVyHx35lxsWijsJ752CXOrnyYl7q8Y2Si7MKc7c442YjBO/xxVo7hsCXk
fVbtA3xE2YAmLNhSeZybeiXfHncUUqX4IA5UDrVmWgiQo0v0Y1jFjQ6Lvbantg0KaiJex4ChvfAh
nionYpM5ZBN5qm1ti4lhHvkFIz6KzZ4hzvTTA/Hu241bVm4Gg+DN//ekFWdR/8+Ise1y5manN4SU
rQP/vHCOtEDbg9t9e97n4HcDbmE4w30slw6/ZnTFjmm48IpUu/L+i4N4VTzWm/41gzeiUl9GKRYk
n2tfrRjC67ocDyV14k6Ig4Kx+pL+2i02Lin4JgSaaQOJRz5kXFWYZzCJxZdEveyiHFbehPXvE1/n
bCOBF4azIg1yzo/W8Qjj1MEG55jLEVDCvFr6EBxTBaUP4nTlcUIwjSS2CQFypmd6V5CpIXMjZ39n
Caa5CeLxkzN1QI/Cnwk9IDYiBXyDiB6gmhax7DfwL7qcqV3e/iMDBzVH7C7WPhaOxN1PUw2kttyz
DLHd/7xcZmAxwfIKgNOjE5fC+b689LoHLq4ZzkP7G5Btb1gWhxT0OS7dRfsodTpyBl8OMnoro+V/
d8I+ld/dXG9+WJ//pa6I7QdROCfDtdRmYod9jwy7P4EDhSSqXLocolbg9quuecNNKiRY8LCtM8BB
gG+ByJbik9z8tgZqazXVZ0dLs6fwDs7drRN6jupC09wVszzktOPa7OHY/iYq1TsE6VCFkzT8zXio
Vt3gppIuRe+LtyQ9hZkymzQ6dLVdcA+IgRyIOrJJ+BCumMlJBj4lsuzOIyNiyZTUu1Yv5/XAAQoE
RTKqCTb9mi0X+tDEXikRwbqIbaglR/CNwEFwWtfN40KkVaKYe10G++8DP9D7jWSJ+ovJe1QSwXCq
kALWWV3uogkXaXrB9qIC2MlYsVLV4ZJ5VQaNZpu6URM7iGOOUuwxxcpu8CFAM5neZxalwHZl/TD8
aamln1bSeXdDmxu0QyogovtG2bQ2Ou7bCoFfVBTVN9cVoFqoCat1bwbkr4dGaIVO+/Sq8bF+GtXg
097L2wsYtiRJ31W9BUvgJq+BS4lwCPNkievwgkFRAoPt/oeG8zZTAdunHIYuTsLJiFcesthAmKKM
aJihLh8MK1+jNQ2Qv7CbQaw5VXO6YvKWLrqwB7zLRUhIb0uKTKFFCZxru3X7z/BkRDUVw54MKcUM
O3Ps1tBUyuX0QKRGEOI0LpVwiqo37NALJat4S2A3uGxi2RmPpIvry+IKJlEKNqE4Oxz1S0/3z53f
uikOPQ8i2gZHeG11IE1nuzmWes04UXpSTs4qRt5qXpS934C8BRZXUA0ZX3L3c5+9HxqOma/Gs9/0
Ar4Cker3ODe937JU+9691kiuKcH8HL9MLSY8Zaj/qUEv9xhsbR7Of08uRbp/i43sR7aYWPRqSQDL
LbRE01968IswflOa/41exq3mUs3Gv2UkZjhkhbbMcmc1GTuylDjw4B1O1NLuv7+8DiqRYq6afCMr
a95VYtyqaS8cpS4POxXDm6vYcy504jC6NyP0bJCEAVjBEhr23COqdwHzLPdKGroHV27bhsnjzR6D
GtYE3YGpyyg+TMPtxnXgiO+FEOGHAhvi2bNF2NFUhDPYoq3FTrywlXxqYAyGprhDccEb3qC6tp4J
qszlKYKHne8rThXhpACWAkCir1hz8ijq9SK1Lg7/qCLo9rc707Pzaz330JgGNIogD9e7yU2GBCqQ
JyFChW/COShIZrjuCLM7ez5SDX0AVXueaH4cg/ypDIqYPK4Dm+88j91V5S2tIeKdDb1OPViov9qJ
SFNo1GaN0I7alpkB6NmkS7d+zR595n0g3bsFD/Fklz1PvrzXZOvBSWnmsHMUi1FbXmHRf++5uEfH
BW/gaNMuZVRVZkl70lITsYSqr8Yc4Y1ayiRFWhVbIeThNP5eXIW44wx9yeQx1r/ptfH9mfPrEfMB
gIZQ/HQxG8MCk8r9lyPXRq02jgVb8NhAF9E1bNYBDT7f9kpk8v0Tq7k7PP50ML5Z4lKeVQ/IEDGr
Mer1qFRP0qcaT+aBXZmntEGUBF3owKCG294OwMFDFpne4TWzJNNem7YKeHSKUIBvgPdcHkrQy71E
BRdqXcW2VCyyJLAwvKeXIRt27LOUaYkDre/7CQ4S99pT6KivnDJHCzn5Cut0ij4/gERaPsbA+vmP
Z5fd3CWVNMKmr7mj9IDwJkESDFSUqq6UoWJVkHkzzMWzqnLRna/gPtnKR8eI8GqhU61ruimHng3q
ad1nwGszN99MayovgVRXLbem2h7rObrt93UkcQMcD0w01VLmUo/+5DvJYL9p4KGloXAfjWaQjT3M
/kddx3H+FAAHnIc/kSf3SE+y3BJIhjRQUrPlKJxgDXz0rzLn0SUgyRVQirdafAXn1S9kWcf5oDfR
qwq9q64/2+2vUNCj4n77AgaiGbb3tBcm35b+Jt4yEisGgRbBFSHSzSOt/x5gEiH6vThkI1nqJ+fh
ClpR0bhAn0/rLeNgsHXWzkulzLIhkChOzR3vtJqFRsFdGq1BXOQi1maisWVOoSKWudfA5eAwXmyI
9YhwCGJ6kXaqrG0vLXc+YCRM2Y1RFT0JqGsjFg3wWNXwkvtP3zzNdC8/gXcjqrEqUDu9a64516P3
kDrHo5NGP5MS8ALD/YssqJyUAlC5I+beWcGpmE1D1qPHpANbBmJr7IUgonxsqtt6fY2zu+yNECp+
Lk9aarceS/USb3mEZY3qxBrs3LGC3NQcy9uSwQmPAlbwOx7BhHSHL4mBCNEFr43gsdpC7+lJI+qb
XIm0Kk0sk2CKVPDLfN+rD6MrKpd5/52e0t+nPF/hPfHC5SLe0NtUOuPafGX/yoXVEVzGUsGIonDz
q/KuU8qU4sc1kaarupP+QK9lv0xUKWQMPPLNSUyL9KlFlEtHmH+K0gZBHjKW6aW9uICXDy2tjVad
ZDyn4i7TD+94M3lZB1PlTSh6O3l/p5FpYv7s89Lyw/Ub6/28swSe/STEQjD7hDxtQDHVwGDP4/YG
IPpihg46MmVfNfRnXrkoyviaa9pzSQfIB38xGZ7wmQhYmc4akNj38Rh/CJUQF4X7fbD52Gnj4zAG
uhvlU2W8pfk1B+oXGnKMBnIjIj/tkR7uXJ8xMMYYSImyegbKsUlJSy43V76YJ+23AS7c4w0c1fv7
OypUXH3AbEoe6YlSGXQPeryAOR0hcUuZ5nvn2sM/Uq1lHSwjqjfztmr94menSKnvGPy+PLBKKUlL
4/1hn2W/ZQjghf5KRv6lxGNzT4k/lIWfKdllYA3e6UHCk3den+Eim5jfdMaN0NIPKuz1Sn2ptDHF
kTdcTsQdIIe2xcCBW4Vh+HlUi8pu105T4XKwkFtlReRwMRPb5QQ2SrItIT43LBm0EpZbXMvqjlps
W1RFMGGwNJcilxJ2h0x4k8CcyuYcRwk560rFBjD7fmKTnmsQxvuRNFINo0rjAzy1BdaO+6KePBpx
KGIRIexKU0jlIKcx81A8k2x3s73ScfBjNrbqTqPq0Z8XCMny0lJjcD1ZkD6xXL88mxgGQzZYUCH8
CYGwBvDkR5VcTIg77tSUv5iQWrZu4mQmi0cK3UYPxUT+/dYi3L+hGsLArwUbcUhSvMNFPHcIPH6V
iTqa87I3g2s/k9bGOBSOIDG7M0QxOaY//BRoC/unvrAX7tXN/7HZy1PQQz05IfFiBcAkdaUo4wcG
79U1B4CL6RGa2mvvRJINHNdjjAJwV6+LkIigV3VjSv+WkJx2njmfMyE3KYBmq6+3MzS+PeVPAe8l
zoD5NxclFQpEF3wkx/t+oaCPSA4KiujpkJlnMnzxEKJQfzKmBrhg0VxApUWO/ekoDn9liZEytyus
gwW+kO+ExoQM1MEbbLu9xWfHylcZC15LfZprCfCJC6xgyH9kwZRQRt14n7bWuFMPBW+nXRrdCds/
IVTNnrycPjolGcT9OJiUuciqUCkasg3CEPcXwpKyMRkotAcNRDfvU4doOf6vchOwrSnNtGvWEgl3
C6NtAMpMUn1UlNBNecFFTWlkUTMhJjwR9HhCdMGrZt5o5eiLqFgMIC2gC44fkFbB58L8GJ0Skepb
uV8jdKj0hWH8G93V2//nJv0y20HT5tJwjhv/wPG6qSSlZnTttcSlpnzaDS2YRaLzhyuowCifyBJq
LNIOSYDkzdcZUqPuNkM/azLiV+98ZNeeR2BuuSNCSRYvlDTBQlkj7GzcQlApYGEPaMejbT21979I
zuU1x4gorNXNANF1A7FsYazHEivne0Ud2N2d0uzrmxG9aTsY6yswvZ6CwQK6uk6d9jB/h2c2EkN7
GvYpA7TnFX7ZnbEUu3/8LZsW2BHNdHE8Ckr7Y93tjibxskQsqGEBv2FzmuQvMW43ORBh+PsWw8PJ
hrEOaPQPLuuDyBZpWUKtz9HxHlKYJVZejoJN/6GpSK6spDSqPIYpyIsAEsygDRvPigzJ5tvcWY85
UxyiaHCyXmEL9Yf+lv01mBKMSoxhzaR7BT/yLtKEoXbcI3sPp1P2D9ZgNjbr2K+wPA4FqJnmQekg
krOP82+HxouFRC5tMHiHRX7Xb5Ov7isADMOnE8j8cFWAYAolaUYFhJNmQg4FNIvF+gjCSWGhEIS3
WvXjmyKjCQOyexdNpSRTTzEX9TPNz5lYcRE8s6DFj4g19fzIrz69wqr5Akt+f5LvyPg97RIGE0xw
E3RoEqDUlRO+XmRn7r9ZnUSu956cWOEKAAOF4lP+01zt1DSJV3fO9oozJAsG8Yjf4nEJoKTgXTwe
AJZh/xAu4V7YTn08/GZDX6icFx6apX2n0mOW9f1Szpb12VVNsd1VSQf50BaYJjSGusPe5zuN2K04
qctluF0hSUb5aChBV+F5tcHQJZtDfInIg8p+HfO8ET+eV5remlHxZ+3BIEbleYUqY/pKN5HpaMfp
2FDHmpm4YAEj59yc2GqAGSCC7Eod881lvA99K3hEPU0ObTlA61hdcXel0uBFqUCOBHntxHqlpVg0
jRKhUlUZHE0PbK0ogdO7SWbyVN2sbPGOfL3eJXd758vmKMin18pyC6UJi9/Rzlu4/GgdTik82RD+
RNkcUjBbiwgQmQEyO0dGzy2T5BduFkNU6J5/eq3g7zfIPsLmglQq7VdTx4J5EPHrkuMos5kpaTLq
PGAS08w0kxwwH3VExyydiOhDWx8uMTwjLV7hS/r836rz3cgDoLOnjMmUXCjSJZvv/0mI9R0waCkP
GZ3OO5bScqfWmxsXFOzHLcQVW+WF88p4DTOMS9+pMHRSgVwN/35zt19mmSkLiQJOSZmJcOUYnPIY
VvPaidsfRqzL9nYzfsICGdSzPzaMe94E7hTkjJXKu6jMH9LPJEucmjexFdB03cHc+xaXH5UvyUlm
MlDpL0lhgfS6lo8oesZ1w5wTkJL2Q72J6RppsvmC4F/1XV1bh8dZBv16IMQt7pi0gEt9WtF1vdV3
h90hTmU0TtZJZbRvKHB7fNV2o/6zwow+AI11t90wNXvODXx2xIU0FIQt17x5vb3zgc+oeJD9JtbH
o5zY+FqFdrYT+v81n3EZ5W3CEmt4DQm/UmFRW7RdZ9jDQwg6yoS49mDCKrWqDLWY7Bk7PCkfdepQ
ARCx6+YDydkmBuwQYaZ5SSp07P/FLCfKlrY1ZArMLTAJhc9nVO3cLPWKlUKPG8HoBNs2eQuc96XU
OQdCmgBPW4LqOyRXHaf85ktNz5OqU/JHxPTxTlbX1yfn++PqMfMfnc7+zYHvkVTCsQAerDPLwNMC
Davgovje1eAAM5bf8uaBHpb31z1ihcTa6JUpfdEG11XlesDGngmKN2pKb7oGhLP6wVMQrScSyVTY
GFMVL9zIpPM+dKfLc5y3l33Pvi2b2tcQTRnAf+WREpAeE+/L+gv6n6N26i3b0AcbxXj5QfQIeff5
KYC4yjRZX2RRMJfeMFAQLSt+bX405gH5UYUpCHlZS2O9oAaGWMmN19iXE3Sz5kbKAFIjyO9hcUWS
0zIkrea9lBT/2wcDtD2b34KYy9X9CvWveoSblXYthFHGatIyifWr2Wb1Yq96LkSWPS3y4t+2I0Vs
OTENxPfT8v/noajCI1/bYShkOlN5zjeAD5szzQuqf40tZEWePVXAAEJbKErc44DF7CYdi4dVR7dQ
pYMzVxT69UgF0khdkqN/yhupDF2MrwO0rBv8tOwN2Bq+4eaVBzD2pWt0VU/Gbiq7hRL5NIdCYrHJ
N/wD3yU7+LdnPgCecZUtvjmxhvdvp00CSMG0fXtDsfz02qkvkdFvzoqONeTJ8wvzIPFo/qAAMG75
WqoNJTevOSA88MyMKyn314Y82rvDkq1zZa4YNzo1lJjq0HTR6XvjrpslhBKqwD86Z15G1c4zAKJ6
1ZxvayIQ1L0k9BP27fKiy7pjKIooMpBApNINQiBUczbdl/K97Wn6OT8mZtWg0jhVZzQ4aqyr3JVD
MejymRFigLM6YWOQmm0x8X9pNVAsjLHCfxLOpA9wKzw3bVkefKF0zCvZArXxLL/r1PLXVB/505+/
fwlt4E0HQxMZ7hQkpb9WIG6MaxLakljRgg3SAu3Nfp5jQmL+7tm6FLeozbS98bh+Ppa8ZTxTSQpE
lNFPqiGs826wtTDx92cocVBx9HHvIo9WevPBde9FlgsQScC4VkPibk31H5UZ7eS3leBsJoZHjF4c
8Q7tO7rx6d21BaH47wfYtBKbPDtRzVrEw4VvK4CV71jjuwzWGi7j/d8op2vuQLuCFgwE6YZ8eEKt
pgWzm6OOUZ+5KtxrdFr8fdHlAUxPOZbN34joOcLzWCCQneYMKZZUMSUv/mjH3WArZcyOnhQfsA31
omGa+xaC5lR0VW4gknVnRtjbpDRPXWVbEJy8kJ3sJLAAFJ7rPjibpHhTZ5F3ij5ICCkr4VZqesdM
WdYnNLFhAvg6wVwt9O3km3UCSvFCQv/2Idoe2Iw70cmt1aD7NIbJJSEtuF1UMeHpNFOpunqfn+Us
ZXQ3xxt5muQ9L5vH017i+7DKodTNnxMS39zGq3KfJNYKQmxsJRnTxrlFevw8DEG9ghYUeMP253Ru
bvgSYW7xQoMaEjvwlb9Mv6uOMtoqukB0tsmgBi3Q1S/lNWreECykDQtwVS1uEsHdJtLEbuqQlNAo
/sT4M1Um6Bf6Hq1WsDwjQgMoAWR/RoWwvz1EpGFGl1iPNge2XdtYrUNfIEYPRmhB7j0dzTCFp8sI
qyCkN7TD3mDpd7pcgaLbhiIyA0esgPZr1OMGdbFHDUGiEQf3R+7xFtxdi7J9eHEICstNzgVbPfPs
gQDR41bXuyDJwK+FLm0jpz7c0UJ8O0oMbci35vEMEsu2zuEGLJGJ143sU+p8yuPADpbR4ivYPYWz
31d1DdEx7stvyY66SeqiEwuakBnekPtF2EpDUfLvvFi9ZJ55gVZv2ZwNa5PGvdCUeJR0W6+dCz+z
ywUDmuZ1RG3ICQAtIkm11dqLAck716brkGOyP9RxPW8NouaSRiOB2kWbQrsJ+gzwwxZykQcOosO6
DnWO4jRka7uN1gFzR/OGQAKWsfePCzB6jXnI4pcwjpLM3mIwgQg05ELds8ZkpCEFzG0HEP4ykRla
AYf22c1xyrNMIEXVYE1y/n1Sd1BTEjDi1MFAEFCWDMo8+rqMiQMYGQ8ukbwByKaz4d4orA2T1A3o
1pIWRQbI0Q0XsxTqkZC9U97vD6Mdo005uRW29u5ONLS8jtt/6jGK6fG1VCFXBhAwJARewDp7Uydg
bevrKOZAm535gczCpy9fB29ABTD3IPqnRoM8q0aBiHnkskGoUsb/gEDmxH2l7sib2QEg1iYNo5X6
kou0DuSCURxhRfXIaCsq4tcJmWLNGPjHG8G3AutcUJ6fvmvJQw8WNu7nLTaJrhPxKXrDoO67mdeR
3omiCiYg4pocWxTixO1xBMwFZDo+KSyXZeD/llcx3scme/tm25UU5sBgF/a3rbziRigDcsoIK/3Y
dDmoTusAcTeRiiEjtZROBohpwVhgOCZ/xsC2pafQYI3/aHhRurVxkOkcz5Nd+RXOzmQmRUx2Mi5Z
lqfE0VZoYySfwMQRrmshTKujX8k/HV8PNlpgK2U/CnxK/3iHVL/lZKctAoQ7bwr1Ui4vQwND/8Cp
h3de/ncmTHCOLY7MgOKKqWSbc9dg2DQ2U/bO6fvZMc71w3eUZrApg6KPSTM4OXZCBM4oClzpWSvJ
RzPWnwk7wi5YZKP9z3TGKq8A5MV5l/thoIzd0Zs/bqvFWiuMaDyu+IatLW1uCvlQISb2aE4Reg5G
j2IsidQ//i9KkH67K5O1EXI9BLNaLcLNRCf3iWgLlL1K9xfuRq3PR/VasvzsAz8c4sg0Glf51mXt
NbqDCWuw5fz5+o0e4cii/fd8Ep+Wq0TWXZPwZmLTVGSFCOyBf6JWCSlqkZoHqQyywjve9cjjEqzN
qD4hUrGzfnpUhNP5RjiJtohv8s98OOdbcTC/jObsZLTVXZEDW3HdGLwUt9ej3s2XVnTTfmQxddtV
idIPfxt/q/M+asQVJNsVdmUy/AfbmXrc1RllShpicRgz9rOmon+uLQIHXbk6JPjWJeW8PT/VXPFm
esHGSQKt5ew9k+EKzrEjGhMO+hNNvuKhoSePIfJaY0tHX7kmCxBdwMRSBppbhHzCSmO7KySD4nGS
0HSLuxfKeaRFI95AC7IR82z/QCi0lRJu+4dEiGuWAdvKbIFPN4jnu7bTXj6FU9Cvhk23gfwIYQwN
JBGa6qK6J9cyoZnhWiPtY/UglIlhHhlyL4wrCysBcAbkt0n12YUZEBeZRY1edeQG24R0cyfDQxCb
Ncd+NhpKM4c/NIfyDJ1PBIYGCu7IP/TlfZ4WZSpvyIpR/hjwlqB2lYVx5XysS5rSuhcV1UgTfHtZ
J15I2pkmRolB1pwzoOfBey8AMNFUTAzppXp7L7el+9rrRx1y9vGg3lb2DNSZvBBMWYI3vXVR5qLN
arq8UsKb1mYUbNVuve3Q+n0n5mEno1FT0xtzLXoO3swoV/OgIPsOZ1j2yPuLC5JqqJ6FH7cWj/Fg
JqYahJdzX+Qo/jYhBH7etXtwqqJtkEoaz8goFC5WNvwyEoNEpiKNzxYVlH5ukW4q2NqgZiNwk5zX
UTrBBD3LtV2CctOxbTcpJYGKQ9Un5fqOyVWNIPDvD2ZAZ/rnLz92ab81kEGQXK7hcUcSAcS416qR
RdcBEoFMWXk1qmCxPCHk04yeQDXlcr50Bt1H/VxbEYCypCkt73bMhtpOTj1nT5BQ1LDxdqKpEgvf
2OplG5FD7SyLFCzD+67pjUFzgOmmkuRs2MC1CsO2qU4Rts1qsjhV4rPCj9twQPQy/ZBdFvmtvo91
l7eviiYC8QFJvqrGXKwigi2rjomzb/tEdHDm1mieaQBwM2E4VwH5nBAGsheRJLWWdSt9UUDrrrJA
iejlhyGtLpbF63xS045xTwK6mKCCu5Nb6hAcsKX6+NCFfk23oUIRb/jT5vQXL5aTln7mSORE4OfR
VA2sMCmXNH+ZfL/M5cbHImMf1ilFU5AGlTJdmDeeKVDJUTpMka+vZck4ELDwxGTfqQ/5uAORcTZn
hRLEJcL5JoBXs6Ve9Yq/f5tKuuxJAFW58bvYP5dB0gdivDgoQahUbQB1hlxuCOy7vh8WZRPrO1Oz
Tltkg9MaRa/dE2EWy0nK3Tyg1WRfC+b5eeVbGHKpmTyJkLL9IjPilVY3I+YiLPkKlo7vhgLWgLTP
TRkbLkPT7Y/OOLYhy+zCzQWXlSG4ZT6EsdCAqzAMh7awWJNHvFoh0pYVG6r6PMZGfTxujxmS40Os
HoFkClWYnuIDy/CsWqdzKFYFsX7j4YAy2fvLR5WyFv6mDDtVFd63wMS0TyUPXE0KkRL3LSdZcHFh
jNa94X3WLEiKeNpMqeVW1FKoyF585giTfutbISyyfh9LahfUZjFUJCAwHOfpYM/nrvrbjtjhBmUU
oqi+nGhwIKhi0w/P+gqRC/GtJjWjIVSgUALRcU5CAlPKEREKKqUYN6m3o0Brk8VMXSE+mwKJKwwF
wsqIs1j/of6RTfCZe/D1Ah0EfTvDJmONt8R6Zl5372BN8SYeWDG8EinFUcFwWe5zZ8Z0Cob4k1/3
GoYjOvoYZKFLi+Q2KWUNMqwZMHHEN82VpdmpiWo6E8R0lW9Bc0eapaTQ2PnNWvh7mKx8qa14hlrG
bV7WzbM9Dtl14wNY5ccnMNGguKzrydxMsIOWZKQhfpoiF9mMLBUTUp6Cloqm0lHpbXrhijUbPhs8
Qjy/aBq+d/c+72xYcjQuZHFk0YyGJ1zYae19WemxjfTiqOv35a3ZuRPgBuXS4kb9V/PTQ4EUXp5l
qtZ/TMoOhqJW4Exfo8DUjR8Epw0YHLg38ialVR7ympam9pqA4WlkUyfzU289OtsOELynh7SdFJyt
7ZvnpTP8faT/aMuWxyDpzvNA8thLMVW2jqdnJA6nRCTptnyFJubAM2GFanoXI7BRn0K+h6jGxmpM
dvFJX0UZWeq2yXGLUoP2i20eR5U/fphS/Hw7RigiNLx9dPrsq3A3P8dGksNDGlFcbLh4hKFKV9iv
r2sxFReoXqToPqDEGg9IT9hU3DZCGVSB2a/Gds1EVS0oMYppon7n3utW1XhB9VLFOtM0VLSSUMxB
JfkHb1rGzL7iu3jwcLUynKfAzhRTTJkS/c4W3Eaii4d6+wQYv4w4Is5k9UfRYYbgpzxmdhEuLo/F
G3e1m4llyk4Vy1s2B6uspBV5iKFYsThR4kBb8vCFCGg9rm4DwpKzCQ8Psp2bBmA+irqpMLfI+O0l
Pkk0jTfFkDepgMrqTZhIgvd7OA3EuOdiNHKDogxaLmiACDWAB1R1WFvuVY9GgC5inPgr0yWYwWVx
nl0pnRnMhqp0ZGyEuKP4LUmA8fsXUELVB6oklq/aNttD0guGBY1B6C2097wIRpkgtL4bm4zHxGG4
Pdz9Yl9ySBLy9V9YY0McERJJ27sEqPm4OjbdBrVCZ734aGA9NmG0FlnOmEqU0Vt88+LqXRJ1kxdP
lb+hykVO73jR3Pi/vrmF6UgmX7d6WNcOaKfyo6UlFxcK7+O8SFPgGvMb1GMFPt3zyfxeK8YChvCF
AUb+G4Us3gb0W2cTmAd8o+NqCZJzFhxFAJ3wvHWSuJK5vnie4BHLHSD9Wkb5VZEuEi7nazm3DcUA
7zgbMQ47KLbG7Sw01gMIVEhHziHFbmeRmnXc1mehM/SYd2yXwSl7Wi/NGKFM6rzd3QU55DJFnjAE
PzRcirFQQc1rinlKTH0X7M3ADdu2MbwiQ3R2/MuaorFe23vfZAn4XsrgA4MJesSM0vgbTpe7ESA0
bRlF/Ih15P6yjScfrPtibdUnsQCM4ZLq2RgoTCs3gMBmE0COsXWwn21mGSD6boG2bJceW+UvLY0d
EatCqBgJ97hQwI3yHsIYyTiZB7VPWDxb6tc/jp12I+FgGqqSYijDdS4cRWiyqr4kpmLQOckcOnrI
O3xlVbVyIpTGqd2xVxAQb7sRdP4SR9/i26SIa5wdyDZcitwrCaGfrR/ALNRGqg06AfL/jIZwmFgK
OEHI1MjJ0xow/dK1O5AgCT/6GGZG2SPanHSsCfdsJRA6QSeHZKt4J5DM/NYWJpuBk30W4KWXcDGK
unPwB1xzGLYSh3elKWcEF+KBnK5iKfzT4Rx+qV4WAesG+cs0+fDZSZEsp0DcvdsUSs1WIStii8jo
Ewl8SuYrqx0sPW0VbyGG3buq2Hs1Oqdn8Lz4iw9x3ynJNVkbHr8JTCFQEFNmwsoMwrnKnE2MchK3
i9HLn++wiwlTRORr6JxUit7/DAVCKKRpkR7ZE7H1QUIJiKHZoxPxj1r0qUlwjdLc0Ij1Wd0jeqCu
DQjneUvViKPhySG6ovl2qH6aPEfOqiHzAriasoOSFLZIyHFo3sh6p8zVXurq6GY7NEdNqs8vBQte
5ozKpFCwDBc1fhw4OW5s6aQuNRPyQ4xAiIs5cz+1hW9P9Wu8EjXz/lVcYsjSYcUbA3MVG47E7TUK
FDngDXbA7C7Eo89hTrQhGCxiFNkd2JBIwGrTD/pkC9xls4ZoR+YzhMrtBPtYmeib0dhnCqzbnanW
XVTVgu830BMgXOokOPSm9XIwgRBb6x9B0Lj1Hnyy6YKwVYPnzuo0wbu4fpfpxDK5j4KuppVvvjDq
TFtKKoodyPaet3xqQOA/lokrNsBc7N97OxY2Ic9e8+q7hTZt785hbaqfvCbPqq2VUgLHQsCHaRIv
+npf8ORl+IjlzqpKchlgtHVhpQraBq3cbplYYTxPpfoSmpn6w/UmfqaozS2MDPNTp+0TQo8Dq70r
gjHxI36z8Kd+QDJb+9OXtUapRJ9tpADhjgMvsevR4ZqQe5tcLBG12NNr3IH3ikZWpA/tuCmrTHTX
BMulVZvW0pPJT/w6bsm1kTM5Wfm7vGvbzZRpVHOjnzWmrF6busIPgihEP2FnXEYc4aUrvV35Vzc7
YqZe75NfMp257gjPf0EzlyKdmoGnswnVnGA7lEyYKiHTK3NdmxLtvG+OThMU0I94aRD0k0+Y2hD0
ADPwApVd54a2lTllKQAAb3Kz4HjApiPsqHxVr8YsZ1KwnBw/L5gyd/Yy22rbMGnfNZJm0IbU7sEz
NIPFpqckMSUMCkq1Ced7ZeDjq2UQ3JZ9IMQO97379sFgdXejsh5ArECQl4q6zvDZzYaamlPUjYBh
+Kv2b0fwd/LpT9I73spS/gYT/pZdUw+imNk/RYQxNfr9f4IbTyeWZ5/EfTLYTC4k5WrNrh7h0T9+
PB8BLHI0b9dbKDnraN+PhIDFLOvsoj0MIJ2FVaR6TrYDVzYNVaLDNZHnxfmbloRyHo9D2W245i5M
K3oypcyNS+yWd54Gbx5TfXd25g1sna/4XsmSUPje1aDg9f4mnHGcmwIsVz6L2ngHwgAqIChHeUvr
w02Xiwoqkden9cO86IWdjcy/PKyoKdKqsP86ZJ80nmddEyl+oS3Dj+EH91xituvcLi8eroHCHUYZ
3yEoR1Gc7iVQ0IAdj7LW3+rE+sxRwI+auY4F9WeKRf+JsuqYlYg+POqb8Ld0ywivx/p/3TE3tKh3
u7TD8ZfR/BQCbZ3IrfNDoGrAwhMkIqZTl8Q127L5xzHAF3XhWeUog5UloFza6xeF2KNo4qZK/k/0
klYKIBUCoIhkEup6vF5fD4f3qRhPwiLui5v7GTjtxXduRktXNajxq6hyyIM0WRNe5OEvFP9Rxtgo
Me1DYx/qIgkcgDHKmH/FuAEvz8UnQ2+kJ5JfQwt5MOkE8+pZLgm2UPUwcr3hEdoQC2cMK97fNBPH
RjNhT+p8CaJPywy+McPw5mtM8mqjxX3rimV8tLkSdCpApP6egG8YX19bflXExnmvy9WDM3Uh2JCN
3dcXMPqRNqzqukRfMLrqk0TEaUqqzPcap307VGU/vffy16O32KxK8a8TZ06K7JYONgNDdF7QZ0m4
asUoqpIPwMs051VW6qWR0AlcLasmAMqaznYs386pzLxZdnVtWCTqLDH7XoGobpGDHkWy7hbFsY/A
8ZpxVdhWSh4AKBzOyb9ohJikq0jqmbgFvc+eMOj/nNF9fFiTcRPJ9qz8mHznbnlCcOWZJo5o8N2x
18/awYk2UbhmIwuM7EaEX5/btVEKwHLl5zU75ZrOd60mShH0TxY00EoDJ4A7k3TjaKCIia7txMam
9FNPnRL5hyU0atoAYw9y//Ff9wd5MpYKZvQE845DkOCFOcvFfr+25Wna3jivRSe+HYmieT92i2bU
bpulTn+a0aTWOExjdC1p1FvD2T26wJxpV/PcSNHz9lO3y3AzcTQVUXjDUuRatRu6cYT6bIiJZBGO
ps0MKm/egNE5+4YgmYBFAu99GwntDjPJXEDEgd7PX3a3l3XPP03eWCws9WM4QHZzCbmXlH9GUhLd
He0SbLItNGD0E8En7SWBnmh/HRVsRwaW2OFEqj731QtfAY0l91f/mYS9nW1DQu29XdyKG0O/RaoT
blAgj4T9OVjir4ox3KrIMY5fwtKYgBBvN+GT8CMwZROpo9C8o/8+K7KocwFtc79Y4losBRmmXNcp
BABegeo1sHSYt3Nm4bLrEo+fGZlQG1hbsb1zj5jdAEEYFUcY/XHfhgr72DP0WU66xoy9POE0XG7G
x/jvKQbJ7rnJt0Qy/zhs19snJVUcIom9Je74cxDt7BXnRpbi8rI0QKPIcLRU2Oat51uf/FdoS/Ma
UDIyx7CJmgGYlNnaVpoZXC2FHt2UlCubVyYUlteeDFHaJ5fhXtmVJEd8huPTSbsL99e/SvI4cImW
zkz17Thv271FfNDAJzI24C/1FgaTh9hXfdcC4jeT5XNMpIORMi7PDh81f6HkSLoCk+S7375uGH3P
Bt1rKD5T/DIJ4Acf6dbkBpH96zs1sjQyP7xa9NXPFY7jwJshMaQSaPXIlOlFnQClciT8PqrkOYNp
Oq/wM2folX/0xR5DN9YXts3ZhFG7aIEeGmLlqW0JHZAzo+KJ3B/XnQgtyurH0T2bmR42400YvybT
nd98XgdwhgHi4tUSxHQBKtfu3zTAA3o+LSsWwaHD2EXv0W7r9ZQBw03ke3eJ+Guh4SBDjvI5B7mw
3+xV9A5/+fSjyWr520ONTWVZImUicUGFuRve+qZZ6pBqkHNCR0pjmfUNI75Sp+Qb4JyP1DEe7hGt
oJ/vtp5aFbFwnCNC+MysbW6z7cJcCWh8Nyk+bn/Y84e/zYL3kcEEGw2z5WruomdIG62xZzmLUugV
X88ehyhNlFO/MBLAWl2qBBu2OkYmOEWjR2nw2I72qq9G2j2sW//Sdv+L3pEL4QjFZKDc/kAP+WxU
h6RJJ3NeJrKIu0BQ/mqlYP5CcSeMRJ/MisM0RY1cFPfa27LhFJEpc2sHhMCA76VLMrUh+5wK6JKx
0oRXHe8iEnqYLEax236kelxmherCuzWygCOVxWCVcc5gXbAIxa/Os49ClIw+gOuAzYWe68NJKXOq
fUTQdjEOTtq7uDVXmWpZ8UZEGFCItoUTuw8VfkIzdmKuFe3It0CFOGWnsJM2UZEa6VQ7ZIocy1bX
8PhT6Cu93kgHmNDN30LNJYwgopyhVLt8DIPpu8Y3nmRBxI/B/rWT3vbtAemkASeSkS+KtZ0QBM4X
m//09/yHc30OkrWrHOraaBK4EMdLWjQR9EzfBgaWMbOoKrtYwi8TCP9l4i14tJkLhzyGGWxDuCV3
w/zoCt52v+qxHSfflmdpl4vDvdoO6A9xSeE7r5evZD7QmeTJJQU6ksxbP8mrokniksMzcLGOMib1
Conj2enY5CjmoxrOx089jwwN7wyQkJK77z5OnJkUMLYQMC2SHFVprZEVtYN7ySkeimu3cyan3a4s
/ykaWsAn7MzZCJgE/P94a7iOXYE424cSkaU8Qvji3zop6LRPwHK23jsBh6vdl6Z8R1QbywjhFNws
x5d5gCmycDOYqE0XJmTDegKj2F05vThdWzVnUAV1f4YGniebDt3SccN548Y5+xRSOyKR0hsAF22s
xCGe/9heuv4m8QP++g+sJBNVhz747SPiLMFoN3XcVvMa3a20YbThZi0wWItDnWII1ZK1QcCwtxYM
wBb69o9njqwqy+CBC2P/5Zzh+9czpee6mpN72oKBD2hdc/dWbLygZAmqzW8usVdkmzsI9IdbXqhw
843C4DJZSXglnRVBi0hM8gpje+uO6cWZJJ2UckzfFsCRCToqK5e/zeSmv+qZgwTbzA6ddCoXcVjD
l58ZHrkOnRkHUEFvgGTUpg/fMABWjWQfESEbAne6H1DztlIWa52fnOTQH/Dx2ueQpQDqAL1x8umC
GHmExrC62HkgnerLgvRIU0+unPjQ0N48tEitxQH3uAv/rhZSPa+C1o02jMBijt6n2srlQEx3qd17
tylB4t8WF7+pdGSbSIbzK1cG1LBJx3YgZQ3UV65g65aeNMnl9KLZ18gcDislV6BdRDN8SMchD7/1
aDr4cGoK1NDM8FAuTwfgKKrbLYVKHnvJpTqBZIpW50rSOqf5Pxnh9R0U2lveP0I/VZSaFcXqHeFe
psPgtbStCYArgGO29YS0FTSHA+29P5qDJxxUInCWf0gISGW8JaCy4OKtzT6o8BzHSXN/p9U9ufDY
INBF0b0IvMANkzJhQYdIZSkyu2/Y7zaG9jIXT/GM64Ceh05dWDCnXkW7iRGy/23RrilSocO+Y+5c
yGu/+TsoJM2BIxdcKKkM/tn1QBtEDKlgI9lSW5QSnHyNLITn5PH7HPJii6h5kKWHlXNAuSbl+PY0
FuPCWvm3/413w2J13C5dXI5VbNcaOQ89gRQnXCuOJe3PSMypRfmMNpSKzwEkwGuKW4RCx5YVYtgB
BkUdIaaTaZt2vF1tlePqoKHpesWGfFAR7vEotH6UF/kDDS7GlQcjolT2YLZoGGey0wwLgcfTOq7Q
5hgUOsTjvIfRTtAbtdYzfJZHJGmCQ66vt4JaQqzULScheJ1p94672/YfzWn0EQGl0kc8Tt7i4YPh
/Vnn4lb0457Xfz/vFGZssBCXM/Obr/SHaF65kmxWRMniF6Xig/4NT+GsQdvJcrfta7YIr2xnXZoa
Rlf43F2sYH/UXkroXcPygP7a19BRaPmTU92yye2Wam/Zd1J6aE5hA67n/TVkRJfMyRzOIjrD8cZR
DtGxgYFIbwHsEQOtiyYukoEGbPSW/Kcyoj2NOOW61C6A/jcK+PH9gJlL5SijiPDGbn9eghrEGunL
Gq6Fber7J394XLcNAMVNyrsRM/jrvkJffvCyoUQ7gbZGM2u3DsP/Qrhstf8X0i8JCiYY8NaGO/Ws
vs8WWtncqq54FHSuTQLmJYThJVe//5klRn2h60Zli82t+dq7Bigis8+MVLObOXDLow3wyMA9knDA
e4OVyB2yvtIkNtVbmm/xvjBcWiq+XiZSvIpH4iV4AKsgSRcD4DAfzFcS7uEtxVHLeIZ6iiA78G0R
Tu4T737COP6Dz14uPz3fKAaGxsAS2mEslY26em7f47BCbNX5vcgc04X5eMB88hLIpamSjFe5i4Va
/LqzvUPx77s4eHEJG5Ui2o1XkFvc9DBRkvHHRt4AB3b9vHAjjfey1d4IDbBNBoCG+L0dJtEDFc1H
6xxG/cQGD9HBdhTyZTpQCqBxQRNY2iAQHzP8zCQpjzmGdALCi/ThUjBAIhrFtKwjXQC9q4ZtmeRr
wq3A5YuDz/R861heszrX3JAXzCMVyI7nYNQuKUEQ57t/rzzVBnY9prnwToB7n+jRGjqdilXrMYN/
vB+SLRg/NYep7sVhATnigHfXHOIG2BtIhuofnbmUtr33jHAjOZS0VJ3wMNfT5+L0irzSPVpmWMdI
cQvsv4VjBUtMGf+JOeCdGx06hRxmhvKskCdslnk7Ar/k/UbUSP2U3JwpGg7CJL8Nv7/LpfCBkKBv
fsgt0dUgBIHWaICWGuLVgg/qUNIIyjYkM2iLtC2DlEfrVYopCtZvmYF0xjh9Yvnq9G9itaQB3I7h
fMKVIzffye+jICPAysFh9L+POkAQW45pYk2aG3a3jAu5YxJhTYpWPd3x6F3cnHMaX2pTHL2wmSk7
TnZUDOy5MQJSgwkX7MQR9MVreipU5RltRCaBSPXvB2G6pJRiIB9oICCQZW3g6+s40gcLCgBgl+/x
qF4jgs0cR3ZQmmCTe3s0jgbO+d0tUwkCiT2uQVKbB4oS3OU2/a5CMfuyn6R91YeUpcNowNZzWxd0
4CMHtKnm7T4N/mPV97cgBLrQ0A1uLiEWJ4ZfbCGY5KfGWfdlsDVxsu+RB4a6GVuQX9AmyFrLy3fG
mh/k+ATIJ1oSvlPnCa1TDFUzoTPVRMoOpHaFF6r0Nh+doKVVbhxc/vTDLtmUZjtjIRMaUTEg41L4
P6LIXeYc1R2A7OVDYy0N6uaOuwAH3QwJXkLKDNhBRIRSbUXdAcM8EPVaXkFUiHCTott6Dn5+Drv1
ptNs8WOadzud1mkU+6Y11p/N+PQqbVjR7K4hGoFVl/x9nf1pQzawtkHvjumUCprOdtT5/1WXDd+y
8dOkn2Jt0TqFauhzvPiKlDWimQGpgrfA8ZRNou1kqFktxnklaC8eUCPV4f56Ebxs76b07zhHSUqc
i0sF53s/Ld99rkjZhzu1Dqi181UGEsWolDrUhhEY0RMYoEQ+z5jfnVIz/xgeea6BuwwHOTJaxveS
xP4NHK6YiqerKiGjSD0QGyv+C9zoPNBiyTojJxmL5bfXzYGDo8KHqcE33TtpPZxGiZhNbuD59sCm
grrMWrULSbvh5bBfcexiAste1i0prUd0JaKTMzjSPYM6VODh9wcsW4wIFWlqngZL1V7tOFQ/hBXV
kW4kll0+OeYb5MswM+rKaJ8zYdZ7I+Mi+vGct1dJgAwD7w4LFHYK7hpBod0zovGprfyGjYwcHlER
+SqtGup5lFU6FfoI37JzdBJsoqI0/s1hA44MA9B5mihj+L0epKoLGSHK3wubqkD4rPyesINqP57m
opz6ltdzSrUL8jzhaSrhO50C97eRJNcFdwyQ7kx7lqyFL/Y7C+Wi44V4X5Hnn23vpA1P9Q6YIh9W
pa9q+LXyePBy9f+jBbMDTwy7TQuHKRyKCtWE9dEpWm0BKYL7QdI7u/uY61ljXj/77sNYNoO8Hi+g
OAisCpGkC+hdwPJnYlV0mLt7sPHF6Ra647/ZacjbDXA88Z5oLHnT3veZiTlk7S0/9ciM9ezisk2Q
/MgEH/KqOTyzXvJ3Z7yHhhXTsFLGicZK/WcrCQ41yxtI01ig0D2vCPE9IyW+wBxHnFKIaiFwtEYs
hzYDpee6mx1Gu736TBQkPpt7jsmQFYudJaNbGJcZgKZXVE1xCmQoDHnhINwb1rla4iHnVXq7P3bt
wAjieMwSOz1aHgGVjlujbmgv7UCocOQBPcU15/Z9h+IJlvJonx2n0amjtq92pJJaQEqJ+CCjg/tZ
PueSwGcIZmE/0a1szmaki3x1xR9zTaTJ+Xfx1nrhBMZixkvUb2Jno70N/BCB5SqmBdgSdgHOQ/3T
MkLvpcUcwnw7ugJCIRBqgu6d5qRh2YfyEARQg9WDIbbg+ztGAs9p8Af8DTZvAkqnF8kUH50UBXGN
7YCAS9xio2JC5T6LBtsPzmGzwQELGHSHAWvbx/pl+ozWhhIdKDHN7n0apgvnKt/KJoGwbfOM8Xho
1NYm2TF9v6fOcH8mOLVqJvIF+tW55IBuuuH9qNCPO+WobaZnmnkC3F7nS18DhaWgTES99aJZkQUg
/oSDOeyEODQOX29elA+/nemoL8aJayDjIk0mwBlT9VMU/V3A98ugL/gt4OTXce9pQkyABTBLlTvN
Xg4h9H7Ayb2bonwEV9D9mrkTaFj3TD4E8F2CUz+tO6GD2oCTSkKNARKz82yi6zAd3JVud0ozxAcp
HGdq/rooqQ5h3seGLTDQT7gd1NcR5/W7miLW7m4fUNGwUczKgK9O7rX2SdFyKPKO8hnBlXqEaw7q
4ec0f4Ko6zSFdG9id4uWyn0pkebtdydYeBPzB7RzksoLVIaYTt2dmtBVs7z6uoU57afn7qbDv+8T
09KB2RZdAeXN8kTgkkzeIv9+BF1wXIlq7exqvqavCk4AQQg6DdMltgU4GbyDsrRHhHnLnEzURIc/
HDJbGCmRnnSPwdl5HjsqnQVn8Jmu3g1kE/ohqSoammV4+8Oi8eQs9u3E9KVbv+0YCwGLYpnjwVYg
gR5u+4vZ4AdN7nPa6/uCiOIFHvKjXdarGlxAC53hJYnlaRScPGRRDaRN5N3fKYfEhJxFn3rFN2O/
KuS1ypWrkgkNA/qv9FJzvJPg9bWWwPfFc/oGLU/bXuVLoJegOBDnuD35GTKEjDl6lTw6LeOZpZ0Y
k+d9bcBrdblKapBzBxL006yeUGfdgsD9LwzNh9hYv2VTV0ACshMT7pYUvpYV0rg9JyR4dgskUyKR
Hl6axcyZ9RTCxvs67C0CCZleeqH6Hvo9I3uoPYWeKdrXsTuNlc7e4E93VahZ2f9A4C9ktA8GbLiF
+xOASkNZDD8nTFhdv3Qch6gmHDS4PCXvIaZyDb8aDCeEn5H5E5o5bajQY8dTtyy8AY3w4ySEzH+s
2IjgVDHcy9w1ZNRsri72ddk1GyNhC0VizFS/VORSxgVHkmaVMYQ2Z2cMNBTPGvw82S63ujHbkc1H
ZMn9eLnjJ06jEQh1oTp/pusSFlqmI9cMh/GNZEImdFtCh3EzgvE4ZAB73+LuWbpG9xCFcyIOy4is
yEVgP0FuNQ0td+NTenAG5C6sBtJyeYnBmFAGnxgx0trpnx8lr9Y9CpOvITVOSX0UxgLjsD+pO3bT
jrEdNyO4+pUii9i0JHWJSmwkYstshcyVBVoh3B0mDuI/2i4XKApikD7xh4PPAG7+JFProleErV10
XqMvgDhOBPBUhsvLzzbASDPUb5lAiqYGj57I//bQP7seuudcHAs7sh9zZiBvN/HMbAPFex0q1HYH
HKtL6ZGgrR8twCY/waE2GFH3u4TL4yXXMnO0DFnGke6tB/efZ8IwFzPvCPNKsjtKqraBJ+ws+y5x
LYmTfL91U3T4WIQ9xzOTTu3r4zTgj1XsKWsnTYCLfe1Y55h6YdCDgVUGGvii4JOXboz2DA2q5U5U
o38A+F8JfOoGtZKMkyjL84gBr8VaMLDfwyzRcl/U6V0tjNbAUepH8JCL7l4DlcN8GCd/D6NYjkIo
9HDacGizvYfzpQUYorH0f4FPYE2JKi/uBncxLk3/R7bxSdlua+0BTtbfFeKsf992u6ynbTvDrx53
cju2fkVTNbYUnB+ZrW+msLvMqkAM3XLv0Z9o9iukf7JKauuS96+ApauLbc0UWiGEmjkI900LY0l6
x0G7jdbsNvyxa5AOGxpYDwQFRD1eWhQktdDW9dqYvT8YL3RgU0DlJdTb+mX4DV0COrir5TI4Ltog
RJanBCDfvvSDQTvEowRvX53ZVB+b162Hz/vlSEuibGtZY+9sWhcAleYd35NfePuZ/CZK8W/2EFW/
OwYMucjl1prwevVjuFQb42GB0XeUa6zgWM8I2j7dfbMBV64URFPuFLPO5PAKd7m5QkOK7A05v310
y7iql/D71+xATEIsYvD7zqE7PJY02VkhW5vtidCwKqGKVaJ+36bmt9zQOj6LHHvU088ZM8583MLt
69CYWyAprT1lExBKVkUx7RXRlCjiJ80EQXNy8ISJN25Yk3e36bvwKQ3GH83N2ULQ23K2UAZAvbLH
exdT0ZF0oAZp7GF++BuOp4aQZA0aH45A+36gEsLrXuclkSVfxd9OFRlqSeFMkiZDmSQVT9J/LUJp
vEAexRNNMfREYUTECNbRN/ZZhq7O3fweakLXOL9ZGOdJm8Ysj98vPwY5zm8UfxbHoi7bj2jlLX9d
2wHY6tD/inCoPEBiJvBbdNHd/Fj3TKKwrlDE0Rk4yjojq1PrG8a5xk1ZPRORQT/sOjT33KwKeeui
UZ8sFOe+c4QqfQ5gL4IIDgYtdPK1h547Nx5jBlzALmGAV3Wt6fPiuheIIF8AM3xxpyZsu0mmLUlX
TScEaTBC5CeBJkTiSK79DTOR8DNGtSuHQBOduNbPGxXigekArc5UkVjwPks5AlfRMG0B/stgxCJM
J4DEVcVGTeZCghnpg+QRs5Pi6gLs6EVSP0T6dqiVw1skcgHqsphPvOwnUGYYYuVOqN4skZGz+p6A
klL+jsA1bcOPUb1tIOnM2aGRB2RloH/DPHmLw/0svY+fo38HUUqs/Pm7ZimDKIF4DoXFqB6zIFby
n3UpTHWY35yG+s77WMJGl74CoDeKGl5WplF68eL0rRxVC0TJDboKyZLg8XSbsgC4qnGxMNC6S77p
uHhP6dSk3Yz8lV0fF/gXkNGuAUjgYTr2Jy98cbYx0U0zvsAp7FfaX+06YEPMAgg064Idu0WSaO1a
VDp26qCPYxqKZd5QMLSJi58hVZbYF5h97pN9KAGw7mqPRXMMC56L3pWEFhB3nrzMqC1LUSYpHvHJ
9OXgKhoQVcBM5cHVNkJguPGf3RFgnhrG02eNaEk6GWtd0KxOS9lhIYR2iOUz5G3MZtnCH4X1SJTu
SFHM8bZImxtfygOM/DDfARayau+xQcBApdLMuVWZEO6UdwLnhnN/LTK2CZxvaXnpmmIeVwWHH2ba
EFEI3HqQjZZzl9BWu4XqpJYMxrXVrHCElwSzi6kSIEsKPpgU3YfVrvgxoEdzxidXkKSgu1ECaqNv
vfQbENAuI2+4sVsROjHsmgGFVz4pJtMz0vJJAchKLQxJqY9FfooiylIlEUUmPM1BL7WjfMLWSfQJ
jT2gFkgTXDxt/vKSJeovIjMFIzlOIVG5jh48GUC1AfsPU+vdQ5qdU+tWyWrJhmbEJkfCNW/TIQ19
7PnAEP1x8Pn1DvDxnZgoK5pqAwmtm3bu6Z/RIk+TK0SQDrl6nvCrzwETBmtr4V70l3F0p6CjeNbC
jLWLFhEw2uPLauMZySTEPieE2VOCLIv9u6B6UKcBzuTCKuDGrlgcw+jy2qMhfW2b5lJ/AMG9fr6l
W1PAtH7PsaZwEhrdOZFZil87cNRWP8HcJocdaZVx+2FVXpvvjv99+Q313JxnO/WKMJiWbdT1mrK1
DMQhL8XMdG2AsinefjjX/PoNTcLRgdrjmU3457SC5lZqS3SI1boiEAx+80XZH08dcPy0uLkCf9SQ
Se/DpQyTLEFIFRGVc/hpBwQZr9uhP0bajQkM/RNev5CR2/42skS2XvYJbcSXoqoNHWl9uI5YlxTd
OL8+RZ8BCZux0GHOietg2/MLWZg/JE/AS3xexKIRBMfviVBhhL1rytnpxhfWCUhjscfvJTSC3S0R
cJfa5bhlZ6vz10JMQZT4URnBNyW+mUxfw8VlsTxfq7fnuyQES0jAdRvYppkGJI42DJCatCjqu3Ya
G2QT7Oihvb21yjEMcaj8yT5mMpvEAa6Y3F4eazclXq4JhvmmqZCGimjKLf8YMyQMFlCf13WKWo5e
eOOjBSjcjkHRv7QH2c2tHgedHyaaCx4N6fA/A35imfGEums6p6aQc+PbKIP/udBCObJaoITGqHzi
VS160VgjjPCg/hK8cs6aNY18kW08RzZ7rH7YV1axR5DTmV5KI59dtONN9EugFp2DbvhXlwxa3x3U
z8aXPWDuODhZmHq97UjU3pJcgH7an/pHX09Vvp5+wC0HtO2cS6ozNFOCiDVALbkx7dT5eFkneth3
ysgktyJkI1cmiV+AFQnkmtGigbN9comvD9rIcHlQTvQTz+iWjuwaOZBaZIVjBIOXxorAMEprxviq
tzgLvb5D+UTjrILquxTGHQYY7Kq0IuDgn+rWdRkkY+WaO0rfpbAY3N0DS7Fmy0XHI7ZNSPeJqE18
v2F5R7URUEzIJtPtlPsmiZdfI0MsPEXLY405fd33by0P8PP8cgOGYYeLM514g3OHZnmUIj2KKP1K
tUO+s9ge8Xuy1BRBDYnWJBs4EmwDFE+b0Y0UehoTqCVmx9AaPV2zYTu8AsVLGp856JzEHIRfl4Kf
YLgpzQz4vSZDE6W7PfKGmmQafbwOvzZKmfwMk3UepoJbDV3mSG/RlThQQW4nmYJ0hocuvseC3iXD
8HeQ63k3Sf9NvMZKYRUptixX5Wwv89UbtWrVW6w9bv+DWvdR89KRCLPy6JjRu1W3mgQ6tUvLrBpH
8YakBLxmIzX6r2VJxCS10MOMyMnEeih84+2h/8dwmi8kbfv9zDOXRiYRT0X6mGKTdihdCyBa8Rfh
4NK9+0Uh0+u0s2zSsIZyMg9XysNUg3YwilJTRiBiasmwFmiIdJmFP2Hd0pHpV9GJkMZWESP4dheC
mHMlHv+ydARrdG3kFXdpFgbQ52q2c4kaKT1j5H2u6xlN7HDXYrOib5+EwoXfEq1fMa55Brgn//Uc
Um6Ox2w1394wvDXpkcbO4lmxCVyr4I/g4XiKoIVX9JsWmYysYSfQijID+44OMd7TyJ/yCh9/W0YU
l8SeipOziO5BG2gC/VCtTadz4DtXMudYO9JVt4Oetszz6azEQgmbh9M+jF3/AiBZxfzMwNQzezdm
yM2BANVpqej5RdHWZ5XSrk9Z4eltRnej8Pd9IIf8u3ykrOrG7jUt8n1nK7fs+TDto0gNulibl1tH
uf4aNGXCg309oHPjIca7wmF9ZlwTwe4SMkBPhH4rOqUJiaeb59S9SLcUou9s+++9gTUb1EBzugjI
z4o84KwjSu+u6Dj7Bdqb8OnWuRBykUUXJHOoRH5gWIKGvsFcXRcLp5VYJFDfwDVUInWY9z9woPRf
STdaGuY0LozoxI17CVW2sMqxbz5WlAxSdjtUFVoS/X/6TRsOY9B5DVqggHANndQL4LGKZ1eFQPte
OP/bRhkcHWL7uZGMUiVjSDefZNBDybHVNlgj+E2K0Q0Jz6Ky32NLW4O8BR8q9RMFV21zMWMCXsAX
elwJB3A5wcZbTlV6dBsjCK5ApgceEosxHL/tP/pyG2t+dAL1R4W+Es953aBrih2pQyAkUTQtIcx7
OepqI4EeG2F84MYN7+hkAGZsc8RFoyzcQFWSSeio5FBkMuh/xY44cNbzAZ3gl8e/4FKNlfgDWr3g
fLrHvz0ESsIqh6rwKaN6P2xCPNaYBJdLGwVvJjfUkBWRvenzuPk/LY24Xoh3yg7wlf7X5R8V+O+A
7JhHOSYqpciscb4b+XQIWds6g19C064eIqytMs5HWkcIdP2IiHw+o0ksxmQxckQr75AV05/HpY77
jVKy0xoScUv+WJ7cnsHTjF18N4YH/3xxcjCbJRX0m1NhzgQ+aBO/AlW4EIgyUcVq0bqFYJ3NG5tU
a4Np48Rlvec7/IwWH0YuNoSW9stn/eAOwvmhR+nMZc+qvnBVQwktC8FFzrxKvRyDhx9yB/vnFQrQ
C3qfsZVWNWGbzcQKi4DzqOTPuwea0QJ6rcwQ0YoB/nWWy0f1js6zjllI6cdecKk9VMSlwLa4rb2Q
V7RdVC2b+h2ni5oXgdH10xIA9QkmQewddeUX6imKHYBT0f+CRFtQiRQ5TX2rIVJHcT8y/N8uAYM6
Xj3Pncr7SEAW4vQrIw9qKzEJRuw5ePMXBvZLEw7F9sayuoZu8BkchPKq59nWQ30G90wBF1MxjWOs
fvAP9L7ssq8ga4AJNpzMi/UN50HXVcmll/wOYiAEqRkwsBUSoI2nU24boCLfQhY/OJu8VrpWdCmQ
RkVtNPDpFNDqTysWcQXps4QMPULRhAaGdL145MSSvLAxHN7oqEWAX/zB/ucscS911YOYu+anqXUW
6QbRgK0zIj4t68hWocxyRLS4VrL1537HLnZOnIIxN/snkseOvYGBUQ7xkVOOP08iWjACZhjSJDaO
dMpdozBaZkiuwIjZowkWIuBaet3lChOR9qAkHLnq168CqREM3+mxuEUZtSdoEKKpMz0ErTWWi5Tg
WM/qThDYeiOaH6XEgq/1MYYEpxegWRPJwAquOp9nmfDzsdj0xQ/TP9WJyJkYG2lq8bwIytNkDPb1
1S5zwlL5vpbsB8DutQYaCFhtqw3JEJsliB1VJ7TExElkfh+NM/uE/IbLV2H1xesRj0N7fkbdSKIz
fz0LnceB7EuAZHqjZIu/oz9nLZwjNFDVsbykLmMuJIokTqlraQYM9ggKA9n7aS4sBsW+25wQwS6W
Q9/x7BIoAhZflmTSSC/PDstFQQ5OnNC3QmrXFwnLOGFx/GZIKrOftWLdEVpMI4/om7Tzz0cMTuZK
YUIfSw30u+lfemXJMs1EmWeyxSyezD3XGyqzpvj858kbFPUBba4k5p+JQS08T56/eyc3soV4ibMY
G9w99Ddrg6PV6+sDLdvQ6UkmkJMED4WkQdtM6Ip5jQgRcxGQW5Op/wh07CnxI18nnCKeivPtfhSR
sV8OF0nrFvDw5F5oP2wHqdCSr5t4GuEQygJfbsJQk4VapFk992/sDvcSVtQS+TWZm8cfNpIJbIlM
UEo7aVvgjoIV6gyUqsbKKumSrv+WapR7J60SDqmVy61scwbf32ofuoxn2uLaiv3vd5Fl6HgS5XgX
Lq0jhOKSKo55KWP92ryoXXJR03E8Evtk33ckLcexP4b6XgMyVFiBHwxUb1D8YGmAgwgEM7mG/lQh
cwN+M62h+VOXGbQ5RfR1Kp7yhFeZsNItlqymoB7da64Dgm0edhZsXAAZRc1Kd05yLcFQC/+9OEYu
WL4IE6mc0/pzEE31u47JVMjx0btbd4qUQQTbrqw4sJVfm0uBvWCXoQ31uGvpcr1kjia9MjQt2b1S
2cG5/52s+gNs2CG2v/4fZk5ujujTdqbGOFROlsa1Z1O086myqLdSaPCzt3dxPjoNzseCsNjvKWMY
MbYUzM+XL+lU2lJPNWW7ygtRY52IFT85wVk7ceCx/dcrvt1/Q9/17eZ34mq3QOAFNMZprYdok425
TWGKBVP/HaY/7M640EJ+fIW5xDK3ww8fjFoNgjOeUU6+eBPJBaKhJZjUNZK0zDWBWWAt6+viQjin
uEx5i+HbHkeVtpxW1idGlrQK5LtzaCth09wLNEZH8YyvbZrff7qdOr67i6SfoPzv0X0UMAdGUZtG
ftRGrO87x6w8Hy4lUyElJObkpSaAGMK+wdxAnil+fNGKBNthWfvAwGMbWUOhvY0zDlJPVHoOf3gt
4iIXXAgtYw+CDkkfItD8oSF57f/dy29dpGyJbXpUMwmSkkt42+wPlO7y2OrNW1dMUNI4/D2pSKYQ
ryStRYqEjHMg5uzD/Eoisacfs3ew2qAfRff+VRE79oV7Nu7ZECGV7FbbJTDpV1ndjbH6NKgj5tev
Osf83k8hZf3Sx4xxbocXJhQdL5RKzgG4jiiEkg59ufoUd8T1PXDrEymTr8FLyWDR3Duxe3VodX4W
nCwPzujOZOaPZTAMLK3r7ctEV1203YiiKl/acIfqHmbmVoH4WDB3ffC7uutJIJrEpy9RvxsEoEgr
tiquJkSYNZGvuZ1HCrA6m3dj1BZ8/PH5ehvHdzdX4K3o82pg2207n93k9PblLvzwbCgRJp7j27cS
wVpHQ/YbfIyIfK/4dkDAocOa2zJjiomjy0POgTrlUFnU9nJGm/SjYAmbSI9D+KhCTRogQLun884k
vDRhiL5YrXbOmtaIkjnZXbNMQsphqIsSjx7MnS18Y16WpHYlfoflp/sSJJQC9QHk5sh5Pj21UfHX
7z/JlVj5I3XETaL9HL9VlSJZw3QA99UQOzx2XB0GUJoCAhJkQtbW31c4ZxdUJmezR7a/yev1LU/A
ak46NHfs8dNHBcfm+u2ql6oja8hfjUDGBF/Ljn4dKUNmA4x73WxPaAA120tGga+nAIOfhMElj7Hz
DoetaW5bDfXbba+dgXrG3MzrMsNQ6LQKYAAWhOdMpyoGm1fyCVlVtlv+2yihEdH2VEJmt/WnHV5I
B+rWOmOumaj0QyprVgc1o0OQWg00aZ1tSpd0NHb6zr+ttRRHWcQRpCv07OsNKtmfeolUX8NIzzr0
m0zmoqADG2/Pn8QgW0anUwkC+gU7eafORdwD6RbEJvp7vpuUu3rdFyo0DSIYEFAapB1aUyg6R1zK
gnOH09eETlf0KZuLB75bKewaEHZV6a5FMvszJwQ/I+oAjqk2e9Vnbi83sZ7FywQueCO2gdikmqKr
wSV7s5gWHjg+umwdycDA9FTd6vqbf/0dFV0CprIeeLO73GP3z0nsamEbojA6bPbgzMeTpKpsFT67
XEjd3A/UDmZs3SJr/09vZRZlhIYB9gG6/ZNPd1v/u0KnZbllKgL5mydSpgIoBHERLV2oytnjtgsn
0zi/fO2Rt++6KXkKlm0IR2glDKaFjTHgoNkic5wD5QGkhWGwie+FpBvmg5Hl2ENNzhv2VJhbtgbB
Uv3oQTnbqk+9F2Odp/DaYWmSB37uWnx+rZ0VoQ2Bdt9Cg8CfI/kiNNL0idikvXH1nPE2aCriD1P1
5Pq7tocxuuFrbAVMVNZfD4JVL+sOQzmrBPPKpGI+8O7eWKHEP2uxMYfkKqbOMeBvOgVw9/reB0nQ
chlHH4Qf3BAoBU5dzu0imb8Qf3eQeSfIUUrEWnn5TGWf71HnvdVvV9TWoIqWFy07ZFMkHAxsHQtT
S/M53b3MDVdoFC9jFIgLWEGg6jzESNdb59SJMzhT938it0Z7hE23D1F19/fFi2n9s2Wqt9Cf2pnV
q7yaMLBShlr305VKrSU/k2FrP8jsz9XfFluLmIKcVabMww/FqvvIdiQ8YUIJqJuI1/mQLhV9GXaX
pXH7prD0pRPm/cgL+rhertPuytFX2iA+DH322pPe+wXRvieX/XPx1fMB9m678c/odZSWmPYLrLMO
17oT0Vpo4oohdSB1tNjwSAxsbZEYEcKClrF+tJ1CAvAiCHef/eR24yE3NqAPIJXotp0ZjeN6Kxqf
v8i5p83dkoHLrTjJa4Vc0jdj2LpCPPaXZuuKcwZyGBQEXkJIjqptDKpShdhhCplldyUVCL7ovNeN
jACmXDRdqVPIRqOYuQv4CwCGct2oUfx9gByPRPdfWEzx7mAd8RvSg7MPx9cVYT1zR/2jnDpLzoxo
8ZFOoWLN/o1i4S73LpPndc/bJesXq7gou7CIWUD4ee1twPCc5w8Exo7B41otKjqgh9LqLOL7vXVc
soHwjwxLoGFXZaDlLAnY2O7VoI+ziU9AnG5sLreABYR/VF2Frzd12SCAxkfYCMwKGcvRBQHQ5n+y
274xCrbfvckUpGGB+jwnDV7Vkzlf7WU077zxpHFSrJOsMfeQeqtZUdfn9GRAVsD46uUUn+K+Boju
Xlzlml3/ScElTBuKARh4G7TOjepruOe5W7v4i2/LQUgvbJxPX3mRdpoW+g0udGX8BCDZWZ3rarMU
tLLS8WigB+uuKdzJr7o1hZLmkNC0TG+ShXHGKTa28VeAl9q+2rGtq4ordlHJD2TCg0bVJjNz9YQX
yiGYQdVg098d09ZM++cN4Eu6QUwAUFcMaCjQ0JmxbQ905vyjEsHTz8sDgWVRrdacTPvujgl7tVXY
cmXsGr8VbMIo0ELw551kuBzStGdbVvDlL9SBDQiOdYh586YJmFfRY+0FEvNNQu7k2eX1sv8BvYti
KP5aEY/08Xjalvm+wAjyMN2IjTYkIQbzRzwT0+Mg5lZnv+t7xK5qL0d+nwAOBgsiZjSLV9ZYxFo0
U+cQ4rW/wxmi77AI/H/KD6+xjXRBskTjZoHWuL5ed11LlxcBL+CNynqj1Gfl47Fo+7laP4JarPva
xu9xDw9NhnobTY98zpq1IbNGUd7AtEbIahdaThsFaQd9xee1Jqt4kO5tgk/hihMz7xRiH9OYKbIX
b2TZOw1oJ/Te/wmY2gvV82xqKU67h7nhabXKvjrT8NSzCNqNWv4p9zorQdiMvg6TEv18kJmVDtAX
YPmC4rVxga32LdRP2HPuOunkLrbFhom4ffo2JHXZuDx/TirbIvDsZV64rY5PJQ7JJ/jqjLU+5u+j
MmwShVddq2G9jULp+xjToc9sJa02DWPIMJsc7HCWsaanE75NrVT1FWdIG93/axhbaCiJgYNjW9jx
vx9tBc/sp/Bic8PmiTkFY5cXjmlT2+qOVRxRscN34xHf9GdGauiOBWjDXd3xQrRtiQ5Pa/YFGqwO
Gg0f+WCgCVnEiUl7YsQ3/rWAHgCyguFlAreoDZBogs3Lu/kINWQK0b5Io06unG6SBK1HcpiwZi56
rnwvru/37Yba6pom2maBT4V1nxeE3QgORr31u243B8Zthb9SFCkF8mVw/ZM1sdiCQQL7cIDeApuR
ZL0gi1IQyzhSQgQ2+D1Tv0q8tC9ya5bR6LSpSUjRkXZbRsFzwFchoG4swtolNwHrNKG0/N0rybob
Ysn3AIoNUa47Hj6w+H4C5mqf8YhEgwfqdsgPecN8xvJxEIal1w8gjwmQMyMUrOiBp51YvXPawCPi
oYhGGwOxKOf7UGJVjByCZdSB+s5QlA3ZzBa2Hp4Us+xZRb9QkQururXygzQnn7OGfnP/aKZkAP01
am8oYgPZuz/1oOBXDMes+fy42GpntlmLV2A/7xqYutDzOnl1mcFDDL6sg3k/GDxJzcwA479Cxf9/
ECm1uGZ2ArL6tAh4AmDbBoaydhaZTIrVCSap6RxZ9q4LvxEFC8oHrLj0/4xXtOnwPqE5gRW79JFl
B2d6Mpi8O+Vk79fjo5uNELrGZ3sXwb2iXrsfvAClIr5hLScRzJa996NGN34HATybqhDniJCHGeBu
zpfVwHdIoRzbtMR+4WAJdVtPcwZSkukXX9AJjhpem7skICGub6cRf+tmOhWCZw9cDK3ezo2H3uSZ
9mOJZhokzP1iKt0Rfbqk9vta5qA7MJO1WmOa13PMR99W5oFryA9L4X7D1sSqYDOPf2ARorlww9Bp
u6CV4HOQ0o/T7vBsEZZPOc1og4wuDw0PbAs/YevT+EPWaaqAOqe385fF93yeQfba13TwUIuTmfZJ
y7sRYu2nisd7+q70RLLm4VOen43JQWq8oMCRJxnGDN/8Obo+y/W1OxgFbzjlR11RmnchMXTvwnI9
Pv88ZfHIuYgJKRlnA+ucnyq+xBotAKguWa1QoaM2arKQyIbQ7E/m4ymOOqPzupK1aBmsw2RpEeRB
1+thEhA+Z2V8ANRMfr+Grio/Iu6OXJJDD1kYGYnw+kV8fQS1FAo0I3VfyxC9He5V7laA21QUbRI+
Oqve53Cgm3H2iMXu4fZcF98Wi+vLPi5DCrJyz7Oo17OPXbj/1NFIHjntS9wif63H9K8bM/45rKYa
KbIbRKPwwQ5Ye/6PN1j33WHbDlrdzlQGtIHYx9Bv61EbgQY7n0g33jmn2Db5iRw5i9eEvk+S+ZNN
dZW15NFoQKVtgIS2xq1BxB2aTVsgegDh6VCyHRoNWBFCKbvebm5ySEF5RNYCMmuWBWBNRVt4Q2Pu
0XtEvLjELpWPo+3u2V0T2HBTXXULoDVMpKqh+D0zpzBkX3BIhn7qz+ONeo3GoWx8TaKrDfv6yZy+
qvA8n7j+KmXQAtH3yV23+qo1Y4kqAIchnsA5f9C5WC6w8qrmArv+GU6ucCCbjAThNcK3eefE+qzR
o+XUTHdlCjg2Qww/o6xz402ZNBNv7PVSngp4ROHtjfXceUtWi7Yh84n98R9S9Q3cQdw2WwEEoixm
C+LsDPWY2RB/90NCNDhWo8thqn56fkB9WUZo6lyTD3kcR8FeOpifs71D4Fj6bQJDBON6OZtKKfks
+qezW44rG5HVnoiauuAngA2LnTIjt6HvoHeoOmbq4HRJ1m/F8Q9dj2NSCQ9LrmU13vyUC3aYqHJU
cHMLvA/QUH44ESnMwyZilixAkFUT6hSVBEgbwxYy+j68M6PSEkKWuUy10wRJgNte42GRkXtsWVR9
5Le0LmDeTcpWUVp7xdHxuJOCq+IJcWOWVZRJKxoncnkSwy7pxnmKwTNEYzW+PWtV5VLADa+grB53
Rkdidfxqe19SK+gnrcD96iSyzxlaFR/aAqy83uVGdIciE2zN9vq7Yvj3EfuGX+3R7Bxdtusg26sQ
U/nrnMneDLlQqO+idJ10wyOfALCNQ7nYtwJWzBbaATiFsUUj4yftvvP8YY5ASJf357vGMInOsSid
vRelwzu1MruTUugFZML4Yc8ct4kYIiGOj67mQCSuf3eNzYWy6uF1tbufB3DBN3nd4KWlmKAynEgl
AvukP3WkLsviqLr+vbe/ON2U6E4ekBievC7YWxELS4WR6s2LjEDnqKbsWOOY0Lk2xLiGRUa6ioD6
BcYd/+Xze4MTz62R/6xcjE4iakl7i4QLYl1/jGoQf+/+biCuJqHGjf4CLZSkqc7Dqkr/+g3+/M9m
ffSEQtNMhMj5NPsBtNtIWZm4yWVi+KhQZzVirgtCd3NMQ3rRIUMYJB4HbnA37j7XRvcx2inAWhdm
kw6sh2BaTKUrZkmEvcnsDn5aW1bawUAJxL35ipxnVxl501SUENcN4mcBTyXIAileut1nuHNMSOLy
iQmsX/cSEhwWur9YreHFhm0kiEKCFkB6whIlmCtDOEVDl0f/k7xwc13nUhfknMUoDYsMVHOwQzUU
HXAvPgadT84b2I9XvldMdKURZ87swYV+FTW4zBdkg7tbTznXLSCiwxjnQ3qTGwVJzGAzfSe5kXAE
wwqTU4n9dgVWNlZZxpsV7E5jiG6nCh4j+58fUvVtTMl4zz1CUXDIv7bDlIQWCvsiCKZBk3Uj8eMS
mngusJl7Ez8giff7n2K8VcC5V0+XMDsHiRVuH7mK/5U9vpehsOJkYwP4MHgesX3Py7Yxyg0wThbC
HTSgIGrE1auQ4+g13jnoXNUvPjW55DAhGDKrxrHM/yErvThD3tfM0AkJhEtqs23ZXfKI4mVly5kg
HKxNwLk+jdDLdwhQy52sI9QNilJsgoIj9azDVj5tri3odl0GTrLuO1iKM6AohjQpwzL1OGDkpQ7b
ll8NVAUDUWUNIE/m6kKL/uOzCW8M/75Yx5xtPIXwmz6k9r42lTFznmItLSv9QrFgQRMlEaqFduvF
ywO142+wwyYM/IHsfjdpYvROjELPtmEqUWJKK3s2DnsQUXTrzlvk9H4AHkXotobOQZl2EewS6QFg
opA79nqj8LXanuaJEQBZYIF/A40rekmERQRir3ldZmtY6MOQnPbuucVBz5N22slNZiA066hrecmQ
R5ABpPeeTP/gaHg2w5/JZFvfAIi5gZPt1cbofVHxy7E4mz/4DCkzBOMZNdRjP1iBLeN/ZJ3AmLKQ
uuRbEAhC+tXhiXJ0amJp/6jfPhNjBHyDkJ15LfyXkOCn1t2vHi5r8AXFVZFwsc4cZuGybj9wTh1E
9nTD+QSbLYZR+Aov741855iq8BH4mitS5CqCbadpOvopsDZ1tNLrTXlUbvUQiVjD6SZ2THfv8kan
IoTLKZqwYBF2dc2XVW4oPymnWWcphP+YBUSBatkmwtR6MBOEhzdUdL4F8fyVujgEyuaadipjOx95
d480SzKtBR6yDK/kbkLTFtkaUcBekJnJ6Jiy1XKs0QmBHvJBybeFGFyey6oldBsUEJSG8H/mpjDU
7pXO3uryC68Rl/oAnllYjE1s/nCubBCfvJpueYDqvQTmBMNUHcHaSTMrJCwKBm9FXygIcEdblMJ8
55JEbjx2qgyiErs0Q2Q4L4XMvMnhI/FEFwCOlIt0dxr0/X/KYAMZV4RngO45QLUUX0mlZlCwSyLW
F81prBuVGKf1r5cLe0nk6nVF/6HuOdU4gqA18yxmUxVk5GJt6/7Bc8qy2dvqtWeBfU3C0mGAk6Qo
anddoSzkDjAAyiKEPEiAZMlSWgmahOl+/KV6OLffKdnfO//sUiy9OlKKdRr3vSfSeTnsRw4dYJs8
PVgzSOpK27qEjPN0aabfwxM4mJSR7JZO5WIcfMUaMkH0KEpT8D/L6ZiPekGBUYlZNUsT31HyFu2B
DjrajpPtbWdSWAI6RqPoxQzIdixE6Ml1lRAva1FlGQdzCcst8ty1bQi1msYHBCtCfCUxrLioQRPh
J9NNY7S1eMyJkkZHB8otXjj4aCCgiVhNb39gO2AGtojnfVtPhlgeJej82vtghY8ZKSUj826x2uz8
gAvjFYH0n6K1qNvVkKcTxo1jv5tPtfXdWeCiOqSvUOZCqup8/6/FZdAXSpjS7cZbQCStlrVJjVD4
wMwJKDsrTLmTywKuTDU2rdo6T0DjFvU2tR8mRHbRoBVgJC+aeZ20T7AyOe/fjEE2dcI0JdUUHdO5
5zKO6nw2ixy2rK6EApWeF2nob3U4ZtshCjSuakuCCwt3wOSwuP9eLQ/OrGhPNPiMlqNz2/s4EBO/
uAzr34rPXdgwujOpY+3Ztkj4UuL5AU3meAwnUAQ/l5jlhf5Q1vApf458Wi0WunhYWfpsiJIrtPHo
Sfrs+At2Dh2zYwO5myXR29nRjcqY+i6T4DK2hHa/F0ziKYCNgQ017MM4Za/jhEbEl21QXdZpotVV
LNizXzspbYiqgF1Tww2cR3GHsPYLGo+A8ZV07wK+/EVoJ5oNB5ntSOdl08DFaA3hs4/5/uuLC5Fw
S1KvAwN+s1PBsnTIpdaMdF0hA0JpVdFm585KVgyzxe5FBKffP8uiXX0UdghBVFuStMlna7ssk8Iu
MwkPVysp4L29n5bbMgwsHw3HYGRN2iM9ssYUE6XshElaG4CW2dFQOZgnq4Ve7ZJANBpgUTO+qBal
KaEs0WGD9N4Nc7Zx0t9+81hWqGpu7U/U4ezBbMnNlNFpRH870Yia09MtqBi+RbqSavzXBA7om0pJ
WwyrmblgzZOTmyu6Gtp3gPi1+jwMLMbnLnPgRWY1nn/LtrM9ySWPqpv0codxlKGvbg+AdDgf/C7L
Ncta2s7dQmj7vOk2TxFM486Vt1NyTKwQePuKm87kZejEzc70IyBOJAfwycFfM63Wj7o9ZTb3Gw2F
/kWNhFWWJe7AiXhGjrAes9e2oBxu+VePX8goII+LdikMVJFBCcvyKGTJnfFq4UxfF05bSTG8q0S0
QFrE/bj7b5ULot0+ltpxZ07MnEdRyDiZCMsZKk0NEKEd1lHL+GEKu8bVqmZdzJFhdF2yHni9R0Mq
nXIVSHMgMTfEHveVqym5y999NDpnETKJ8JI1IL0QYersjIoQL28DshEx7sqGlq3LEGJ0IcL4/Mt/
naWCCpOvCW3vuqjjdVMCLvKk9Ik/TpVWnz+1MC0tpSsAXhxhivl6dQ34CPFsadeUs1B8VDkDi1xk
/kPoKGRCQUrCn7SgzwTixC4WgtbabrN7qvKC8T70vLOulNg6DAap5pU7BZ/6dGNI8Ft3UoVDuLhG
Pd1tLSPWDVpoZ6NzM4phxn9dQIaQzdKb77MbPd2H4+hnMHZ3+e91XNpjFrLo9qqVISgZGKjtqcph
HTOMPc4S2mIClemP83V77jGJXIRfEtyZeg02NEK7w7ebhKbKHz2MYjw0b9KnsLwCxpmnSKJbxVhK
qZbCzX9Ryk9RX9yiRovFiU+d077Y6tlz63sxfUPFW6SJZrvUKUTYb3gbJLgOr4UCx1VxgSrcBJhO
Ee38WR6d92UaDMBZIgIAQjvJHG/AQ/n3xGbI9kH8hD2MlghCbGyXzbyY7kBR+Qu2kyJCBOBdiewS
knA1DKzMXKfElPc7wNbYfhrPE19ms71ribidi3Lof3rA/IqUdROv++UM7exNhacORZuSNna7fR05
A9aQMxOPGYU48xEpKcLwqLVoMN/BRSbzlImRst7L5hZN/QVRZKpn2xxddL2KNdc2MD3wnrEH2/I1
M274oz8OxQgQdqkDBKOToux8pBkNOahuHsdgrpigCZZ+l5DNtLsFYBuLpxvKsFZQAntzCYZrSxkl
viO55iVlwqWCB27YPYu/tylT4cMavIirtNeAU8RekMjdL2SiJpk5SgYLBySWSP5CogPuc9L/AcKn
wmXuMbs2FI2uoJallfGZRjP4Ja1NC2lOGJ9Weqi4WQm2lMn9wAc6J9f6ibwCwE9ZZAOHhFz7GXMc
YCQkNb+VSZ2r1YwTpIq8X+NvkWpS79cotPH20g+kyHsmcJQZX6hEW7D1FrCAfKI4tNCmNfQVdJH8
Yx7ooU4k/gUl2R8ZRRX3mcMgAa1EMkZqhVa8Q5HwFbYLW2DlmYVw1Qhz1h9Ogm8hIV+HkqgOZhcR
NMDqqls4UaBMH5BtBKc0MFMMoqpQmIwOqpOny5i/lkEvNdLLO91CHVJ6iZqcZNdxCc8PuuPahA0u
CeQ8u3lTK049SWZuP596SywqEXZ9HxvSDrra+3IbcmWEylEGsHPeRm5TOMX1awGzLg7KDH4DU+Gr
33H6OsxR/gzQZmqJMDF66l5Qk760x7gVI2wnw9yA6DBRXTB+SjTiAF672JMoMJ+QCcFu1swpETqi
GFIbfEXHWSUeFZFEQhyporhVDzRd/3xOQS9wrEV7SidTyAZDlGxNJD4xkDYotN03S5mo8CjOWlOl
YBjy53baO0z2DIsg58p4iOA3LboKrfFlp9ROuUGXmoLWwkhoGSZ2OLYF8zRSv9pSRrl0QszoOEDQ
qFi6/msf7zqC/JUpII3LTjZjahM+NI4tePgcWvsrLzhXa1RpzWBNUeMFRpUof2UKhs2tXg9AK979
BS8VlpABuSOXbjQJud0mKecChF3UmZXoP7eibP1tu0bCLr4oIBu4GfFjj6He5lSpIo7/AVDZ0Jji
MV/erhzuOOqSrAjtrgP9xcj7NvELCLDzb+1OgcghenNgPmNFFf/g0uoPVy5l6UvxuvniUmrYyVAH
pT60Kta15ZqugLVzWuEMVGO/0fiuwgcggOJtPe3ppJkyLUvHutu5MLcYW3jX3WfiMMZ7R5eu7NiE
rFwvXcBrcNvUh8wk4TcVFX/zzaRWlMSEHsAbUfe5Q+NvFLuexqH04zoT5B/ySc/cYIFeULmyt8GJ
DwEUa1vF/61/zkXO2PBfE8PGNTisiMQN/SRiE8V1U1kSs+/S1UxUqWpOB6MXrLmdk+kYz6FdSuGD
0eNjZMe3CsA1P4W6E0zyaaK59Q1Z6JiMaBPnf1hej02W41oPtj6Esxf+weLAGzP3nyQf7dnfTHrF
3FhYl/OvsrWOot+meSzMzyHKepTVwBgoHNekwJm3NOPF8tDBkRweXvYrjzPqE4YjTFRNYSBXl+ro
e4ua82aCDZ94Q3Zw1ED2VsOS0kGj5TVyj4QEwxMU7qOrInjJVNCrnEO48voumtNxFREjxGTXEMbV
+IIIVi2c0iOfN8nklaxeYF7LXWfWHQQGTWiLZl4BGTpf7q3+In8SzLRPqgfR0gpdaChtT3QYjadl
miVI78QFWUPjua1Ufz+8RnVnkRDRK4w+5F9sC4DOz/hjj1hssFXR3YnnTZgAjqzmUFdppCi4zsDV
fXVIMdDVPzOYTYOmKfptuKN4AHSXkKyFYpIiVDN5beQRgvba9zM11qbzaJgl8mIgXMwA0XLPyidp
A4DY5/qLPRjtQQS747gCIYOH125i/IJvHA83L24MgITf/bvP/UVLfOdRbnlYE5gvA2tCa8eeIK4x
d4yDLg4AUqh+8OZoc0JdE5Yn7VNPnhE6QFd1iwCzuVfQ4MTOhrtjcxisFC/SCn1395IHoyYnflfp
OTdS2HOkoicmTgG0llaDCTlRHghGZ+dmaj4chm64dr5Y0y1uA64VNoFndLY6K08VsH9FwJsCKfHr
vSJIio/lEtQjK+WJk2sb/Im0epuSxwBi9u2155SSKg+0Xfqu+8aHF6/T5ikZV2Rs7E0c6V9X8UEK
6S3zasdiwEw3XuuiNNq/rtEmkTfRhNUzOpJ/jOBGhpE7Xe/snoSD5HR2g8f8tTY0ORi9vlaADDHe
7Xq4n8CFG15QNfZflMfV8lLGu+izmPMiLWlOQX1aPm2hSCz/Mwcz3R2VvnbZ4jfA9Rcl4MPNWgcy
dUjYCdtSoIM6vPhF6BoceN9NIeOegPj2ObIsPb54ky7gSSE4HolPkOEnCBYsNgpmYiwPfJAfohRy
5o+4FDI+M9LB6GI+U1viCH9DzrudnTTGkCvyHSyLHNNrrWsVdSZw8vIMEDfRpxqA8/fJ/S3tUJif
JK0ejc+6iGR8K/dLpOxwJXuB3rYE662GBGSExfFFS3AKOpuYnlQcohfRubD53l+riIXtxn3/pZtt
SfJ/yM/PIyIReuXRHyEnS1quYCPhRvB5iXGNnDIEC3+sVnJJ4tPZ0XzUQFevlfhKMLlM7BdQcJRU
P5OtA3bNnTFZYhNtQahLYiSGsVi/ELPI9F75TZPFHPGqYnyzamYlvL0ryt4e0DO/PygBkUlK1kRc
Z+c9VzlWDrTqRhOYBeU6yX9zPe1NeJ3HCkmdm7ix+4q1sO5TAL5mwg8V+vmeTn2EzkkDtaXrOq1W
dqNlIY4POXa/91b4VCHAV7Y59qwH5oAQVUzv46+vAvXMcBYGjlsYVsqjCwI61Wde36RAeNIkCa74
ixYXaA5i1RCzpJE9c/qZV/aU9KPE8uJ4Fc6P7t56mmDzfUZ4De+4Btf2SuFp98Xsu51DxGfBBi3L
PGkQLom51v9UxdGykZ7M79Xp0euialhMOKR0Eca6ZqRZSH0jl8vghKZ7FvisxyO3uMTWszOiEl8Q
wcRvyD41pwyDDJzKdEErADLuyJ71GdtY5qdHm5chlKKWjLZ4S3gKcBtTdt5OQdK9+NFPuotH5ewp
nAsNfMWFI+J6Kj1xWpOss5AS5Yo+FAz/TVR9yRBoT2zUFpGNmyFeCjLjpDZINSQ4Aexunp9LeHMH
/RlBOtquF9RiRZVq2NsOeWAc2zo+JNMgjpjIqpgB0USbs5R4PbkIRNjHsylPCWx7kpXfX/g9MQlI
7HOHWe3W7So8jZPHYVIGCprAtWgDWXa3U3C5UfOl60gUmos9iSyr1qHO8CmfKaxmfUfSnNh14fwm
EkOYup3UyQW0pa3Z6u49yT1281V4HDAHV2MQSg/x9OmW/E+EiqQux4WxMpkAWtmpGrOq1pnQJ7AJ
q8XSE5j6pBLxuS1y/nx696UgoXIw3YlMxLOIB2t8Xg+D1myrFvga3QRWzxbnsW9uItR0/rYNkDGV
n05TFyKXBjDBKv2DXD+KZ5vM4FtMA3XTQA/HOqetYEtR4tNAzeXLKjJ77E841dd3+g6ozqDEe4m6
AFRInNWPRQZyfcL+clwB8o8JUKggGARU24XkpsV0DZQjQcmMv4dN96DaH+BVjlB2GxyEAzOq1LFQ
ssDucAgwtSZbJGEsXIY2z3ftxmXJj8ef0o8v86DYf9hSipGD/iNbzrt2PBmXGpWT+N1ny3xYfmaD
4P4IknhtIGJ7xH9i5MNLyWrqLtzAAzAmioX6GOs/vgHh8MFysFz3pGYNLKzfFWfvjcwi9qtmz0UB
rMpctr3ezbUKmvvDK4WfbvyS8Ugi3lL5SsRqjyRCV3seGUgeO7VSGU60bYjOKvOl2y9Uu9b6Badd
5I0r0RUXf8KzGTJuWKo4wjR8G0XM3hL7NXVNX4GW1R4HvJ4wXmEEBgIzvwpKz84rW2GXGVfD6ha5
JaBoclbTR/Fi23ivoeww9QVidtXC4Q68rCEwSuhzljSQyAeJloGn6yWVzCLckQN1OauzVY9JBrDM
/UvFnChcJRAEZBy/Leo8MBcW6M1RtXI8dV9HgtivaVdskKXJboDY17jo++CmBDSxAsEJYTies83k
T00sZ1rdmMw+uv++Dv3AdZCjvm2v1LSNpw1IZ+Jv74ZwpFgtfHFJ1XS5JrDSlux38kICmpS10qF+
Nw0cdsAI0rX2kd/r0bZekbGSTK42eCsfMrlsSb9mB7+UmsQfeUe+OlJ/q7Id65fhi6nt/Qh5SUFS
apdGttJe5ExePOEkHKQe2ag23xofRDWpHbYeFHpgnWvDFhws1ITqOyh4QKFFqT4WmwvTt7zXcDlW
fNW+yWSyFwDVopv8u2zb4v4kBcTu5lutbEZuht7VqNFDHHex8a74tk3evHPUeziv+tRJIwaGeI+b
G5APmiH5gfD6VVvvNsYk8qTkFlIT1XO3mTfzjY6s33t+M82NCJpIySB3Xdn/+kxxI3NWQfld17M0
CPDdVqkKl+0hQi9r2MStxXvpkTyg75bW++t+EKgvahKYg3fDX4k8yM0HT0Mj8j64vU3O3wARxT61
3SjpEy/FoKhLbVxdnuKTO3gUrYbxP3+L1e6HJvbq0AWV3DUpqRyOEsAjZolYYHR2L9qJ9ihNatTG
0W68gZWI8rI/ZjCdIgV60iRO59G0J+PP18NxRpGjAaEm89ieghIX1hw5HLLjop1x9Jsa4Uf3n1s+
f97ChDbYdEutJhGspnzupxS0vH7JrDP1ctk3xqAqlomnhbBT4AqkAW5ro9VWxmdRXcWBj2nQ1xnf
rFLADfThOi7vymB4mTzifyYNsCr1F4XD3bXFqGKU4TeMQ4FHWr+JZvUAaIAis15Mm20T9xSlHaBm
Vk+G8Tc6wZARyaOBx3Q0M0K2iDwZmsxTJHoyHDH/A8n5cYuHzs1zmL/CxhPWKe+XLMhmCnICv+6u
ilNV/JieqxIKN+/2B5d3CD2/89TWtJ/s1F7yCUCMVUbqb6rfPag55vQXdZ8uQ4wdMHn8/zgpJOgO
1DDoCdh4aiH2mZuVk4H00bO5iMEz+LvojYpmzSVFTqD9nyWQktcwqzdq/200uf9cZeReg7tim40i
guWFgulbg4Gb1EV7wwUrqkqCzuEplccGU659XeAs813746wufsuT+Hqwd0/IHr0lN2RWgwvRE8AF
2da/1DHQZDPAWPyfDGexU6uKFvf6GJiVwC05YFdXgta8whgi3zu/uw8gs8yOyT0QP8Ktz6El1wbJ
LJWdE5Z+/BBzZziV2s8bgNo9msxBHaMBMgLJEWG10GxS85pIVo7nxGNOXvOju83IgLUi+IqaAA2u
hkqCCQu7zEellXAzs2tYdwZkPM92bn0f9yJNC7kUAT1fJdO+KAbTTP/ULv2vwTv4/yoUHXFFAbAK
G5LUUtYivCKtz8FPbA2iTx7RUCCP7z1K3UDn6XIGvuwhEB9ZEPOZmbI/en//H0NhMpXht8QNLr9V
N5PZB1H3lzKR1W/v19orDrkkDkCGjWZD4FDS19rp+8SC5Sh98wC8LLlkKnjqQTu6aej3fvPO71QF
GtrYMfYn2SUK0qPo8kByfeOYurg3YhDqsmnn5JY3MSigjfNw3nz8o8SUJD5th3WuzFu34KjagvvK
oth43SlivN9hpLZORq5oZepJfnZ0+a8xiVpv8O71UFpPTgYAN11H6LZLL7Id0Q0B7AvR7Xd998Tq
zDWCUft6A99ue0jUqSQxlKlja4gh+mN7xeelC6oDyu+9stOVltdKB2SjpRGKKG5auqmlEoC/VCle
/+MpRLYcSLspJRApIJsQ6XfknJWTnPLbS9t8BhfiI9zylywkZFZgfl9/UQL/OZqSsIFecuA1CaPA
RaYtG/aWi++jVyTb1HKQy2y+5dEEScCurSmfioV9kYDDPcR1Vgql5gzzcI0GVYxK/rdk8TMiNUY5
zHUR5Pbfu3udgj2DeAWDq/CzC33IFVpMUJb1nd4HpnkVunayvwYlG7vE/9ardGPJIDMU46HzOqiQ
KwJnM7meQ275+SqYrEZEsOqycGzT2KdDpuEszLBeXHtee2R8KHOc4JAJ9+VeLPldXOPkAM7PEugC
XzkUFHk+rzeQ/w76x0KxrfTzlWuj0SRxFCD931PNrTu8RbD55+JyRZGwtGW1hJM3C+Qt1ME8aZqd
bsoT3x5MEzbjHLT3WUp+VxV3QmszY4VldrBvESDLNnjvyUBqM1otp/vTkktn8E/dgJwWie4CyoIa
09dm/BMXbMb8VaK+EWYEqQxyqXbFtAdFbW7xBlUlg2rNWrZeyPIuV12WSIfsomt39wgzaXnMApxM
SLlLAz9U+GNDCfNeOqW31cxhC3i4Z62UL2/jMRsWfwN3NZRlUdX71jEQK4AIidOBU4SoFnRwRZ8y
w8aDw9tBdnTXILmXpy29ieDAePtG50a9KKTsK7r0qf6msqiZslGdPu8J/cbM32m2OS9wuWF7Bo9K
QxhxE+mv7CdssIQs2/DkAbAxj5l1GTfLRZRyizXJCMLGQwPNOQXUgphYNl3KUJEKNmcig3x5GVkw
diDl11BryfUcynG8XG4dH2t+JHn72o8JfflvOU5LA8oE2h/Du16Ah20OkHroWjz+LJAhqtvqOFH2
OKVnZ8ECqnvphIIwdNwawlIvxIhV64XAqH+Don/pegbKL5DwJQR8v8fO1Dsrns6iPJRKjMu216gX
gh7IaERvfXkESgclvhaBBXmMY7qMv6mER/9cl9Z/Tr51JngaYYhkm3xKlWZ4MOmFueXAcJoE5ZAc
EIkq3vnt6caOGnZupsZTFUY0CgeTNSukVaxzdfCjAPoiYvz0iihlo1NLSGNjv3I09144KCJ7O0jb
RIGy8CEbjIjex7r4mJ6YHg0oWugp+NGoPJHgeMq37KjoW0MaQAk1szvSSv68GyT0Xz2DeLe6xdBE
8LkhR2w+JYd3Jr7opB2A4smLPSdxDaIy+LcysFta4SylzK5Y9kGNtC4ICr6T/9xf+OIrFWlfEUO6
wHFmY3q22TvKWEHgKgw72Qis9/h3bjfzITuUJRGEO14/1FHRSUuU1YiaZ6wLJjgrvGOo3Rlid5zM
P7RRp767gQ+ttiwhclmZOd64n2xmt+m+TeYZrSb6zFhYtUn+az14FvP3LSBIQX9VeA6f5X8oZR1Z
ploiXjGw0WoJ84ROhbWTwINWddUwknvAV6ZMU+P1sCehqzIRB55odlxVdKT+PC5ep821iGrOYmmn
CxbTilIAifcvQVpbDKWu/Aiy3it83ompG6hsRnV05OZOeNU3nbCIyZ8BGP4dfmMcaSSeq4ApVkRx
TInoCVmdBJc/mfdmdBaGY2f7eQtNmreXqXgcAdNwNIjKvGPv4MQRqDu3G6xM5+sOTF2Cm/FWrW2O
TWLa4SsHUlIZbJa6dwDh7dNycB+OomT+np+/z2yZ45Ax8D3eqxvrjdXwZWsEbhuJ8l6yZZMlbZuy
D3keVc30GPNwtwonQc5fPr87u+O50TevRPHgcaF/fYQ4ENmqGHlyXbSyOpdFqM7ePWh0K9Tss0CJ
zCshVgperl9fYrPhEStZvmbc2RMzAnvGPTwrfF9Kg6SqMw8969Dt1S8TI+S9ScztQWSNVVAEV5py
z1ccDMqFtev+FNLCp4x692dBKFYdFBCwLgLLqkCscyZORFNQ7zQB2VsI7kH8TqEIU2mJSXJC+Kbm
Ztr6h4Dg6i8m1bFJR5JmbJkES9kYJaBgOftx3ov6iVmcbl6kdVsWplSiWUo6pCsnxIF7I6Y11ZHy
D4gfXWRC0JuBCIbRYE4a2H6Q1eCPBhsLG2twPsZATQRGLD+Qr8/nn7usGxng6DjRjkELmB+//z96
xKAaxQpAxOLwIGmynqWWUz4uxhIwvCkQkoRXmDtN+RHZRZsG6O4V6wY1IiBG8finS7vvCRCbovj8
+3JmR1ZBMLgYPTpmY3cqq8QxMq6X98JafuyM86RlPfxvj5JzCi5QdMwWIeIk0y7kh3ukctgN5qLt
ht/zDwLx2vj0btG6ulQ0nOWY3SwOZRpNYAZ4zh3CyZvLX+Jx0YECSNderwLrvZsOPFZttWNx9EIo
pjlKhLXa3wXS3RUN0RVUXHRQ4Kisif/k9jrMFEwauwXkntKIjVjjcxGAYLbl0neYEHpk97LRapJk
gaFgCA4hdg8Winj4gaaeF5ccht7C7rKfl+VOMssd+ogsUwxAHaBoXEJDctJSbs9YcDf1n9JBlOPY
G8/IwOD0GZtjOedIYOhcv5hmNyUENVhCpFzJbSO2iFW9jkxz9h0bT9cDNRQqsKauavCwyx7wxnVq
p2w5Qkv3fJhU1i9X9AhLAWXrAauc/JyaZ2kYucS3YqVd9lZaDD+rIgouwu49dEl0IOlPeU9CyrPu
kga0178gw5ZtZykAer3uG2e12u/I22UvALVYb9Roru7mUs7eGIE4mpvSTXTtUgXupF08MM7jB8BQ
m4jsqKVCnBzIthM2vT2aTHhozLxweMLcRuWP3C6G/9xyGcD5AGtctPMf8TEm5T71vCshPQXdWNAH
JwpH0ttcpvUKzhLNe6Tnb/raB/LU1n+EKlROjjl2aW2OoCKyoXJguUCmlkmqAznJJ/gdaEA8AYzb
XKQ2P8vi0WGH9EevZKT1v2j+eHVln7cW1OG7vuGORM2dh2YkWD7J4Glh31ZR0Lv2el8rkSngb7uT
EbzpfcHRIYqMnTnti5pyqHWj/Dkx+0Fto2E05ftHW9xiz0bBl0HNyISAlMjXQaSHrQ5mgcc/0Od/
9/AwZ+HcRN7RGWO+O8yaezL3b2hGMDFKzQa2uk8U5JaC7xmSsVv0WKqDIZG94nyDl79wx+vCPOdU
KKhnWzkJ/DY12GY7OiXAZx7Z1lxnG36xjJ7qsEKGTKjQm0VTpC2XxYS9MWSa+18RTzqRxDmPA6xC
VmtBwTGwA49h9sH3tUl/ItKhp72LbNP+gBsBLvradZ7ZxXzdnvCC8rqsoTvn1fXwkTJ8RvGS+2/o
4i+2g4uvZnbbwbLiXmMmTWtN1hPEHDJ7MrQvq0scFfhUvCEafNgAVExc64UHJOBlVgvP4itgmTi3
mymsqAiKE/CtLbKQMSfvOzR5cGaQzYnHOcP7nFJSXUrTRrKdbRwaMBnY0VE/o0gCr09xu/RC4RWq
G+Wqcjd8KEAb/w4Ll4p9Ts2E9xNNRY4/D1FlehhaiSzIy5ZN+rCBuOSP5c5P0Bbm3GzYPS7+czme
r3V6uCWf6HTWlxXF/CjqE9fPHLAgk1ejvdvcpAG3qjV4INtxvvHwfr++WcFMeQ4HgKpcWOIuln6b
EPzZtu0znVQ9NSjhwM4v9TZOtn/ic89j+xAVrElZc2tBOlSqDmUHHKFSdVkVheStsReyCdi89uRF
mK+lGlmYlmNcyW8Q6qctsdsLjFcg1KpEQ+cK6MmhrMAcxYnwMwoAusOqm6SEuOGITwS4Od6cnlwm
MeZqy+voB3+1J0RkcAls62bfP4PVryUntfnlw31leVdvQM7a1/8z4fHtVXPVDREjgYj6lPDUS8fa
Ie557dlEpiW9w0w8V6cZd4wCLgMVd+kqdyPOoAQSfPuhgvZfNQrdidxBl6ma5g9KI1bValtPRQc7
w7mYL8k29Zd1N7yfDXyczi4ZbqghDo1d5Ds7Jt+gAnxCVDAgZNS2f5rzx+T6lTA+IzWnQUsZ9YhC
/GG5QcMEqxoBfXe/PSWRryMbowq2Qaa/a6UCibWDsgOs6hBMdRS8C6QEd+eixKbbSfyjkVkuBdNd
xGVzj7EKeepvXpfFlR/vNStxTXIAv0+ybHuesGD4VCVcHONDL80FMEuwijT9pggqsJGUjUpCwuCA
NR3TB7LbV4ZxSj7smC7bcseZfceyDArM3sMMvbhowFH5ZdSiU+pdezg+5dax5wIFnuRlYFWc/Uw4
jH++qzolIeikiTxLN2pK0kCVTas7eCynzNLiAKoyhx8GiFlUAV/KLncL9k06/KNGBza2aJxhX17K
Ctj/gExVrO4Mh3Zal1vbLgRna3ys5tqYg0XR+R8RiF7jH21t58n6qEnaruyFo9yGEfO9zKr+7E+d
ivnRVMMk7TfHLngnXm1bOR1GKRxFdaES0dpYKDIwpYD5noR2LU4YYR1qASsMtvtCq+MXHg5yfmhM
vjga+7bnzxqr/mkGNv9It2qNiUSYIMUOFQa5MJejXjA2QXEzQ91v7V+4ae1UXl4+v/nh6GkQ/F+9
X9DEzwPeD7sE6ua79v3VLHxvhmt0dr48Pix5LJ4ermy/Uihzr9BhCfxCpEE9hfVwjig1eJj+r9j7
wxij+7e4WveY2j0KZWnZY2/2JlNqBVTRJAZx4eDYwLmICn9awesL2iqd++y773C4dX0ge4McpvxF
ToUNTrKkOoOL2jeTrt3I8WA9wvDn/jjhUg2Hm1oREPlziYN1bFvTw41Hf/AGYBXQin3BL8FYi4HM
vpOpVYz179w4LyoPagxK3MMirlfxuIERQns4HgBX9Dx7fy6GYpZnWGJI+ncrY5X73xzaCn7AmcYe
TGuBW5Y/xwRf4kRA0TBRXgx9GkrEmG/e/UVQXT0apBRrMmcy3I0tvcfllDRaUhw5aPUHtOfOHjmN
E21Vv3aUs3D3TrdnXmUh21QGivDnBFMbMlcjW7N13j/tU0eYXuNCbDMG0KYKOSWq3h8etLC2REmE
BorfzTVfJR8vETgXz9TJBzRM54ona7TjvhrE8K8V6BhD0S8F5d0bY9Nrz1HRLafPfhOifUoRNGK2
MElfaQ3YGsHDclUiHvAZ0GY8x90WMZmZdfOpM5LA+1qDtRab8BhWqH4/sr11l2IAwr8sQ8RwAEnQ
9c3nT7KTxULZvo2L8Bug3oqJfaxh9PJr7O1qPTp67+drnPzmpjh3Qr2fG1Y7DiRn1PDbBa+YWFG9
Tmm73HAyH4npCbPKprSRkpraeaRlV/bjXO1zYS3L9mEu3ab+UiyxBMme/xDrzA0ikHTombVQJjCy
2Xiyjlg40rB5Ua/hQnwpb/F9dFpY9ScwtCMc53suMacHsigdjC8X78WR98HaYqv01/JpdI6XP4OX
tjjqg9H05ooVw2BoXLU8RHtwDXc+a7etOjnqZphpT0czTNzYEJMNYLiz8ojsfKw8Mw5ObeDEIUWQ
Wxr8Xlvs9WuGMaJQeUHdXXCnj4nHQ00Zgl+fN4TMuObEf0Xwfhzco2EGRWD1Davusj5FlcaHBXnv
R5C3+JzkjbBEF1lhjqc3R1tLmoimIhofAyNBCOZE+OTELpk4q4BMJ2/mo/KRjeYeXV4RtQAn9WXa
LTJ7Ki05eeKAhPMAVfW1wVg2Erkw9LedAasqinXT15KamEqUxppOMHzTxjTurPrk17kTcOG/d4HP
vHlpjxvIdMYi0xGXM0JI+5tQ9FNz2ly8t5U/dwgBzFyROU55sIMt2koQuxYAphkUxTXB6F1rYjK5
xOm7/l5fCHvmHI4cbFsW4FmKInQNGDtjcGlCMnL0640OeabDGO+okkPex0CoeiKyJXRUWQSe9C25
CsoWl3xkJDISWHIAWLdT1k3zDFot8gGYErmUy0JVyEeIdR0mRajTcQq45mFS63UebXAzbmagnj1v
ttR8htbfM+qyC002Gwmt0VanyTYpULWgDXsy8klOiT+zEMBr9iIpKrQt1UK5c/NyR7XSWytcU2Cg
qBRwtrXL3S6v0ETu5xHJgKZ+XI4oe9Uqrjqxcr+dEb8wZuJDM+HYnIX6epmhUsleoyc6UJD+rdd4
R1kGwloN9yCYkQl8R+NFq5PoQViL9tyC/JaUyXGpwhm+wlNVwdFbpU16Fugis9LVA7Iu2qRiPcO5
biVjJi361E/cC2/nFv5+zAqyJDBo6yEwJ6IdDBmu2BOqPY5TEQnorJsYIK09giLKoTqHAvN+OqWd
p6PC6xbgd9Npt+IYBPvN/8qujCuyQlNqwV/f9iUFZU7AeeNzc1KY/R0vWz8rIDxas6HLV7N5beeU
fvTJb/8RzLcGopeGZRVMI8HicSyKmNIVDTRtYkpd/5rpOc7vVkxEdo1uhN8/hKRHzNrKQpxT961v
aqkDWjLGAwu/X+d7gtMiSqsaqCu/epIU6xxmWj+1KL4En47MlY7UvWtGe8dNxDD0AJo7Q/B8UNWB
J+PjbN9Qx6c4KMPK4MX5wFDEcPP+EAFZ7H5DSEL+gHWGRKwrToLZ1nrZ4UdPwWc4f1Es3UHdbDj7
JZBJoCTjSLRUGMqKgOjO9zE1oy77oCpT8wcFk/fiWX5y0yCQozU5/t6DDmogTxOopEbdYedJcEkD
UfLoh0S//xLcVOEPVGXRoaicVhMzloSrP9nVJ8G0xd18jyQ99QRcIDuNmZJMvWjVyK1+9Kg55/v5
SAOKRAgPFu/nmhbZi9TsUd440QZtpW0e+1ZqCf7qy3ggCpLNX3YsoyTyxYW9fkGlFjcpm6JIX6LO
e1WV/P4zeGclCvyIV95UHj/cz0Hqh7pKdfO/8YdJOUVtuxiSm+KL7hwsuydT56QCRH+SF/Yaz5r9
/lANyOfoRukfyVJj/34wQ/XDSfzNE6GPvQLBijMrZeLpOBtSeOcSiL1kx59qvKUH0GoN6xraZx9g
1ICd2Wxr2pzAvN/vNt8TMj6P2GU1hFkWwswKxCqpgQW7Yf8o/hpK6nHSVj6B8AcsIY64kXcpuz5X
Y0x3gkd+3NLvIYImxJ9QTfGj6mCE1roxHFuih4NP+D00r4rUJ0e32XVi5bDWez/+KnVOLzAaNvh1
Mke57LZzwRqNVwz/nHJ1flqJcgxU1dhipvy7X1nu/o2ZzKKZyN7Lph+aEf7/D/GUgRa5iQePs6XZ
vgX1KqwtWVGBWD/rMwiha3+naGyAKtjmKSvSTG/mP7lo/AAyVBzYf7VCz+2GpORPiVcckZ/gA7PU
4M3i5om+kQDZtrGLxdj7SpyXkxxzvMY/FhJRa0X5tH7p+aw1SKQCt0SV6XOnAClaGyqHWzT3anL1
Hl6AnNGbh4oDvV98ZmZno8Jr6yAvLG8nw5WJEYiv8BOpd93cTQBNmo8cH2huA+rEO5jNfauAS/eu
P6CYTw+Ps5plfmW6Wc6KSX46yDLLURh7J3U/o4p2veQOAOaKgYdwl9AEwzptdkvm44/90Fivb58Z
thhuRB5pDCxLGUCLsmnnGJx+uuYRwrlH8wpJ7PBLOISbYA5DwmhtDsmJ8geObkZlEgtCExdBz6gG
m4OR+Ckk/Fb10jK9oZVVUzeX1pkJpgiyjrsYTI082a5sFlUmC0nd7WZ2cn5lOUuPHbPRmpgBXz/K
9cjZC5EvP9dOTBu0ZC3gRIbwNwkKaktct3aIYPWoPXdKwCZQoc6YkMULARZW0m0JlBewqJDURECb
OFuvxT4PvBS14Kv+c3KVG18Xy3VRrNNA0eQoZP+R2psz1fSJ8MyUvk9fvrPCx9zxt+MWsAhC4pyp
c5MeD0Vfdk6VHEZksD67CFmA3kE/y2gJnUh05e9e2TOssLX8D87VmWnuLh2fiexN3ocn4n9i0rQX
h9z/JUFfPu3+eUj/1D0APtKpD3uDoTmr4c+HlqO06BPg62RMAf7GmmPY9FBn/rZ02wTuQAnEn7AM
mpfRzyojV9q7Nz9RhY9FugM7QUjnhikPIpwqN3gqJDREvG9IIN98IHxly5c9lbAEs7wGaJBTcnE0
U/EeYEMqdfaP78SW8PIYm1tAlkTmeIqpaq4ks/EnXC/6o27c2OUCar4SU0afp7ywv8S3lttsJbC+
J9GBB/0jUXuoJcQJlNWUfFJwyrq8nM+KGGLf4RtQlZsUF6xcQaJBtJoFXnkg5jm/69L9/SvWlvLC
GGgTiO22ZJzyu52CtinSH+e6XpeVSc+D64a39nN2bo/i7nD3Js17QtKni4w5JYz9pk742iUgsy01
KObJ+aHSewK1ePIYN9wIZ/j+h5GSgvwLba1lICh0rtQIU6mZYxBi9JQMIEJMeBWYsYFa8rkdZ4LD
el0Y+TTIPCYVGKxYzJZJv43E+8DzusHRxoWu4dJ9CJCRwBoj1xgJJjZoG4BqL1cYR+sNofmg3evW
dp8+AeZgKoJ5xf6+/5HI1X5l5Qd+xaPF/JYp1cRog5aVziw8rvf7jvFpKsIrRML8hJVFsQrUIu22
fMZ91mYmQ+CtlfY3KafsK7dQ0Pxm+6JasCFpztXUDz1e4v4plXxwU3qaHlwLT8mNEPdC5rJbuPRY
VCkz2lpAwffF0dGMRNviNrftuTWOc75oZXnYipaI4Bf26tTCy5XcYcEMJORKqY13WisFGvoB27GC
f1stiE/iFbQOGGlMTlMn9POrfjw4Iqhp0+JeCd/p2g0yCIYlOD9Ebf9eahdwcBJ4AAReeQBbQc8S
U9+OQF8GYmsn5+EOcSPh3My/vZkCdHCMGqVnjQhlp+J286AG/EEtuNazIZotW6gG8iyWzM4TzFnP
pNJ+yF8fqrcUx2RnsWueJGdFfsfyINcuDAUcOUPTUtn70EAK/rnAbaKObCGe7mt//p+dRP+Tg32w
xrzJja3VkuZncYdKdkbIH5brpoiPW8WjExKbdtU0+KHhvXI90mmhKHteepb9szoi92cddWe9HoEu
su7N5GdGMHkKKa+/Xx/DTeImx6NfBmi2cotJlKzNK2JTGd+O+9r4KTBlYMFZklx+F9mTD+IRghUW
9my/VUGdNPDyQvDbTQjg2eE08lqQRxI/sgDxH0Okrv7dFU+AMDJPklJEQXCGDBVMXUR4Qk+AavaG
BtHwxfUMhB022d55IOI00P4ySj1LiPWXznZk+EuNATizIaiKjENUOZ2aveN+I/EW/sSDfjZA5qno
Ftut0F4DYAB1nfwNFXS9VfmqjEDDfrfQvuzt0Xr1g16aFpF7cBXAzOnJ94L/NoItUsvdxG3KCjUr
kvMLxh0h3tSruYks8AruMFCYSKnNTXTjnDB9eX0eXb0nM8gb/a4rCwsVJp7FJoekxl8McpCkpify
vu1yLf0NPVbOoLSGGU/+z8R8Z1JqvVUe9Gh7QqgWX2USCyycvHoquKmhugfP8oiVdtOfUJ79y0Rt
5TQOKginsZ8hA3hfnATVbXMm2FRMJhd/p0u1A+Dd50AJfjBxuqZNgSMCvfEIQAfUBji98K4tpyxS
ffj/H9V8J9v5GkvT3GKeBU7lMD6KYgdpwwdpqUet3gl9s7KzpGsw/5YM8wXyVrgoWiddG0MxJmIt
V5TjPAduyIOS3M+tvgbWquC8y6Zw8WUtWJoR+vhk6bgCHhtPKbsE8QJVXEK8/cxd9Vl+yo80rI0l
8QIlhnViMMa5Qceo+QTVRO3lVOUMSuSBY8B70Y7JojhEeaYRwD11yaBti3Jf2rSTTm5N974Ze4nc
4Cc8/XLneVLIEn52w7hiLH4yGIcu7xhn37MStxdRLtBBD2t9rcgB9pnAJIV4Gu/+oB0LV2jew0Qa
za/BsyqGL3+vr4s3cZe/h2U2HVNCdzJzy19HY+v9PI+P45rGkqNgqQdzouQDNFd3mBVPWUMn9Vno
dDwcdPmTHFlTHJyBo8oqDxg3cuZMg2yUQJx5MDD35nRHNL2v6hXgLEKCgHeE3JwKOY7fuoAqEN4j
jU1rCd5baaSE7b+sdZ6K5SGp6Z1znZl8z0j/2LuBc+rUtB5yMQnuW0PoNz63zwpq+YhrmgLysQBx
+NIZ4Tgiy/ppc/8oB94b8X3XMSeItOx5LPMPXtbwUnKaUOzXH104KagIzhBkddEoMv1YZDx2eXG7
xyV3PUWaniW56wymKrIg0De7j4EqlzMxoKtCBAPGLdf1t690hDeEbRqpcnEi4jvarluKzusTyXAM
IrhcMGU2vA2Bq3U4p7TWnuzJgJkHUjQ7npeKlxZTLaVCpGA+BGJkNGm+zSABcIepXgvCdFOA3WRY
Pq5RQbbrkRiYmUdPNCI67OSEu4uq47LJLJ35AYOlq110eCAWpL/itAZIeCqTox4EkjStVjibSYi4
NZOYJ9DDZfuG/0DavKWSXoHMtrfNzvwV76UHjDZf5z8Leh5LeFwf0NxcGoYMuoCikYImcKzZvWbO
ksVlbqMB90F1euQB+6WRomiVMwTzFP5E2ieK3yPL8HMaL1fFaHNUC37yZbhgXd0VeLFLpmQlJyBI
Wv33XO4TZd2pEd/ctiGu9QaGFwJQyt5PrGk5hZb6wPloRDeZ1EIkehwMvV5oAYKB4X67DePKMkH5
/T7vOu6YiaWX48M93nSkkFNGWsSNOpotWCbihNzolgDDzPyvvRgP1GiD3/a48AbGpBiFJ8vw3Vxg
cCuwWhjgmIYotdB9Vc0FjslmcE/M8JPTmCsqGw1QyP1KYK6/qFP2WPNIGpTJAWAi4JWeDoGn7CtS
InYtglJAThjXiyZ7BDd4n7bEzuBF9HONDZoayTEd40lxYxvXKAR9eTwZak6eq2qkx7/TH344jixQ
+V2FEMcFMzMiU1WX3HGrSttfclOpvSF6jBvomi1Mdnoa6h9MSatt6vtp2z7IztkhiidGv7QIDTl3
75s3R0L5Peiq6bvzq1Hiv5IICve6HwsWbwZ64kNKX4spe+fjY5TRRHiFmePDNfgNJwjlOEklcr3s
t4HpQIFdIFMT9NProzXs/5XCyeV85WVfmX549Ky1MGTGERDUd5VSFjZL25DDWeBCSdPcGGpZAOwB
SBEcv1XbReJwTSULHL2Guq1vQghuA/gljjnn0hnDLpINY7c+ZFT32+DHgXLJ7sSOWGyrBMellyaz
pD1DABv8fAOfB3NQnltV+EB6WsZOe0MCixertdam8I6PbPZEWwQ4jp8fCOx3pdi0yiICkCQ60CKn
quM5WQD3p8ZJny105cauGQK/+829xUiMSEsKipiau8fmimKXZuwVhE1EJ6JyVE+UcW7rihcyeU0w
cdtCtGTovTYVPH8XTcab5MDlaixWC7m0KMMjqhEpBMufGJZ2p+uc1tOQMtb7bMg4EZ5HPPb5FZUC
9ve3FA/ZhBMDeI4WPcMIBe/X9GytOuVmz7u72KgYEksiCkwhWLmnOnCjcKN2AI3SkRButNHFDdD4
BhfXrY30AE/FqMvVGCpQL736/LJIIpgrBiTRJV45UJbx5AEEQdaQnMYKoLyPXJrzvWGYbbv35a3K
WVx0jpfYITs8cPOd5/w77B+t68QfMcArjSQTZ7mzORJ5reGvZ7xuh9GOBPPyPpuFrxIfT//A6elt
clg0LjLkefdKfd//iWZcWBo9mJqJs8ZdDwChA9VYtHOHbgou6uLzdoIaXlLDMvJfCTMqkPomDZFS
2+WOclfwk//N/eEQ948PiOhgrRzdtCYXIyBM6LmGVL8LqdgENXAoAX9w5jTHRxKX86yfuQUYTy3W
vy/f2UHc8ut61FOPuaNussPW1lBPvtS5+ICq0cIk3qYHGJ0pXQAWW8d1CIxvaWP//9b129jw1cQB
j0+TNnSzM52ap3Muyrr5jz5qsEb1gZ2bRoJcM16EHPdAjBnSwCxoZTepuTDklsz4+4pUkITEkqXb
SSFb5X/dr2BnClmIXtraG4Qf14FZmR3v1uVUQNHIf+G4C4VDfK5dGwzogUGeXHQYClUVKkSMcMSs
m4Zoq+BLJj0aPfs8QITMFVZGhN1QNVnjwpKtekC+W5K6EvaOyKPhgPVpyB9wSFzYFU/PYziY2Jpd
ripaJgsIB//xSljnP/eLEOTuf6ggNiQEAyrzx2uRfy97rMZlonfd/RRyMj1w/Ez9SjDIrBwNPhUY
RLJVrcugM3YsKSYosfHnHdRaKqnVi3ksGbCW2rXZdX2bwewtx2WmG4QmCYQ0016fxV62EXq+GnNX
2OStBxkPq9HY3BSajqhdPSnvQyxcI6mfojjZFIc+WrpQxiRnqTRwBhNLioZa9d/jJx1KP8flXh2x
VLFBw5hK7tojK71Y2H/j68R+YM4/eJM/k60J7pLeZV46b78D2VwUPtuSGpcMUH4bIbAm60yqErjN
8UNXZjxgce5oBUNoLo0erQ+sYGV6ALMx9oHqH7Es0QCoKahJkpsjLwgzw6b8gEWdEmKpTXfe9QWo
e/V6HImD0kd/ZvRrsDW3IqsOixfdYBR+9vpjquEstR/zJRlmAkQpt+XmNoaD1PrgD2zp7MD+A4F5
FgXf4/g5s3xgIadU2O2HDAdFWiSqayOF5H4Tj2i29xy737tv+i375KKpbetrtjdQorlIWGD3AtSy
mxxVqHT/XLxajFBKwZh0kWpJ+p9cg+9EdnJj1tQjqaYqj2qdZWPe02eM/hcUumfi+33gEBYb7bMH
odUoKHN+R4e2nMgTsTU/uTHv5uOy5yeDLU4kMT+3frMbX77PkNqXd043unhTKa5ZAr07UKHpyOrF
eG7DNW9rcUqTpHmopcK5HPGnKNLHtPms1MA1+Idcea4KuNtFpTCDEs+XUxEg/lfE0OtAzSoTXATD
RquJ4ruv0CuTyQPwlVUI1R1pIPZcawHPCIcHebA+cmt2e65J02Ll6y9CFfW70q1QHTFBxHF4Q7OE
M6bXvIya/4dsPRW8Kq3BRl+ja+SzBPV0lR938U/o1NavvKscoCJO284MSsNrcFdOwty+BeV+hNvQ
8P/UIMfaalWUUqfOZJ8gr1TWHiDulNJSsGqEakmjjNlI4aOru7LekLBtJ98uAyHa7tbCV6FKWHTO
qeMnls/sXVQ+0aUJyuTluxfeh45xEFK9mULPNuDTiorA5MHNEO9DZ23X24ntC1G7j4szQcdOTMFM
YpBxs5VgCueaKZYW1MdtV4r7pQiKACtnEJBI/5+dLLoaKYqRDeEVZsq910EdSMdTc2Q3fKKac204
NMJyY6hy9OVkXbNuKZS8BDyTc1t5KuxK7F4Ay66W8QMPkL1b3lg/DwKEFAb528qiM8baoqkcRK8q
N9+Kg1QORhfBVq1OeA4XF741sLHB1mOJipGob9RCFZXUEeDSNi58eMg4qNVkgHfR+ZCL4gBj9z2n
DuLmrlBpnykD/tUUVf9naUDQEV/vxGp31CPFCmObq2ZkKV0vMPhAHhWrCnT8PoAfihlgFMuu7mJO
jKCN6W+Tcmel73HyzA4GSOpWT11wpruchge1BdQsoid8CChsA4hMbE4fs4w4qrzxQMH+BoXjxxU9
ExwqAl7R9DxU0xme/bbgzbr0vudueQVFQYIh1YVR4j5gt2NuQYzwu80h8+YpcqZuM8kGO1NN7frz
E5gpZ6tZ1eewjMnzs5//b8tdCKf/JHV6ZuUKUGVLiqEGxrej3r3QsEyKWl9gPBAEWHj6HIL7Z4XX
fB1n4Cw9SZVV1JvGjiJDKA2CKiZxK84U2yJGDgfgEjUfWcPTbUbtq5851hSsdwpTU5TcvXZOVv5c
SJ2C6ZVT0Fw71OFwBJ4K03QFLfnn51FASpmPFHM5PBtNXDS1UzIJTj578Uptj6GC9PufaPBmNg1k
x82BQHRmGqtgHmW+yLF+pDLxHsj1FgkksHmpXv9IhI7498XmimZBfvy/BdsiceBbt5h34PYsD0mu
iA6+AzihSydWilHRTOco7okrLmip/MvPUoiSZ1PHDAUzHIQVjnclwS2lyBc2kZfBOnwPHfY0SdJh
aZx/9uZAAvT62fTOmKhMT4QeJHYJ1pkc7sG2HWVKZZvPFiBI7gm9nqaQ2n85h+/SRj4dD4Ha3oZk
VBHU+vQhaHHXw/V2Ue7Fvjw3OqDJImy9sjZSu0+qiNeLYKopbnD75zs+vMs6oGvnodkfWmZAj8Qb
Ywlx9fii18XbvG2s5tyIjbhnC9Q2qsxVt76w4tzsHT1KH5sMyH75t6b2hW94ruhzxDFK5sWbWTz7
h861icAmi6/90airwrcJ8OWcLqcZg+e6v5PQHj0uk3b1kKq7pzQFEzCxU/cPl/7YYXaw8kysASIY
HVuucdjY3KzmXpJPwLNatDhEmOdbzgyd0sTTvgWWtBvN8h4KeHE2oxuQ7lCJw74EVgupDj53dTsi
xeAICCOiwdHdNlzE3t49QDzT2uABdlSG0y87FQqndpAJx2SBhSQ6LVkB+CVqMFQ+d7r3pjG0iXGM
DyXaBCZ44GmEdGl9ntD84Ogo1wBmLh+VTRSCzXbDyc/QYt+a4VO7fMKXYy+fHzUUSHDw2j6y/0ug
Icl0Zw+jxFVuDY+qFzLrfo8NDQzK1cGO8QfuLFTtfKtUrgQsdCezFGyO0R/M7ZhM7G1Cmj4TANwm
YSwWaUUeEsJsUp/wd4TM7VhvAi5UF4Fc0I6na2MoUnYPM7tmzqbkHUw4gv2XDz1qso/8cs5fLjcm
ttpCV6ljBwSTgK1efkJGz8s/Tw5PD5FthMX7sWfA0NRelPvXa41dspb+yY4WpyPhZ3wypj7IS8zA
HmcBnVbgxtd/5ZLt6qsMWfNcq7D3nKskNZGXF4WvhPNlN0636rWQw6moK1akAJ2jYPfvUZyaW2uC
XQTbz3TdmxgBArUsXM4+QfF66Gr6t0SpXoKiP/cizbXgAZTHKHFGTXL4/kYXESdmOfVA00sl/7U1
TfWxifvBTZgzra0gDFISZKe6Un+PDIvBY2eQ8aDEI2bUBQICuwDwYYC2Cjy0KNlPnmU+PHDDPorX
F3Yz0GNsp+gAqvCJGzlsbOXjyQkdT26hCxehm7zjvWGoehgsxjVmADSQ+1NHORHTvHnEGwpPcP3x
1dQQ3JMqE7BpwqwTK3MoR/+HCOymOAfCH96l2TrIL7aL3zN9cFkK+joLhjTJWVcZ8nmB6dMhOdAn
RFfCy55XUj3GipwGBjACZSXNHX17eGbs/u/rSTZc3wjnj/+rgIye5DOoVTLv/APh5sty8yDvTwq+
tl1VmUb/VLlvZklprOXrEM1p12RBTeqCb6fsGZ7FKr5LPySC2xmvNAYh5TQ+tmXkbrU+Faj+kFoM
UXnkVQFko+Bx0lFnGtA/tDBJXiP2gADPky7r7CD1x1pbpcDwV+8DU9iwCvd6gs0OSQgklz8ndQYS
WzEnMGeGo6VKOeNQW5v9YJBBArb0x9kawta6mwRFu6+ait4HECDKHsCPmgu4SfUfFpvp5Y4ARjWY
TCahFKy/25TLrDDBt3E74r+OSVj4gBc2YRilEbYkm0DklYeGBPVs7/IegJYEBN8JLHlNxRyTary3
/yPPlbekzC3RQaW6ia4TQG3SJeiJFk0EWh9RJup9gPB5aOe+Wq8sS7nu/CtifBUpKY5IPAOiZsCe
jWehdpF4kf6uN/+X0EOC1sHl1ehiHecWbWLfr8tYdk5af7p4m/vN8r/kQJZZmOuROg8Ox6IFf2FH
3hMk6SeTuS0hafjRkWA1Hpygve1HlYlw/8XwMszGgXBkZE9BcuQId+FYaLRy6ZmKe1tamOBWRosc
gjTVj2cPJf9BSqOOGnVnByKvGXyPatgubQOyJrE1M2E3wszu/MLtEo9qGkmpJ+ua0qh8DLZPfxDI
iLK8kxnKy0tUnpg6Ba3H4+7zU6kifYWjx1LEMTUP2wrLhaKM0K7lyn+4Yvvsu3lhYeq3j4xFK1Ld
B1ALdz6iqd4BdH0rOm8u9LOKovTp6+j30Dh6YTmYsEYOSA5uGE7f414AGK+hoTOoPAaUntxmXXMg
cfy5Avu97knkNAMDbSGO4x9gpxBXQKcOASWqC9xsyGilMZwV5uvxt3u5nBsHfvaFxOW3vIa9Br9H
XaBnrQk4AlYxyh4tmk1GIAi+K1QtJhf4UPG5beIPgYCgQZuKXM4AqRHAdAnidRvpW6u4SVEm/ago
jG2MMbhjuOjwwrrdHtRWhfZmuGfxPRJePvo6pbRt0xRL43WhRbV9C6Od7/iYrZWXSE0xUQs2ebKO
U0dZQJ7hjAd3Vq5Jen7zh1AqjQ+kUsAcFgHgrAzdGD7wRDaNTRy2+2dEX/no84680dZVgTJAbA9N
hGGwM7WmzgDxNE5XlyAd9S7LJnYRHvlwsbVrf8RimpqCIuzRAhx5xRKCH+iENhrhdRhSYZ9nI1rI
KFo61g8mzjTndouYrnCTnPI31rWqXwKD8LIr89JUNuGNCgza2eNgKE5/nBE9pQoGEs+rCGkvLZw+
G8jB1Q8pDAGNBNNY0dViTHoCkoJeOaZ2diQ8G166BgbrrFvdsx3BL6Ip6GYLwM5c/m531dB4Qt9i
UY7J6xgEV8iQjmqEP+ebSp8jXiozZCF6Zklga1RMR4O72STxK360UQQyuFJ6Q8sCOcsE6GosmBQh
0zREbxWSP3YWOipaJXtEmChttKPX3J/3Hd2MgYbI/FDWyEk68dAVxJF5Ldqhif6kUgh5aaanwrIN
9NJAAzm4iSrUx//ufD00BiyawJOVLauOPCH68ZTwp3O8b/Fl/HAhN0d5Hz3RpAbuGLBNRJKVmm1i
l/F8gdU+NOUB+YPK8rWwMa6kXua20pAw8kFKHvKtxMk3Uajon5sFiIOeLunubuP8dOwcjjlqJUHB
a4toy7MTjJjimaq7+VkZUx31VOf/LDB3PqDkg1rgLeoI+a/Pd+D6hCT93IIg+EY47MyWVFbH3m3j
gYYgNRuz6rrN5HfMFeFG5bixVkK1n5+o94VpnxZYozNPLRV4+ZcqI4NjuBioG3eSZ3JF2lyJFLnR
80xEr/OEPJx54vTyFluadS5vHNO8yVU24AdIKWkdDOks2Jn/tlZow1Wiv3DHMBIIcJeEjrrOXXYN
kehfE6ZK65OxjOh49qZYBSZe59yxD+xmDzDL6kVFYRMTghOMYqngHbiYldwgl+ezXheUgbcJs620
8lZonyJf73UY8PJIylETZ5kn+/XxmhiALSqBtwau+vg73EW7us6YMGGtArv0RdyKl3Vn4Kc2M5yg
M4gqx1tDcQbkM2+eAMkcuH497e2m7zico/rQ3IsG5iPHQ4V083af9IH6jxJtCyBxzZ/magCR3GIx
bgTf2/EZNW9PRhrbZQVpe4aJghgk0pSBSNLmMgZNPWsYvJFEVTIAXHmhDF96KPnZU04wwMGwoIaL
2xfGJkiel3ckewz6c2R91iy2aaOhTT20EyzXdTpGAIKaulpBlNkdgK5w/v8z96QOEQOGk2Mby53z
rBmXrchFRpbdcw19h5cZolqBTMnx1bwDPou1Yh/3NPW4fafV9DbmneaPIB9E6r0XzJ1VbvogwoIE
oyEyXmSj22s9Q0PjBKrP/v1+kES80gtB8F7JVZOC7/SylkDqV5e0EQ7uLMC1e5vmATrPyZ24a6OE
G9JGoC8b5k97tXtFIC9j5y3wJDjKRhfaoG2jv6YO9cd/dHrr5nMniDzZNcrPAe0nn4kcpLi1Z4I9
mCVCSxkIuJs+o2Iu2IDncpyAca7nslqKZAtEH/MSdIMrwKORulBWvBQOry9RGb1WrXb02XWzqOHi
UByOKWxuTO9gAMk7cWuMhDg+2By5v3ndu5aE0JeBjvQiYwuL7frOUzxy0Mvsy1+XBVUjq39IAUsg
Ggb9dSZwtU+Gb04hLcj4RWu2JqyOhar3/XIzBXAhtdw4irXklpawDskiOCWUpfrsnlVdJ6SrJIYa
80VV8rBmD3/fHw8YpeZy1CKtpmI3vBPT/DALLIoe/IqaWZgELJa7N4PnVTFU9dzlf3sXQ5qtgOhA
wPWy7hq3ulZCGqK6E4vK+3XsW9eqbckREWwIRPaQjqt/GUwpoJAIv+tQjBC47ShlSeI5zG2+wWep
HqF/b7N7liwrYTacTPdk3jGCEP02w6eYySjitqWbHJiV+1L947l/U1emWaQYMt9i8t4dWw6C/HZo
C5o3OxokpHVnX0aEnu8NYFSRqUIQrrsBdQMc6fvF/W7F1SSNlXjf/3iD12hL7QLHTPuOQPnp+Zei
fyURCEGmikO04FJNYc2kF8PVQ6qu/VcCKTp+YxpvVdveY0WQRloX1qZqcPTInw/dduhzPRb7wDV+
K9wYWK5GO7W5tm/xD9fuLYw2YweLzBwowlYX1m9XKQYgSZhZg5gh6MdNII3WqV1MNFT+jTK5p58T
3oIScoebgzH0VAva2A7GOgLjw6ZaUzIktATZJIffX4AsMjIlYuMIY9z2wbc2EDmn6hXTAzJ/JY3Z
j7i0nuo7o7pNEbePoDuJGGmkWauU+WqhfL+wSnAPzZpcikKDCfLWfVr37bi6YxourYB68v+VqMfz
H+/CRW/3kF+uRbeZReoTsieJ8NPqwjsB5r92eb5RFT3s2sKc3Z3KJZdHNjGx1PJnLjIrpGs7EuoO
pZEiT4wmaQKloQpyFle9SpSotMIVug0WFz/d0VQHtcfu1MO/hgZ+mOl7KS4QDGPiJJOrgyB+ftNq
i3ncQUG6CwOgEiWgyGLVCpG5niHFofcFDiu+Ne0nE1i7y8k6rnYJeUnHxlA/8fJwLJ6vGAgJ1T3b
OrsEv1rJ4o04t3p+rFBb4inJNfEuGulfZZ32g3rtBurOPvcVWNrk24EiEbV7EXYfR/eSDNxkfHeH
RNA7cWWDFAmkehCFdo6OWgIlfephoUK9UabtII8xHJBHpThkV4ccjwB81nNsZKkm/uy/xiAS5dJK
EeWHn8+vRuHFr51YiErlEV6iDqDmwEUmI5mTC6QraD1k3ZZt6evEeLaPEoSYCIoS5IiAMeL3dpEN
KmxkzN6tOXKYYI336i87hmyW0h5/POUyFTHuCCZZImDxmnkmGlKaLHelUA5Ju8vpS36TDJviTH34
nWQVtQRYI+t1I3W375m8vP7ASwAmqXhqwqlA6IO4cKt/R+BshTFHkWySMRYJ/kdU8Vyxb0cxemg5
XCEVgzVAcZR9xcPkGjDffl5mygMhO70pg0UpvJgcCuAlRujE/kJExDgYRWIyBwcOrvWtwT3ctORC
f0HwxqmHzW0DNv+1IV07/MldnfyPffUALmHlFF1htLLoeYpBT+FPdiBiz6a1Gok03SXFcp62xsk7
AsGqPS6Pk+Y6BtQmQKb59vqRa2ehMsHhoL6gy34jLTUxndd6omL9EHgzaL6qFoz1W3CjUybGwZC7
1czPdzePQhPgCU1a4JYAEY2OywchCXw2DldPloPHd3LAekNMkMCBXVP9pmETIIQIFyeglSAQBkMw
BZDffMWmtg58D5LbC0woSFYwf25GqTQvHyGs4zM3i1Zfwjl1XYzn+MKbR3kbCwPbU4rQgm75UWpI
5vCG5UN0hv1MsuUowKSHeYDjYnJ/kCMHCrJkKzjV/P7j/kh4Y7cLzFhkh1+1jtzJHJG3bB7mSnXx
ZuPdNKaeqKRgnApfkzMA6vMZ1nre6r/QyGfdCMFXDDO/ZXBBd8xQD5BrcESzkxQQORQquqF4+6VW
1yyEH95nffFc86nOMjRJ1RTuBoaN9ppA28NuQRXoBGVshtZ69kTE/lpGmS+7HS7U116cSDfjRHkH
ocX6cLJ++I9Tk4vsPXpf9PIkiUWEFA5G3hd9h4bhscgQyaCe9Vi3gyViga15SiD56MIDohZ9pHhg
5sqmnQgUbiu5N/bwacyVT7qpeDxLLcxpXyLSUGGVlSj+II+xOfiE8ppugLr/vGQQ1CLyX4ApT+VQ
fkz0P36bYOBYJ8jba6J7Laog9dbCJtjqb0Qilbu0D6SrCX6YUPP5CCja4wWCk24t3nfDQMB4NOMt
WelU1mWYV3WQlP+moyYzidaUluVm5ZyFtopWu7OYOHwmu8HzLCd+nWnGyWKXF5cNrPvLD+k13MBD
RV+E79NsyHHlwWcGImHsbyI9Y+XX/4Uw7t5TEDKmlOARVSI0GP34Vy8NNTx1ouTHUO5FDFfQ28cj
3FZ86sKrtKZJuxofc5ooE34RkeWTIulDGW5clVTD4JL0CcotVmEL76Zs20/BijcbFDRhk0WyjksZ
hruSKn2ZW8vIBwsyDJQCvtEHmGFM4tWbAmRVHu4vBewrFxoAj64KyeRfmsUjbKSlPiX6OjjgdH85
iRS8/uLUsoszgS2KsTWVVIWcIe+3u/k3fVBRSPWpCHhBS+xg5hxRzAMm9HMUgXdlCyXCYdRO7o8E
PgZROe+L75GOaVVdRwNJfAMw7XZZ81xN2/MTakhnYoRCVgj02bkgYUA9xjDCrhNIVEyA3znF/XPT
8d6KR0Z/nkTZQk3UcRsaSxOgGkQBjXZRhqcwl1JrVIctUVOQNi20iKZebhEZCbA4aOqBI2bhnbCb
nq5LpR5iux7jZY9UwHj2kj87cemX5XypqgnC/9iJIK+BTCsavEzCreVMV+CBq96cniX0dmZl3SIz
73lCr8j1l6NIGjd4m7ngJ39GF9g6WvrHRlyrWrs6FPvsl4oT/9fIkWVLkHee8ngZFTTOhsgE9Qam
+6KOZUoUU74ieuHTWmJgUEZwFkmkbavYjnSovEayooB4mXMtDaPBaSwCN43Aqf2WeTqPFwJznPvv
laziRfXcIF+Dsu6Ta2Lt2FaTPBODXXyHzbGoAFT/gvvTZZyrqX+MGokyaaOb98vA9Dg7HhOwwDnn
1SmsNu6lxJvCdJCOPbfyiwkQXHntGF25VFoYr/Jd2cUbxuz6EJhrkut+crE1KzCn8PDkLkYjH1w+
5xFzSvg592W1xFgRbzpSSr1FkSIuokMcENYDI/RWv7BN6H2L2aSEPHDzG6oOnhzv8sMFHt6KUJ43
DG+mYTAw/oDCM89Am1a96LAKCDyPdwA3pu96jbjOzrHtdnC+CC5KyohwaA48p1kM80MVlvqfldmk
/Qcx3abZPGtncrNFPhdWbO9+Lhdeq4UkFG9n06h485A2Ekvz4ao4jtDRBk1u0sIgoFjfvRcgh5mE
d2JCBV7Tls9XXkISc2ilHt2sdIlwDftDy6tZ7yPqFVYWK2FalQc9Sh25+1loo3Uga1l3/RvSBY2B
BN3KHZpJ0OyifZMcvAqKAJM7z0NUwkBX4C+AgepBxMHF+sxECndWtaJ0yeX6BuQIGphLce5oGGlk
jne0hHlnlkYIOS7lF4LrcV1eA6x76iWEeHyt0kEL/Hs6in/hwbipzhZfESNHDJ7N9JZduZAUQBw2
4ciNxdTEOZ8HZXeZWgtwza6kCXI8aIDN1PRmnpkrW1Sy2B5fldC6PnNoYD5rNWe4ZZ0jht1Vj8dT
9kyEcMGAM6W7GoFGreaOMkrp+0q4wpWsiwsZp+pykTCz6RFKLD9iv13dAI4sBRgUdBSp/PBdWA4b
V0w+yKj8Mr3ghWhvIY3US6RxnqTXqsBh4oWz+BrV1XSx/FKm1iVv35jp3tZObgxdn14E1OddaRod
HfzBNOwGWKRSe6pp4ZBw+wbSj4/R1E2q/zqJDE4vtq1g6R2lUXZoAiDe724lHpMfvKMIMLqseWQ/
OiwU5+3v5FuQPnMhdALY/w9zO43zobpziLkPwOQOikG/EcLb++JxLk+VRQdhv2bw3p1xM6JLTxW3
OZc9kImq+TU744NhgWBGffmuGhfN2hp+Hn3hEfmlo1uJvxSb6BUdaia/hdoewEUCtPVUghGub+rJ
Di56ua9tw3yrJrc/aqtVP76rHasxB0E7Vv4L1s5kXsrcUEOz6xBrtx1a8cJj35vm8Xd5j3q1FHvj
wJk/x/0pWGL0nw5fCXTyKU9TA6tEHOnbA1EMqVjal600mVjhdE4R/k8swx3NBE9kDcxbH5nz7K4F
EtHLwhUQhREUCKlosl4TrkiVMKy6nzi+Kv5bMsWUXSgEQm1R4t/bMlsBRUf/lfu8C8u7OcVUcF56
XKKrdc2MdOzEXn8ZXHqt1vnG3zBENNy8EFAHs26BEJEyqSMgQDSX+KO3SpFvEo3sJR/yWppyd6PQ
Fu2b8HiDXf5NDn3k/CjIOc2SiMmJ45F0+qfcJtBCpQEcozd5+XkqajzH0fplbtXtAYmfIUi1uf9u
Y2Sk2FlwkS54Cdsyd8EUAVIdBn8Tk59mzDZkeB4esSLCmYvrP8QMIx7Z/dYteWg8CDcre9XrSBHD
abcPwTH68OaXaecHoyWjOqpOJ33z300IG8jnISntaN5E1+fWsLxumcdJdKcSRtTGg6PCCpRfftO3
eHoOOlzX3FydbZItW7X6f1GzWBWuK2+gS21sChPea74NkQpk5+xJT7mENknYKxEt5DwgBOgR47SR
3sBjvNaF/dktEUWll2pqZT9BTr+QFy/2qiPn581416Tsnx3HVhyOTfQGV1sDeIBRKdD43czGSIIT
Rs5mVJt4Fz5s5ohmQMwlLm2tPFXoNYzZ8AqWNcawX/HNNqmP3yQI+fEcmNI5o/WZDwAi8/PLMCAe
I56n/JHTD2vG79yd2o6VSmhZEicU3HGK8D3ilBlQQzfDlmokWs20qYWp4WEAZ3OBWdejyp4s0qm8
9ewksFpYwwy4A3VC8J3F9UtHth3jKrsXBJeQqbuS69YugNlfoGwXPtxcqnWUKjn6C/9zOfNa+U92
IVyOsKvqlXXfQSsUi76bO3jnZtL/hBh2pLv51V7IFjJObyMHXadUydrqx5e51vqSolCjyMdWMDVq
Ziwfp10WW+hAloGzl4Fw0XXgDpPczzZUb5kZ+lTvtYJFT5tTm688XTrNPaDNuo07vovNJVJur8sQ
DXz2m4nO/BsHgVOTHVAbuPFUHIfenAhkWvXHn/hNOeQAS8t75h59p0ADsNGfTp+b5+wFtlJVOz6b
R4LKMBRxApB4H+ye0QMgBQGZkAte0nvTYXh/b+YAjQ2dl0opIQ+zhdnw8X3J1jDKZ0P878MwPf37
/XsEp77C5rZlQVEhTeGS7gRN17CeSMTd9jms9Ci9vC0+76M37DZN3kaRenDKXAZFmYJTnGCFELug
fhdEyywQ9Gpa/6aRPoNwBXdnEBFL9Gq4cD70lZjYc1GN2p4nIQfFWmyjT7qAr3SOB5z/m+oPRt5G
p+lfEDxQeUugDEXw3JRklZmvsoYCvT3r5+hD4T+GxofEPfMr4X5w64eJMosNHpN5CwJqfwVwpAZ0
Q7j5Cz9bNrHUOE8Q++8bfVWKjS4kC9r6u3hGMgKo9ZExdDEpiVUifyVn74j1o7w/FMQZV2CxP02W
YUhQ5jRaknyyM2hZAa+ZyvLqYWSj9lIk6ScGLEdyhEG3IL0F8roBTkdNidgQzwn4P3U2ayYx56WO
RdL1Eg3h3Gin0jiOral5W2Q76fl1d34Gl1188FxqStcrSmnO/7G99MKJH4r1l1r9x7hbS/7rIGoy
tD9lV50EgpBG7kAzlTY8grbID5togdxgA5ou3W6UvJmdUBXo2HZTDUzfdrv/sK88j+JHEl+p30Dw
S4CAQE8fXx0fuGfzPTt/SEhLuKych67pWw4XV7gyhOHq8jqQzdeInycEXQqCJvywNCOdBooyFagh
DcKdod0679pfX36mcAlkTmXVKpkjLLlJ8Kyc5qC4Re+NsmwrtpXcvdTabRBmrcmYe3mlbGGElTUG
ll0FGqh2GYyBJaofOVm1gSa4E1L4aSfaGJTlENz042OXb5oW4iYIiY0mzH/ir4XbZelWoey9EgM8
AB2JFtk8mgX7d5Wl+k4Bc8t+0o+x4LbQyJCRWI3hhIBvsuqHF0YNxXLiyKC71jP6d8spkufQb0PS
IItXnO0EMaoSQZydOFMVn92GQ5fPeuazJrmXU3OARf3T/K0XuLyZKhKlMvI2vWszIFGHKkUr/bue
rKPF6VFcj84pn3Fk1AwIy0kDF1uaAgl5eAOe5UCfej26cyci5QiMq5n3yPNJiodzbJs9QTb6LrWR
oMdw+rKbYxxrX6Sries2/r3qPNNlo+0Jo68tc4ZPaYMUA6I2jNJyUDhjvOSODDXVrt0Fpm9H6zLQ
O4DF3WDr/KlJ3tKz/UAHE5avMaauKw82icg/4iL7ZgxGBUC35Rbz+ZYKByOr6ubG83jBkRUe9Int
5Z2NtL62f1I0juQWYjP1yyVSDvv2cB/QkbrtAKfCRpVSuVmYmCmpYGExW5YbB4e/PzqWADRtCJUb
07N0JBH4ojoQG+6GQsBppir/02SzUfwLE3AzZfDXPwPDVx5v62xB1+pWw7937AQlWaA8tDmbyiNb
Ys3rvqGGd3/e0iUmzs/mdjZKSjLOJsT+TNuaMCr5SEg0pmdYU7ccyUVgpoJFWp/dHLec6dQSl8jV
W1BrphUirBiC34WaKJqenO1s3n1C4zO4HJeYn9iCiQFrfbdnaw49e1X4ZkjFsBbbvJQ6YoZ3mW57
8so1+U7AW9VDhGB22ifuVlEsG8rf0BDF05mY4IPo6Opopvg1wpS7aE5fqfWAknd/CvLTMmHb1faF
qIyFSyqoiR9XpRBNpyiQ/Ek+yCCcfqL+RL3xEB25cB6XDuptHyv9DoZ2u8Ap2vpnTtbUikpDcfHf
9sUjSxlRHBJ53iTA58mFp4bZdtX0D7h9onMuIST+Qeg16H8AGNllYWHP5PdrkOwLRIOjV1PgRnoE
w9KBknigMjrXnFwjePgOyU2lB1rcOAUyMjpbZ+z+FXJV2DKuWPLGWZjxqPXMn4lbJAia7BKjy5xE
5B1SWMU516FcV5eVx2tVvN5PlvM+DYRn7LHSpOlMerSqLE27aeETH7l+TgRBHmeBxWN2MjjMeihK
cUDV9Qy7/CupbDVcqvWa6qvWm87WD3nT7P5NgnqR8xfyPOvtnOhS4pPO50s95VBwz59hqOIMWNJX
1fiMXjmCccWF61VCVKMaysDupLVdo77ebpnCA8Trs7X2mIzWcrSxRfsvM8I4LtXb6Z7yECON0WQz
sLSpfjjjaBuwe/PYm2xUM3lwmiV1SpGNMwuKFPl/lZbAtNl03RTdzeketRYuQ/ptHFsLtvjLFYq8
DYPD+lNSiiikopJz8TX77t50a5pAHDUOD4wylBkzpgofbuiFg1ZYaEFpMSaHWvQuoTdSYc9WxPmj
CTJ0KzASurhi3OLo8s7PC/xDvVJVbRoH+DKcubqug8n/QRpxtIl7KngykJkKgzEWDpgSd5Qy6CKk
hdtIVXcr64OGW1JMjBowXeVPvEfDcfX6hLuFQ91lGnnbtyN3EzcH3UlM2+TFi5+7BCG927JsvY7J
6a/A9/l5VOFjcxQFwQTtruExglO2QyE5xh6XVe9BiZAhXKPT50gqmNbJh4jZEQUf+aHtLSYson9M
m+i6Gv278ROFI4nkZDul74cnVDeqgw3bqqS7qsnd8AIs0T/omgglEyK7+l03eH3b/VF22Gbg9q3Q
4NaCs021Yv0tJn2Mbsd55O3b7GeCBAZyQX85j5R5wboEqBtngvcLE/UPUBnhc56almXUr5qTnNDs
Ts1Dli/6RLJu+jCB4SAakIPS/NiSSQ+76tm0dZyDk1pxOibXU0ChRnntsCsDweM8k5HqgkfYX3xE
6au9knsbbDRRMs8coqHTFe5nLHMFP6ZUatm4ey9HMyI/eIDJmlOITqFJMvXC9KpSy/OBlKkm9nkA
JvKdbstaOXC/OUvIQCvZgEoHhu2KTuR65qFKMQWVw/LdpUX14eCzgjFfoohq+JlBA/1prB1WRXJN
88dOWxdvP4fxnd5cVZ9B7DopCi63oyhqkEdMaJgySTFzbkSC09cIjb1eXIMdXv1YgAB3RhXox+ul
ffezI5TkYhKBVoI/5WIOXXykOlevZNR/CuZVclE/UgL6csAOzN6WPebkENAbzjomhVncFv1q/3iV
2DpJNPC2PLrMwR6I0F7BD5aIQXmLJZyxG+eSKWD8MpmydLHS5ZLTdSScvvQz+k4EdMXIaTCudAH4
4Mx04TTKeUd10QKNVUpnchkrv/lmAMu1sh8HceSerUcjEgKXlLS4n+1SSxD+NnZKjjqttkKH4Zht
udwnuR6XmQuX96e9yUu7nhtcugCeXdUz1I2jTLrEKkDmZ/6xAlJDLvIVUTRicHICqJ164BQmhzYl
2GMd+7IOlA9Moq79ca0OvUxyo49ZncOlt+2JZ8HHHrQ+eF8BuyNXw4cUBNWF7Bo+J2sswCg5B6QH
YL2vh97TGL2Cc6OSRQnkeTtel9TRQXXydX5znpJ5IY8I4jYpiCBSXpBKr3MNo82FKm8fC0IBF3ds
V53lIndUA5Wys47vovxirtWubtw3HhdyTvghd1k12QgCzxZSLsoPpA67XQSXZ7Re9HequzfV8Es3
4dVaeV8UNb7NG1eTvcFia8BEQj5oeID+N6dD/9MGQwaqHZxKxyIn949641b6l0qktHi8lWHtTXP3
3q+vjo9Anuy9hEv931LUbSt4kPgHyL7AUBezXIvTidwOPxULms8yFSRMVdS85i7hltBqRdGzVfEP
nzsYA+uvzIuD9bETdB2xAJ7ov+BF8ajp0PsIhPVlVS8lhd5LBrIt6zeeEL5Vbrye5MVmPcGW7bcd
bjvWkAXLGka3GBEd+KCJ3aXygalJqkPSPW9OXKdMbfb5issKM3E+oZodiWDVCL0VItmBv46jh62c
qO9/UMuG8QXO4gU3gsrgOO2LGZQG/0b8C+Dg4tuNVpOHahsqWCYsGonV7z5V4iPW6+3ZbZtTGCFI
ZeOj0R4zGQcnUZGlNc7Mw4WaTdS/W5KS+3nHm7491O0EwHdZqyVgxiGHTstg3acRvrJDHjePyhfV
Ij6XizrNHS3OnjRFObSXBhg00V6iln4arP+2wEWMugt0WMg+asspgXAY1r0PMDZWvXmqaFDd5CuC
zyn800K0xOOQqEF65N2aChH+WyKIgmd7nGFs1n93I+a58AtaxDWdnH5teG1w20V+K9j21OQHBEH5
8NBj8Dj/AXrBVQAnY+gTiw50oV1YSkRL/RIuTh2R53Hyu8ZFoAZA5FGEJZ8w6Coi54Hxl8sNoreR
RQHynW/9dUTkVZna4eH1EIdE7fFcOwsUYXug3VSWYOSVS7g/MbXnUqTXLnERozyfi/BI9YqlT6yg
MopYsV2S7Bbf9OSucTloduXWShZsHBKY9w4QidTn2RnZuwCdiYjxwuBJJU2DW3vPShFwew7KxL5U
8U3wMlCFU7VZszxp1VZ8qK+qdMrCLrLbtESj4KkdCL0u8y/7cmvRzLUzMtFqH4MYC+cJrjw+n5dG
Ccu8PsTlOPc0Nh2yE8QA54Wl2Aal3eayzyy3oM0UUjrpUNYFWheYpcd60qm4gAJJU72aw/iBBjGR
19shQHXO0T6dKjn7RO8bJCSd4x9NikvGHRqXEv9dlJpQlIpadFhP8EFgDMBUB0aMJW3PChcNpNnZ
YFFXfX79TGqt/145sBJP59zBnyrn+nV2YF+PntP3PazBWzznGg/nr1AltwqT1c3+FjskMPs0AAER
aAHU8mz5S06oDTp3AG51A1C4krDIf7zEoFQraYvwlrq+SISk8uRV2zl7T5KoXXHm2H8jkmjTaSWG
r4x/kmGPDCIyBU2oYMZ/a9zqXIBlivLVr14tqImwKVCHJ4BjexPs5oxq+6EifEHXuytNzRad/mX+
WpFJohc6/scXWBrOxeakTDCDNzTg/BsLTVpeaJsjkYCoQz3qkX9vUceSrFw4ZFau8YyIuup/L1TZ
VojYN8betfTu+nGNLCOxiGXapvrbdjWzk8xY4xqkvHsVHZzAzJE+fpdOIB5TwTbhHyKVvjBaDuGY
evBoy8QnaEUZuyEO0a/vz1Pe+3C2cLas4DwtWdqjW2zzze0suBt0nMTclub/r+Wz4uImZdBZttu0
fbruh6BGuGVMYMQbOksQAOSRpjZsA79l4gRAa0PjCLFefLz4zngSItHROBIGIYdGBlMVBVtNDFhw
WDf+EKBeu0yPKcnOimeMX9LIkdtaXDM3Eufjx4oENN0pThVblKvXm8TOe3Fu4magI+Fg+uI5gGpZ
PoRPbbrLxJZgaDdIYsVpcOx7giT3CtE3c2xoHf0I5dPpnyeKgV4LURLwcXrws/OjqNsP+9O8UvuT
BUo9/9WTWLILXSuJ2uWvttisWHt82scViBsF+S7k2K/c/jomU2HxQOTfQno5HIl659Bujl/CGKhZ
dKar8PLEtBxuNq5vlf1B0RI1ttjOiQC/+jvyACA1wIgCTWKNwxC79PVGZLA8xQdo0YUsX+NNlheN
oSA92cKl4fV6P14yKjHmxZk1J4KAYZWDEoD7YZc91FpNxq+WOKIcBDDkyDUIP3uK0j2sILzI6DqW
KY+2Ao+/lzPh5YtMvxNp4p+J4G4Cuk3zMHonka8fStNYLbqY0lNMn37VqyoBjjeh/e8u7E9LAyCk
JKTSJFK5oTG95rLcI/+C4NHBVQu+BD1zemEBmquzzFaN8IZWov++RmRqUgulGsA+JqUGwhRfOcF4
SHt3+FjUytcnd3OxnqvCW2gqP2Du7+/6me8o6iwHSMqkPsm17wEmZEW1g969HLf8zW98GQOJM2Ph
cSeho0PgBDNY8OFoh3Ktv1H1zc4M5/7m2pwK0vwcTCDp35TPuyPvnedGyFBBmpp9jrWCFIvhi/Ao
7G7LUfU1x+IV3mtVu89MEojKBtst3oYmjHxzUwVWpPWZOw++xO/mfIJaRobFyNt01KH7LXa/HA1v
ohG6rDrrk6+RU8kCbNh3SnGMv0bJCIMKw8+vE2mTSPX91H79oAacsWPhPXfAafQi9OwqWSpyXrVn
WdgRYLsv71ahrxVd6NMWTl27lYNFGQB/38o+7KH5i0TEXxbBslqu2nx5rEOdYyauNiSfXfPONZTj
HZEXFBNK7MaczAJbN+02Ejz+uqqzEKcNctvkbOgt2sUTJMSDdX9r5QfKy2jFOW3v14kbSIQUFzrA
d0Mkm7snQohbbwiFdBgbI5PUERXtpbqReyt2geZpI5xnhVOFJnqzX0+EiimZ6XpMQthiLFLfO/Jg
3N4avtvvS1jp38kNGBh4Gu531VO8CVgPR18B/in4FP8tNZWNTi0TangrWXJ/UQ2q1CqaDiPgcgxX
gbZMm5sqh94vmKPhKFK/2AdhigDL+ta+4V53bJfEvYog1kqU1x+dJscTaunEX+KkL0mhqqXOBIhw
FYuodKoXZwGSwiCVi2L/tsyPqzTezuiNoiP1aEoFPmkOo4FT9tMhHK0JbZ1OIvMQNiuewibc5rbz
fnOprgXP1oYmwE7iEhb5waQzYLvlRxvGvuUPVnVjmYQ0bhJ0QMRgOlwJhn/7t6cEg55Q6el+LeFC
mBZokmsttku3b40x2dX+BoawzbchDTSgkZzB1XaFbDGhUexSJavlNSWgD6nH4+KGSa1gVZHw3bEJ
hUrNG6DDH8oh1eH/R0bFQQWaahYPmloYrY4Rj1JpaYRAK1sNRlJWk0Bk9egedNUO5HLSSYhQsu4r
p/A8US+cZI2kZQJMzespxl7AfmrqB7HhLbLdpMKc+ZPPdZ7oO6naXxpVx6hOp/pnxVFyOFRfbC7S
8SOGzZtFdSUf+Y2rDESebNchxob2k0yB1Ax+LWSJRDgLgGps8HDK26P7J0qkdrtlpVmP7t+2eGCG
Z45npInnS0E3CvCJ0lXnjB51RHAVtHTgXTbQ9RCbivt0Bs/V3fqMoDKhM7IskLhHI9ac1mISIrpx
tGIH2YgMd+h2q6kiITec7d6YtQAUXQiQxUGoiIhcS9LOxzT2SdNlqoe+aDK/E1w6YDyNEZ6P8LXk
CobcI2fFmLv+dOPG7Af9mTHlpIP+REMAdJXDT4Mf3N8vQomWVkkk6vM/fwsYXdcr9QMgMGYMj/T7
O5ZgDjjyupa4ywpgSo9qNafHihE3UF6V+t5GGywxfjvlIzyLQo2yg6P0pm6lZNt3G4KEh02jCiv3
RxOIiaCrYldJqj+/gULgiFImfZIVY5eGAucGtk8XxoFizojw3T+9QsY1XwER5bHTT5qi7o2bRnJx
abXZoCon5qvTNBn0SSTzhTb++lzdy9bt/I+M4xW/zRh2NYjq/Y6oqEY2BUsCqyJXtAv4B9P7T+Ip
7A2xPjqz2RaDMJxpYBzLKUIcwTmCR+mCxy0MQIRvbAst1yhDsKdJTyHHTuIco+z+0wUrbV6YaXIG
ycPrbcrXrcjuZT6Iczzqejq+N8p+9Z8UAf1BPvMgx8RDN0a9wIK76QgI6JE6RtsQx1UFP7qeehRw
mihwu8uOQRxWRy2IiGllreVOU3nBshTyoodJYvXXhgtnUdr8UwqV3N2ijRjB2ofvLUdEYSpNRx6d
fZyS/nJ/KOozXTdorkUA25v32OIICg4kcTOx/BwBVK0kKrkloCQa0KvVka3cuIfKwolumjQjO3/0
ECrb8Ap4hindO/anNLq193wIOElAHqs2CIvMGnAFIvOHnYHZrTKPwR+BLq2UQrVOPJoz8GJhBPce
KdWZXs0KMwAx3rbv3rKIE1l4xC8l1ErLQzyAcvk5LqI6a9Ak91b+jw5YaElnFQqUHSHvl7lqDJ3b
y2ViQl0bscpwFycTRfh0K6Qry6kfNDKVOL7BQAPgo556IJ4bplqkO3OzQld9CjP6Qr5/3duAQOCO
hUHythiCY4L8c1sDiF3dCCcCof72mVZORtRFDQWKyTLdwLklb0mfFVN+Z+FSOhZn6PugVYcZKeKc
3sDmF0o6jXeY+OxNo1XeVqjpcHtyC6QLhrZV1FxOeGUuq77pGqVfdXdPfXbrVpO4IGR7h1rrr1ut
oKYh0w8RadVM9jNaw/y60K/J+0qNlP+aNTK4PuSJMJRcfc6tWeBdDfMsByxQG9PfKK366iRQQDkg
l3LdIwVg8MOReNFgEZFtONl4i+VTNI3obPj5UPxmtdWGG9v4FqyEWhyMLAwos211PNOB2Vk/Je7O
1/2tv4CVZ7CIDCFtrfu5OBKZcXNeC1t4mQnN33kreTG58ycQfZGcZOBvaEU69lBafRdgzSxT3NTb
fotJBqxJIHMirj5IGAeGrRG1nBaoxDe3TSUN+epXpYbCZy01Fo5YRvnhdMCHYccfDNhyNP7vXMHa
gROHAUCPj7joiLMPDMjqUzgznthWbWAF3cQBIwMvkXe2yFl1pH91sC5geUG3GxgoIv/300LvoI0K
nyw1CLiClJ7U3W7UD029RntGAgMnLZ7+FjGJ5OqproiwYc/saofj5c1SIPpKBPBwSVyHd0VqyOij
SRfGNx8CKpqzE/QkO51OKyqppXFjjcK9uOZUuviYN1DrcMcq3l8eB8JJRLH6/hbDMxC6+lQ2GP74
5CLjGisaf6FHJ/qcENd52uenTh4US/qayUT/bdfvH5fagoHkeXNeAK7nbGgbYg5f+lo7r7dywAOJ
SA/IajdiDNnW/l/HHis+s9PaAWRJ0gokGBT6AnOcbEa8XmGv71Y1xYYS+qNtHigkdRqCQbKvGE3k
+X7OvPjm7N7oqGQl0+hcFii0re4b9bJYWj2ygC7XMZw8lvy2UwZ+erDYj8m9qOS0k53o9C+FFSKk
YL+JRmjJI/1b+FEw9XYbdPZmNYstQM36HQcPlgE2jAcsgr6q2BjFAp5EfikhsY31gwYj7OVOt1/c
0p0PpOKcAoede+Og45p0YnIRAi+XgWjeN1/uvTfwGUCu2WBCHgInyEVXzp/zm1O6t9oRhqulAo4p
187R6MwNNcOtvlOeZmsABLl/oWqw4s4eg5UG2z7JIt/IrqHU0vi2jK9sstncUvwMPgyi7I+56PEb
yjkfEUCvVHDiNmC03oh2aOBVSHTBZSDam1DMZEs08MjwmUXoXjhvRCasyJyXRHdxk1J5wP0vONNE
zb4C60NTKZg4x24JBKj2y/kD9TstZY6Dg2O7EsIBg/6i4Fm5sJeOIo0XTDYawLEfIlIOTifnaH5i
6Jyx4TOxZaTTOWng18EmWmfZpPhG0wYmjfxyH40j3dTYyMkfbVwFL7vQvU+YgYCmWvOR6VglwSe6
9GpP740DQBnyABQQZEjcKxfph4L1Jz4do8+ia0nJsSmYFB6R0tufA1sjZTJBDKpN/7YRwSm/ShzE
isuP3bYfjX3c5y8L+z8Vns23j9uz6NeOleQml+IRGHyodjzZkmPkoh8QeHoDx2cMqShODZCvwRAa
X0tKiZwYcT1FdQoZUu35KyHx1kh9lMfhPnp2sAQ4YGOJiqMRbFccZ4tDzSJ0mgCYAiBqGkt1kgcn
9TRmnP3+O+5bVtCnu9htzO4s/YtvQ8GV7me20X84bf/kFQcZRRcL9vROOC1un9Hh4RvJOJsXPFZY
T3oQkwcazSTo3OFzLjjuyqQ8YOyMWy/Q/u8vWC0wNottjJCX2SYh5MLEvVbBFSDj6O67UGI/PKrn
v5pyVh5NP680dI02df+8+SraLFc3eYj4wWcTkff4r1AVhVap34+ZNaAy+7XirmSruSjgX9fy42wT
VeIIWFLHfyTvU9i3+yR6WMhw9fJdbz9mU7iOwFLgesMs8iYimnAvqJVjV9wh60LoBwGdO86PV1S+
06pBK5DEwKRGar15Bv0QeVJ1k39vgN0OpfZR/88hT7ZieQikwcookV5TjXhdpUtSiLqARNtUeQqE
QoEs1bQdtmzCn3d2qgDwK6Y5vTzgWwPlUP9C6jDFyyLFdlLaIX8tLvwLglxwrdHFXwd15iNua4sY
26s/QIXdOxJtEzLJQbiOLOCjZJtI9Hq8C43t71f5/p5qhxsS+XCLHFGf/M/RKwRp9jL3pgAJm+y6
I5bZCT462sOReolfdFo89i40jWzyJ218JJcaAk74EjwFP1zZAga13w17k2Q9pE7cvxHBER0tSXxO
7DngiRBbqvM0XEr9BOjlNmaCXxW71b9BXA2UBijtsZNzirzZnQpwR8N+dyfQwsUzSbkrh/4eyPi9
vfyJWHypjxQSF5hd2sGcjFw1CB/qkD+oQP6//UX4v6i4nnOifqymYlkKxSt8yzHQIEtd3l0yObfW
ib1MqvH2p4TlYSOTDv3uwI3vlHdsX2h7sW5vcN1Zw22pp9PTc7C6Kf0BedrIkdpSUCFG+1N1BdgC
rFV6XNYukFWmD9LsPh2fKcvmK8Sry77IFIzkkVMcdI4TLgP+NZB+5RUcsz47FrFIP28LMB2LSAfs
JprB8rmiwg9LPxnfWMgxYlpQEKqAHkhIT9YWz8uqYftW0QyfVrvLs+ewstyW7cfSGaunFtLuxP5f
oWjrmw/YtbcQ2lKbV3apR/2Vs70zZVE4HYlSpBEqa4aLLwnvIo6HaBNWHh+XTENR77I2ZhmsvU1F
ap4HTOZSbo8YczC61rRF+h8GykyJIO/Dpy3KLYT6/dGuyE1r2QxfhH4nae2zdlzfiCmTH8tEA6Bb
hP2FZ+GJFQ2DTVohZtijlyWwZW8v5AwvSXM3x7AEYsMCcAxc/JZLRyqBcmh6w310P2qxQA9g3C3c
Ju2XarArPoAv74YIUNjr2H44BUVPGZws0xKFbnkulzxI2LpFexxRsuuCwX/F0Q7DVSYmBNR7zIZP
jCAxj4UqkLiYEDzcrGD+9fmbkhmo/vpv0QyVeGIbUs9VVauZ4TmHmTqP8r/2DHy+up66O1LCsgPZ
95V4pwaXOuJvj3RQZkyg6cIVJAjDlcb0Lf8cPdN0BqOu6bGtghQP7jadP3Pbey/2kwuTGdGnPWd6
Sq9vC2aKUMoI62HY8QV5yIET4OLUGLTa75K2ztS1brEJqq1maABT6LTZwKd2pf0Mv7aMFV+F2XV5
AodjmdweO6BpdEMUlbL69bf70YX2pExTjONDhubp94pdaCxekEvj/SNsbli4JyL+Xu9CU24hW68D
pYu5xtH+EEYRXMvCoKcgkOmBWJiS5OlZl8hNi7iHUyYwgSIQujFu/srEUesxrzEmikjiSREqFcyi
BwV2gyG9gmwkOu8FXidSXauBnDTIc5kvlJxb5h8UPASjGPfGrAhgxawV6i7AIYTp6co3dHXEJn9S
RYSh+Z/nXw/wkQJOimv8sCXEmOgWZwgxcejputQMi5W5pF5c1rP1MjBgMJUNMUTog6+UzXaogons
hNkg25HJ0i3B5YWieOoznYnH6Q6zSGFyfaSqv+dLa9F7N21kOYGkeaixYv+0Bp+H1pXytgdq9wXc
+YorPq0h5XMC6ZkSp0IwgpvkfQKNSNGVThByVIHhuF1U/Y3YdW8rDCtAsYQA6slTGj8ah2StOw2d
X3+SgEF4n28ocwUc5ENEvwUjDtx028FMkGNCRGQsLg9ume1VrZjLYg3ZFDgDiU7rQf/KhZ///Jf9
G/7SeZxt01pw3VsS/2L4sRfXrILJQGnY2VGZeT7WTx5zVl8DxB5R9+3ZJ9TP/x7Yte6p53MfDWn8
C/z7Mmyue3VGTaswv/um1QkRpLYieSZM7ObG2YkmqVuYqBTrED2/rDXmd71TKGi9aBkCGhSPyozH
5iDRd65O+RwS4HZDnJa3Z0+fGX7OKVoOmJxdDqmWr4TmuRE39qJkhBtWS2FUus/phVWO9dWikAdw
VqVok2BCK9OpyowLO6zamyS7ZbQ3LgscSv+pBMrxgXiot5XxhbjaxLSD06p++Uqr8FhREJ+eKIF+
jN+3ScRiJlfmfD9ONI9smkNhGOogiuN5BSlW0nDPp6z2Vbb0FolhXkqQlwjUrONWk9KKwb7rKY2y
cwnnH5uQs1++RHyi/wdSH9B776YAuN87NIWBzUXIx0+c+lvlpjIf+pcStSUEHx5tGHm+RolwhLYz
HGUn8H8Pj2veMtlPdF61c27PeoVvx6O9jfiML3TW1hj8qdVM5yirLbjj6fge8MwSoCKDmmxM7AIh
lM9i9TETlykU6t5iVE4la6+ARVss5ItGUoMT0sHmDllBEpEijm1WGq1xChfB2buAEUsTS1VD6TLE
3sgRgI6z+U+E199Ta3cyEdm4UtamHgzPXApAbJEbodqlH7kJf4L+O1mwKXOUOdS6e2QLkBRIdzM7
6gzmz143Pk25NqxlN3kK1kI4adrG1yARn8nxRry2B5i3AQ+1GrkcElapibbCWrAzWkjTGlhvgV0W
FoYrLJUgn8OcX3PkaX2JSKvP/9dOwMEJsyNStHUjaNycB0Q44wq2BE5/+4S/d9eRaKeua3Niq4h7
eNLoOmvIAx1e3CvAgXU2Eg/ylgYLOS/2XljM3CRRTve83DIlUkzrVid+1wouvlF9NV7jx7delVse
uMNMFg5J+QQGWsOsDC2MtvljV+MmY2HmvGr2kjfw/4CO6OjF2BuWm6GMKG2nkjFSo8N7jO7U1D0p
oOBZXeZExVqRCUZZWWQllSwA17+9C12mNj2D2XEVNlWqvywRtxvsKIbS4NUFlf1K0798sdgV7Zje
kyXUJblLQEOvFb6N7bu1cdqpE8wsfhTtHFLFxXylVlL3Wrr0tshuhPrkJTgWw4uZdNohAR2oxYUa
1rNvB167KNow8v2MNS6Do2Yo6W0Km4eNG8W5hmSLd3NUUSVG1t2pzsxJvgZRYmJMzpjR0nwfWf+L
AqlGs7eoL1V/5l2B1sgYxgdIV0njPmSfkkL3ry+Vp9IG5H7xdl0s9XqWwY3EZ9ODvugPxTF/QYPB
c5J7JoSi/uE9Cu86+q7bImV8+wEoGYtSHbeyb1WPQyRSd+7tJxmxqchxmBQG6dSxRXkl/qjNJHyH
jfEcnzv7iR3/syZiHy/YO1RI6nXNMok3MHKvjb9UsirhIZIC3xW6XWuR/t2/rMoWH6Sz+BdIRk0E
dFLQBD1jluFOpwCQWbSKFfpzkJcJgui//XJ5/5Y/1kSH00m4APCBH9qfPQDvEhiWYG+YY1MBLph3
b/cC/ruoXu51k2rjEEynTQWUtDPOMRCk8x0akfLFS0pCLj2dxzfl4SBjRtEsI9i7E4F+1Ab+6d80
RKxkYLKxzJQl58RQpgnzQ0K8lP+hs1EHHR7rqYhQfUkiEQCSdu3DK2+9L8Po+6hOXhoQxzDS5/kL
EpP6xTYfGSFTR1Dj0QypzWTLRL+Cqo+ULG061Sur/pSz+ocha5wDCAKbTUXaI/ykT7/qWbxi/c9O
+rr6UVioTDZ3GBM/rx/C6NLf7OrTODPQuQE5pjy848x0nuPkphqZeB+i0wS2iv/rw+OfDy2a8Tmr
6xPWjXd/dCio+ZZeR6m4EVRyPoNkKLWYOJjJwQ0VWJrfFul2CEjAZh3RjnSfIsXcB2Ddpwm9OIOg
CzRwaEaymw96fBWMkrrAiXa1cJ4zmG+bFDkT3xPTGV0e44Ms9P/OJyLotiRKgwjWBtbbprTNWgv1
Tt70P+1G2RwspXq8PUR5cMXoZPdHnv+kEOWMgr6QbEIGFEkuh8vsIQJHRiDnPz8uUng9jF6T1j50
APxS/o1dCUClMj/OzfspDt+V5fUZCcuaDPBun4QJYkbguSGF2/izANHlpP9jEMxFdqwGeIJg6yhs
b81ut0NtsPhV/Xyp/0vj0UDIgaXf0xJE1uRxEjJEwM0lYF82i5/Q0RCzz42M+grq0zUuuK+Nz1Rm
Iy/hIKJTxPsVxORYYq6WmCaQRv+mvUkd3OYstH+MWrzAPjEtIFVSyVfIUZpouIUVLzTrGhdqNMGP
lrIm5h/BUP5Yuv/OdL6otZl7tob2tqHBNMfC3n087Ytu9gwQRyecFk9ZVFhmZ8D1KuYs4PltEXUm
7/r+aGVJGhK6p6njUCW6T2DfY1b/SK15YZC5WQ8nkOlTT4qJsMDnWdy1syYgTxFgezRYKb8a9s53
wTSUwuBcxIqWGPkZCKiX/QGr2I5rS02krrxOruDWvHQ7D0PPLdkbOvj8f0RVL0294xqy1BTpW2FY
A3CUqOTLTnC8ons/wmjpB2u4KMEPuLLltYxrUzOlzuLt+mDjxhstUlwJGoIZijivYivXqljOBxCc
T0CVnNcYNQLdWYvv4HUDAKI6z0Xn3OjkmwR1q7iC/oIvnJijf+QGVq6pWW16IgEtglmes11jzaUa
AUOY+yGAQ4xcqsa46fT4uxDS7NqDFxIVFKO4Po94/AAqNe+ByJcaA2RgScLYAsfkcSFUqtDtD48x
B2HrqSPy66duOLtmNSGporc76MCXcW/5+UqDt9Iu6wWhHXM+9GTiWvJa1R8r3MtpuK1UQjh/YN55
JRVVSegdJR0sJm+s7lWU/zGKuUAPUyYshU4PImpg7QBgeYGdbNXGOo40nAbsFdRCPQqCrY1cZeRt
kBjw/FguuTmjz24zDA/9ipWOOezjf0py12LRVenfV1QxMe/fgn9NxszvyVrzV1UF44moSYAacmMy
vfEqYmA3GCt8Q8e8moPP9SfuEg7aQ43OR7tJlS8FtKceFiAHIb/3EBaIRUNHOzQ+Y4OnhmTLvOaQ
nwIYig3rj1qmYzCDvJcQ1Gtq+nUV5L6y6HqXCGYiUaIa2AMfXYPW5sTmazjTNaAhFsEhbOs3nEZr
wGuh8JrwLR4HxTQL8fdzrldg5yX552/+YGdQGjKtPAn8pgEJSzw0/TTHkYmOo4CUa1SigKjhYbHW
xF+JGmUgvt23tns1CYohU65R7IU1hHatc1Wqzp3Nxm8vMoW6L2wjxXC81yKvsTE01jQC3eqj5u6b
UoGw3YRhfoWIEkaKNjdigzkwGZzIVNJEiLUWFfQwhTF3Ir5HxgHwwWYpSQmUP61iTm57pgH+CIMs
89LW6IjJ5TRRRRZg417zdQIOvOP/RwpoZs2q06Z6NexW20j5q9ENUEUCZ+1jvbnx2B4KYiVKbMin
lslUu9mAYPiZ/Xgxe7iXiXZOTlhGlOqQLvOm5APhGASpkcokQC1S0qsbuSVTqoDT1IUq02qplaj4
hX8eVYefib9ZQPIHi+xGO1IpFeyKwDn9tkLDdbpIEtUgpBMHkDRWTd7AGq69XjcN1IMOJazBDYT6
LWBDE/xCzWSbnePj++T28wX/swY/SH0V6OshcqAFDgSnDUriFlKSdcF5zvGYjMsaoEPK/ss+tclb
hTDW29MeNs8sICCH5cgqTv+24vsv6z1OcZZdz3paQzF/VPI/yHnRRhqsE9Pkc0WsOnCfmU9Lw5FE
prTsznrzdZTxuPk8aku59WENUs3KW/vNhaJJb+rYBGBjSX9SIOGEX1LAcKWdKua4Vt1J9PvsZxSf
yTvv8wgba9L3tAxJpGeZiAvVVxwt+j+A7dK6EqGXAF3K4bgTk55Hu+Jh4TKLudiJjAw8jKivpi2F
rjXamGoMMouALBB4ByIvTqrUpFi4wIcH62m75aB7KPcrhxXRwmLwlYvrtfFdJ2cQMSl/2e/9dur+
P3H+7yyiHmN3R6DDA4T9xlTKMQmzqXz1aOum/iaVaBhw9YKQlFDTYyjUliyYwII5SAMq5I0uw5WJ
0A8p3ScfJbQO2Mf6GgCWfpYVBJPeFZM9aN6LWFksy34xYXHFZm+xQ4acPi5a1xFTyBtKv03JURmh
Cf6SmOJiYaLv0+sxWTv+5KzHIl0tx3EDtmO2CpoIiJwAmdhT/YgEtQQd8AABY9mm/nl6qpM23nK7
x9r8Sbe/4JgBNjmQhfS3lrIIo/v6p4TEfzrCjKGoL854pL4lJ6U4BeYmRFkzshtgoL15ycB3v9YY
mX6m3wVKw5tigqTZgQ+8vMaAeTqhfmzFFFPVNwfeG562MqtVqMEE9z9WcwRU7yWRWJU19UGGTHmD
vqoGm9SgJFpcpy2LVHigHxOAfQQNbhxhSIJd0YkOBJ4FfsLQGN/zLbWeuOquRv+d/mcVjk/CXHcu
TLa2388wVGWR51Ni6b33IZkgGAfVkao8+PTP1f1LkqppJ/2SM8r/Z+Vb/bdgxCVxAYxPSV6KPzPQ
jWrRfScnZZ9wqDA0x1BT7l8yV9Lw2j8Z+o/UmZzWXnyVm4FaBgIqAzJ6OiPvZO5VYs2R8H33SRfi
NR4JanZsQvR4ItFGNLwqBM5s6h/dkLc3dDXuQON1jVZgnLg8/bZKch44vi5J6F+GrlTDxK+sdapc
dNFZgYx6MlqQVe+PxCkYIXCkC538XVuw6Ip1x+fTS/IPDm+KN5wk2XLyalfJ411+YjlPnClA2/ep
VcKdWJJlwRUnjyJsdmw4GZb5GClZNvMmqUUngR8au2OAIHhJbUh8JFA1Crxjv4uwQ5CcX0p1h5Xs
EtkiZJcBJUglxCukKkgQt8/1z1mTet1aSaekv8y9kDK6RjwEa1TP2osobhplEeJKtBqqIOVmaREN
Kvo5iPkTIMMsc1fqz80LrCoYiChm5skg/jO4XNEthlvlgxE0nN7As/dh6pV4m93lTqUTSfRE1yko
1SnPDveZjAi4TTl5PJ9TFuhFsFZ7eJFt1O1XAKNha4at1Z0U1uWcJG3eFsHJSBZUfye4FXpJAvsM
s0XZLw59iqSX0GFwhSyq/u9FoMTmk5o3anomzffcshqIESzbH7Xl/OAzXR7JbBkhJKhM7vWBE3IB
VYMQuSugBtRU/reloKpKrf0Ec9xB5vzot3TKDWRVnjiG+xH92/3ApSWmYUVF/37BdtAi6WqWukoR
ReIpZwq1SKDHcRYFxPGhXhsKznRJKaE0BWhwCxwFhTG79jklVxHIXZigiEiPecjZeCYr2/30xld9
CZSYsCM99nGOsu1XmmuTfpqBIqig0QrD4EiryHcQ2R0PP5T34NuvgiqDBpQyeF10cXSqrkMvUvB3
aJgNUL3CJEDwCEhY5jlrLa2b3G8y7CqRVRkulFyphqr3NUwA1VkESdEmQ8X5iGYMK3TNaqkRyvE7
/C5yvf8xutsihgoO1mTT9OVExRMTWJiK6SniYzCqqUrM7pYoQEi/r2NXTNWuQin2eBh7uHIw6cTA
OviwNl1Z71f+7/hjeOzk7nPE7mB4Ya4AMuksi23Ur0nrejnBsKw4rjphkK1mHKe2CbLGTH8XxBK8
a6Ug7rSWTufrbrHy37dDOEHNMazZe1SJJXwQcJyulS3k5uNdOcbxHQ7PFbuF5P2SG/dqFHrEq60h
BTSM4XkFf9uE9XQ1q5AxPqaZd5FtFj+4t2xImJKYGTbnD7N0EAIGldU8lFxRYNwOlNuzPAmouZhZ
TV3/Ss4ECm/SKECIQTezFfteQ2j0QLiyYQHQZYHgzDsoo079Anhgyaqkt3TSYyOK+0X51RjFgBa0
UOQJyz1GFbkzyDtoMAQV5tD9iN09aFK2gSql3/Fsr+1aHikPdY58ybmY3MeckcO3SwQsQvvDtqsm
ddH2hgRX0sbSRWZlhfFcGI/O671B0ZWy60dpn+7Q9TB2r3uLZmOMQOBbYLAnsdsvSbQvD1ZrILUt
3Np0p6FIeGRGcrpHbgcVnoQgxITKC/FCs116LVM0L4tTGswMsTPOVEk7nCOlwqHlk0B2Wctdkwmq
fB8aXd7GX0RGReKj965ZSWn9j780ljzncDN7L05uIwU1WTFPLUY850JzMGxvOPwXOT2sjXU8a2AR
2hCXQkS5QKa2MCXFBnTyrkSyBBlUQRlbBJ9owt7TFs8xrimiBdrc7RpvVW1kfkAaIbZ53UPomX7d
/Kn2378SpSUSgdhH+hjg7NAxhCWDLfFDwXOSIT86OSATRnwHyyIzjInn+tqZBqAy2Jx+ZzanXuyV
Aub+F3tNnlEsx/251KnebMI/b+uuWMPF2teTd/Zw3etqRy3m7ztgN/MwnnYat5Scal4OCwCnlpAY
UaAWB/jsatdM2hajzeKBilbvXcnw+qCTIqdb3BgOJgYI+YgCae9/uFdePJn53SlYPYzj0B8ydlGl
vqk935yKKNTM9JvL8FOq2eOaj14cbj9QpFtmcA38P0DUoVp7qt2lbs1jggEf/tiT9+Jujjvwb49h
j+8WDiTuIRAlewkep/SfWm0R2SoOlFPnzUS2dufLgyCv6gXuNa5TAahyTxTpdcS2hVqz1v8Oi3wO
FoVOUd0DpS7E2+PA4BOfQpZ4upfNoypgiPJVGhGoOVQKte/E/JdfeS8VWw33Q3/oiLZeyQfJ6Xoi
1X1icfCRrbl2ozW/RkNmopemDGzv1VUVdiYHkmSOd3HFHtFUreR2RLfp7bX4jQW0qWl15smJO79a
hNF+J+vdSK1XSw+YzIBGBbb46dzCFC37MIHreRaHtYc1EbHzdp0E2D/a3oiDtVw6wSPmfKjI4VWt
D1e3wx346S5r5cOtw6P8hWFiena7vRtd5LWzBHGYAehOsKSgIz8Kq4O7rEDyFqYx3IEgMUg3DBhl
c2AuluJv1CmxF1mirorKT7IbwHCPcAlisDhlpiP9Ra/x2YVEi3ROmAeC2pVsX3januQNa+DZBriv
ICuvNvzrV7ryyo4wDUARcg3UJMp5XoR7jhJJF2jfGO16TxRQfL4mj7cl6POWU5Vfhn0bH03sj4fG
euyIXWU47Fiy7e1pd3TUzw/c4UgOBSC0LAwrf75fzmixp9u35W032eNpTrtrQzAMvwlrkKZTaFvR
jVWfBnmtq/RhFP2Yjbo0UmBmaaDKhLDFmoKkpf36IliDSaEjCFXND87Cm51bkT4e0by+qfERgsmh
GQp7K8dkFeXAsS5wg1OUJ3b11CrWbiQJqBeb77C560otzTGhd7VG5Ok79z8nkEyqq8VR1NlsmF+K
6umIqOWCEtalm8QFGzFu9xZ1RVEP/5s7LrTfPzzB4rrqLzN7DTp1eOOoUKFsffQngTM5cC379Uip
po0yGTFU2SpJcnvwIJ44BBIRjBTjPR0N0zhRsM+7RPqip9lSyFusRuoW5yRbjeSbO8rlrpiADRHt
59qcIV2cpR1pUIkBoKwUAybG+10WeNbYBmCxR/U3UasxBtQMX8/im4SPOdYCfPq3sXcxD0/m72p3
SdQ4B4wBhGVPG9qaq8gtFbj3qDFsso5GEO9/6eEUHDcG/EcWYNeWoBzZbDPP2gA6Q9HHbSMvcSVV
AcLYy8tCqCp6eL+PJv9b/1x9kLVmnwrnsKGuoWWYvL4UVhYBQ65jUqgsN3Q8174G/fxm8amtJ1Co
SOJAt/uNvxOYWV1AD2X/kwNY4cIwk4J6RDt07zqNdl8qoPuLeRhCq+G+UP+jiKtWrbIHu6kLfp5z
qJaiyvrheByP5o/R0eWXVP8WbcnHOGwHHNmCRomh6lbGwHYvE7ble+qw9KoaIVNXvx5NlVfjbK9/
dcaSe8FrPRueM6yeh3cHrWEMoxVLGfiVd8yPM8Vy8MdrRMJgUfJrRHX9YwYkrxaeigCv1PU6X3zA
pWe3Z5ylLLhe05BljH+olmXpZnW6CVQeRVqI6eyj1GfymNNkUnwQr42CGA3Kuym+ZR/Pn4/ln8OO
APxw2PObWrl/k9aJy+gI07iAdfmBRVoH6wUsUbriksYDgeUZbUpGj+vcPWF/EUtkMmPfgI4iGiSp
+0GZY7VjkvalIAw5rNRmn/DJr25dKThBxmtC2Z5V6c1yL0T0+iNpNFCs94fOs8omeZpip99r0zFM
LXRx6IkAd4N89yHcvGFDlgnejZRGGmmzqdaYXW/6rugNpCac7R5azHfnxdE56d0k6cKxGw7xZPGo
uuRJWrH7YAl2BBbMWpc5MpUJJ4a5peL1c90pAIGeYqMelczUXAc8lizZ6XnaWzx3Yma2AmZwu9hT
iCSWRgx+7symTmRwqUI63f30spwcohIKSfuefTQPwZE9PhKGSCr8Qj76AKBw7JmU3XT6QXHASwtc
vS5SAi03o0wMGCMF9p6keZ4pmlv0c7QmoD6LlbgNSquG+KA1Z2zXutgXwu//u6HNWyC3O9BXwgqK
jtIs7L8eWb3UUx+J8LNxvU5mmb9+/mNB5EIfMdgyE9Ut2XxirpyWdNM3yQ4ZGVsSZpxGFg0NU8nx
o6jZ0wFwLYtJrCBOPtS1nYs3bxF1XCTY7C/TiQQhknAUN1c7DaAaj+21qAFPgKsLJvdZLHj2ODLj
TQQxhmnxsA2wuS/h9jtomIXAk1l4g+3he2MknB+OngNC9NvnzaMNEfguPeLRWna4OBaN74bpPo13
w26s+3cX3rFTCrvbsgmblq1hth+MVYdnX6zeqUuWbND4QdlWO1kA1Rgb3ti/AkMhErf68p+Zx9FO
1uOjJ85UAJqq/2nbut6WN9vwO8G8oQUFIDqUwIuDywJDPZA+2HfPWA6UL7TMHyjpAKG9EshsYm3J
dMVN3C60Fwlh64j1/lybTq15U4q/b7FOq57nrxYIXAOJmeDmoFPaqHXinL30q/DdtLvvxmNQIsOO
xDQFkURaDtEpAKbW6TeMzQGZNhGwLeTiq3xEk+kbZMQJXYqYe6mUwa79mfKocUCdD4eSbRk7pHY6
ah6fGHW33pWkIYz0i8gD+wjSI1k68U/1dTj2MYpJQqL/2jvosKIs7Qwnb+ye13nTphOi5mrru/IW
gIWLMW3AeV/vlxLKL+iIwz3FV7xU3i97GB+qH7GSLjImLd5+j11NJ4Vqru7RdAoMqc5lHgf9BIoL
TAUX6g3eJjVSa4vuBdje3pwUxL/hc3rYHgBwetGEBHKGwXGO4KRBIFCly8Y1PdwA1xHmF3TTnmAS
UtS3NAS4JhYBzLjka+gFgDmQaKjMamU0UPOAQ2EUC7aUA9MuqbDpA5SURxHupykvI0Qrge5s3CGP
A4rwJZMOVI20LKtxDOeIEAp8SKptRP9o9UCUgd3C61o49U7h3KMWG4Xt6/ritO5LnLSPLAns+QM4
lu/oLOaucWqsXLDR2WxcgQimlGyrRm0NpmP/r0a2ffrLnsIB83ogOY2tX4dI0XXu8jbxJMfcaX9/
eRzokY+AqO7+Ic1jQ6nU2ESBedmogECcBxKb7H8I3kWlaRr2XqH9oNVEwm9odjGXmyMwHS3HRWfO
zX83Ovkxq7BDvhe5kS8As7L479c4cokfAEs6O4KAYm9YQbSsJxWwgwHfGtZlbur6K1BzmCbIkqq6
EqWzeya0vnMYqw2hjMw+EU5ARHTa7QyQNLY/utOfPVHJC0nmq2zj7Zl2OkwAghCK2dJVeVXNXbly
fGAOA+HKIu63NdSbQdNx2aDHRmNIuAWl1IWghtTWMtZfeAZOVHvOPMY0pXcqSaQSxegBtEgWpSXQ
azPyBQpeAQlAmwblbDtcWsq+WrP8SwCcs+Q6I3F5+lIU4eZ1V0GHmaFgwBZ9XbJZ85Q7+gfR+urC
0PTLSeQJ7JWfvbPfqD+hTxANunRLdPsJIwPE5qI80V0vZ5+UFKis/RKyKo7jDIiO7EXwH5eid/LH
pXsY1y/SWYE/wjb+3/qxpmmJucAO3RQb+f1fLANat93Bq9t5w6V0ODNRTl9ceI0rfEOo+3qeAO2c
YbQdqIolzdkUrSp9j0vGQR1yPXAH3nKXX8RuPx4RySONKuM5aidgLEpvXoPV6LXUcvGSuvcwfYAW
eAqHoadeEXvnTtJrjZFrwUDBxOlGl4BfxdvJXwDv6ximwl61L6rdkLo6L9xbdIlNIiNfgJnACK/M
xheC9Ej20wFplu+Q5tvLkrI+XmCjKaOt/64IroZtgkWNX/MYrdYzYwIYE6xDkZ16lJyiVQJdt7g9
iwk4Wv9gKLZAZRxDoJxuFzif04B4kTwsWv6GhI216Kq76DYT/MB/5a8U3I0LFrdQvU4i/MvFXvtw
zkhOWLxdMB9EF5KpYMtaDB5k71SNZELzRIghrJrzaj7Bk7rvie0gG99eA8fS5ZKNoQs5ZEBhonYL
8ROmm7gndk0UYGgkpBwkeUMOPZg1Srd7BJ3xg2ksaD3KMnJboI+oQLQ3AmcvZAfGnI84neWbWP7N
UPOxbGzuZY3hc5gD5P2XZdHRfTOdz4BxsSX2OW/HyKWzZ/smZzdFWrOTU2DMd4BCgydRm2k1PLeT
/ekvysOaD/oXqNl2rGlHrlTOiCN4N1USsuMIMzVynwtXecMisl+3LzgQcVfGzKbBhtDnwVv/n3al
BhIgX3n0Bxk9XiOj5uprCDfaf0tuQ/pI0ZIGni2ZD0cniTyMbnMjJVSFfJmLxCdgsFo82YxPNWWe
0ursViY5MGFLwLHhBvnub5IZ/y4HlQlOVOO/yAJn5FNagCr6aIiJGEo7TdhSj8tCW9KxBX5+KWmO
3pyA+y5dr41GkLzgfNvUQi1ZEGkDIm2d21Wa7Rn0HV9mJ2Pde5XMzs3/TViyJ4vDDCmDFgLEo2dC
JFLuAV8y9da0qhD7CmU36ZlLGHw8IPqVD6mBvvp53bkoB2oSYQrM0eSxFHeTVtxfZ4RYdy4VPtna
KthX75xR3g+FoVzMvRBqQh/OsiZYQRKuc+Zy7u/SnZbWt6QzRLrt8buMmB71oklX8UpO0XfI7DrY
3yHJhEqrwMFdaHtk8skz84z5r4MAHLPS2B5Ek1hFHyCA0QDpdF/OetkjIYOFZdrGhQpMKMtVRP6E
YG7zjYQIZNgptCpfT9QV9RhFbkyCyLYNQHYqyy0FwFBLdLoMmGvjhjQOIEViZWZIc7jRLe1XL09X
Wog7JKZAGJ94qfDL6Xyg3YFU/Hyz3EtEmLL25rVDt5XrIR1kysZrOWt+RdXuXlgjbD3Ql4vivN0r
+bxHyvI14bH/h3YwmtaAAiWBe0W3PpozOfnmA1FcvpO2eLHZ5I0Ql4Xqp1cacDs4+nI4ly1plLci
fbxDNBUcf2tLNiLkgH5OElpFvLKZjKtDh48ER2UbyxQoB1DT0FJCUsK8JI0mPN2lEyvhGserLv7N
jkIOGLGrciaHCDSpA93UKR/sE3AR1QuuQOexuWN3BnDPCce0UDMAzr3QK6qhW/z5RnB9b4EJ2/Fu
3kbwEZC8TxVmr1g3nvMMlWL9e/Oisx5iQ22MWaDjsR6m4JMVv8On0wxH7yxRE/4tzs19y+URLYXf
3i72SxyDLUf821wvl6Ml5YalkRCvEwXmjTqLJl7L+lYrLrDv1Ikwsf+BwDeVKPvTptGhVfuu8VRo
H+d8pXjS7GcAdTVp/88U+dob2WDRUBPkoVeyU8JDKVLzNTiNE1mU80T0u9YZaa0/Aozfg3oX07KO
NQQQi9AwodWrA5WYRoX4I50zoRA+YSTnWxj/Evtml5dgiunxGSbRR6qMYzwexDR4ZuqM6vM/nDgy
wTik3bObXib9cVNkQohhPpH0XQ0lHb01ojtmokt4yWBPM8AXQk+5sCVP5iqdBlO0ZLHoHgB3bEx/
MhDXOhh6uLF/nVRRZrAG0ssysGlZS2JdiUTIMGqeRo8tRydefiBFBF8EbeW8yx2amyJzlz1kJwRX
oWZuMSf1YDLLOwX9SoRLvd0ovHyIURFG0zSnHYn5iYirZGtwmp+CAoM2ZXSbZPOLAniex67OWXnh
f4wv7N0hASAs//tWcp/9WkD3CwjpQiqKim8dP/bFQVFpLwtHid+5nD4NAZYoR3TmSududf4tVi5O
Z1NIC2QzI6gdtOHSt+QWuVtX3hAsUVc/d3suBbCgH/luvAWxMm0ZWsxQyq//SJuRmxpQSgtj3pJ8
T2EO2fQeSbPCI7n8GOKZtw2YloEmBvy64SC2FR8jseCOxh6PHLS+Lh0RZkXvhH0sR5yOnaRsy19g
2nI4hKuTTZZUjEGq/ipNKDkiEvzEWmBE8TDqA5LvUDNHSwQWGt3BBdt4vOudFaIHIX/LStxYaRK8
BpLrydtAV9++HSK8Sj61Y094B+szkhWY9a3prZpawvw/s3L5IoYuuBYN5DS/z+bocuH/UyGXDNyb
ZoyrlBe2/LVJF45gKwDtAkvTcEyAxsZbIgsUjtmr0sDMBI/7TANDZvI8BC3w1drnqUlUJMWv3kPq
nvlWSHvcaLTkraijfn3tW3eOVEmPmGV/VJSsFOAZIwmBbybdokf6jR+plC+6s1m77H/OKPCccXdh
e4NMRGj/G2npd3Umemvj3Wp0Zjn0g0JeSTypyyjcixhcbhEhbKJGx2tOMIR5w2LC5uqM20gYGsDP
WIERfSCmKsDPn9iD0/eOkt3Z1m8yunc4qVm3LGIXv7uCsW7xhhpL6d2dIqICjVwc7wUL3O019Fk8
BMaKYoYFJ6M05szNDYr4YvgXR7J6wIC+9Rqq30/YwalJaQXtlQSdPU1N2k4cccl0kS4Sz5q5WqUA
vPo8nacbsMICbIYjniK20Jjs+7KhJv0bN9x3Nuoa4R52Mz22S9dnxJDKwpI5vdGtYwKV4j4+VnKI
3Cjogk6s/xEk55+53OjVVSP0bczvVHynhweb2Nl8aEZUqggS5dEwLGJWIyfqzzW0W/OJ+XzSbCF8
liCL5w9xPVm6+W8oLBWuR8gxCiCEibsYBV6EobRKNAnFlZJt7LG/6aQdfksk3/HWO8wDCoF3026i
xWvHvAV9KBd7oCfaEGHfzQf+U9lcqtJu7SjUsnU32b8Wj9MZX0T9mSDGStSWIIkroOcA548UMq2f
sYvJKNVitV2jKM8bVaciQBFvAe0GZl1VL/5XCVIQf5kqDcKAZOQBiBgKEMqhZc/k2yHk6zEC3j/c
KznPN33RuNWIjXhInduLxi3yZgdum4aT4A73TlIsXiV7r43WJpMxMO40N1HtHsHRa2Z24Thraf2P
T0h7yGPVylU/yCFYX0/Hjdd9GOpVUPh7LEVZ6hiOHj/LdW5xWwxrcPWLbOZs1QnlAkDdduIZkBCC
0yulgi+4lwOUcJ57Q5SKpp6KsEnEmJIVkIZ/Vz3gz2iat3A5gyEf5KtY6o8B8Wy20U9T51vbNfEf
CARXI/ZYInQww2fi2XWWx/hvJalJV3iqHoAG3KXpgtZrNClVcoHFlOyxcoHHLz/apHUWAqYgObgw
5+N6Gw8MaNu5AkX79J8Uu6jr/tY1cnfHisclixZO289xitC7jrW4Mggh9uHejKY8Lf0Ci868ayha
FZMJRACCuyV2hqYzqEE5d22eEfjnSayECcqmeBO6rdqq23SMua5IjOuDumMohChdtkFTGQAd3Ixa
BMFdRXmtEl0O2laptSILtqJEga0ZvoUs6/EXvHNwbp/PsXqDjF5oUMFiDRPrFamE/kudiOHMIdg+
uLxsJ430xSpQ1HcipQmv1dXO+77qc2fL0UbOAeMbOmDiZWTdJxWI1ANQlvZGp5yIodcS0LYAJkr1
h1716zfn6DCIpaqWXkjnjhpogIrQD7nxKl+BA/ewu4J2lMgRwsQ5bL3KUfmXUX1Ws67JO7xai4D0
1SAu0KDQboPVQTvAD0TIZRbEsYMgsxRyJrLmRBuppvMyyRECBkuqdyGz58EY6IHM1ag31dSf6748
24dsfaBjgFT1Ja18iJWx4vzaEWgo5s5kvyQzGDPA0W/9vvYZNKECAonbkLNPq203bppIvkKqPM2L
VM/+CpzXD9jzLQGMrDVGsV9BQtVnLp00id+Hj1eyIhZisnNEqzGHc62dx2m1l+D9QsX/5FpKgsej
9ORDf4Q/tUOtj88K45yrLpBmxLq8+Sd14vXVm49cPS8QvQsTLUqYO74tKMdyggd4xtFZH5HWr+GQ
iRrTrG3364Ryh3g1rIL5HzU+iHOKV5MOH4HfiFdvT4+rXFx2oEoiV5jf/kdhb4YYWlSwC3x8dA3C
OJ3PKwFi4DTKAhiBhlLEeHiVkzOc1SSw/fwq45UuqzJg0AaStHM/Q2JH3Eg/lOZddRKZa2kWTPvv
R2pvMpdbDQNuBAtuZ26X7XeVhfyG4CqAEnvvj5H7YIf3L5zb5dlrFhZEbgjjWZlRix5aGGTcDDVb
JMNbX6fjWd2rynYvRbrdBWvuOldWRPf23iObHXevzSPbw5rqkNAEFmJNtGfg0XROmr3TWBX267bt
UU4oWgUik9WbN9JeCHJ/TaNod8JUJePjLSORjZwgstY7/s7zVwgCeXM/VxiwOh0uLqCAATbcD5At
1Rg98+xDrhJypU1/+Au2vSyGH3U2F8WkGdC+oEzFIAFhOsuaVeeNT2b1u4GGLpfkWxWNMXZfMQLA
CcWwYR2IUvUH+mknOUw9Df/GSqKFkUSmQXUH1aEYlLGQLS+2sEeZsuxI9sQuiHzuiAacl5rB8A7K
cI6ZFK7+VaghO11IhQIapjIPJey/caN1L0fcHrtEN065W95th6mDudR0lmqOkHsqRvDxFZFpDOWE
Buv41TE8noNVBEV+x3HiqZikdOH1nXtLMUf1LyzkkmflnwNmyL2Uumq1hz/oHeUiHZbz7QJiHpFL
bYm4nGiGpd5wsdvREUmiqOmDXmuIgjyyfPhuWCDU6r4OvZ+8GuEoCcRvvpZnqsHKJL8a1ezZUM6G
lnMM5uFdVXZeUNGKdG+nikgPC7gcX/56FmwRiJ8S2LZjmHG0UcA+3F5snG4X4df9typZlP3+s5ww
n/u8G4xn1/PlkJ7Enf+B1e/lxOH5DAe9nM6h1HwjiR8ASkrgnqT9531ricYAWahK4Kt2xQ8zCvMs
g6IoSUEjh6RH6c3LjDT4Vuh8Emcyo2JKjAGdLCFex3FcOkBV3qU+UtcvMVUq6KgXlEW6B2vPaEz0
sohS4lXqTAngEc7JegExvxehPoyW3wUh6JwzvASjwj19OmhaxOy6hf/zUyWSNR5jFNjvedtYtXYV
V4VPhUhmIji8XOzaK5Gv7OHU82H0eVd9CwHk3jDxRBj3wtiH1Y/x2kf5/b2FJNcRQGXkNeFWmHyz
4sJlZchGhum8K1nWoP80YW0VYacFtXknRzMJ9qPdLpyWCSrW8/0YD4RtFBNCShuyQMpMFrefm9ic
LtEao3XU55LP02hukk7ck4qzCbtFZiFrWGCDiD6bRCGjE9S2rPXlR/aNnqMVgQSwTm8KdC7boDjG
JXG6rdBNP+6V30eauL5lvi5iSJJhXN7F8Xy/zBQgmXghQrPyheBvlj4wqRPMrBrOI25e8EXjHHSh
NKmqUnSbLIzC5+Xd3903cRwOvrC68vQRBydczECXyP62KUvdenBpeXI2wA83xs+zIHgrjfo2Wkf7
XRsT5Lobme2uHa5MsfZiC4MU8RWuxtElcJQ6QnVFBmK1Ge4jeZiqgbVTXo1aRGSTK9xiSfSy+79x
7hXonVqg7qA+8Fau/uUMV8f1/RFrLFkDJWmgYYqc17uEgpgwodDUT76YOI9bZ/8zeUGYb/EahqeR
mocL3aZOTzQD0jYUEXEA1P8U/XDgP3fnO9XO/AznsXvGNFqT5s5qq5UPKKOgGjjQ3TatefttD0jZ
s+EAdBCjSjWsW3HTnRcqKxiSEYU3jCiMDHk8DQPZSf59BrX9Xv2pBbs2E7B0m23WLWi3f/HzVBv2
tZ+5eshCfkWJy6JyV9S+o6eJncUshZPEvkJ8LVolKe4xrr0OTOmq1PcHohfEeSsybK5uQ+JNtKP9
b9jOln0dLFOO/TPcNrwPFXKubwX/rlgzC94jPDDwugLV0opX8M1fRcYGZ1FsTmx/WMPl3EwCGseS
zajRZ+0kZNA4tXa+z7sAt1ksWHhjh7JEuODdZZnWIN4D9l9A2isEhQtlgfBukpOhWBj6pYWXNjYb
CD3NEwQ4Dh8VXDQdtGZAcl41Y1ECdJGjkk1eq20CNHA1vcxP8sOSr/cY2gvWinQl+R7tgKPPlho1
o2IIBb6h8foTU4q18KjsgYQ82JZHsYSSnCYUCZrw8YXq22i2hVM3ZgvHXu60/0G/7f7QMEaR6MgB
V+TGZWtKQ8X/gv/oas5EpEwkKgFiC1S+nGyJnptn4g0gNR/bPTinLfqIk6RKVasibjg8rFrM++83
CTEcMnfHfVZ+XUhoTeoEKS0SpToZ+a8jhgyfEui9pCRMw1ZRxMtpLOdF5roImj7EhlLd/ZQmSmEF
uf71/Rvgk4V/ypLMWkjNeNtA8BY1TbYbnHmenxnbTIZziA678IkSMBMKhOY3Z9X4GxW+7sx0TxxG
zf9c11dMaOJvtHJfR8au5SFUgEt5VhUx44DSd6cAU24f+qqGIsgn2xomvuWsS8fjHKFi3k+Jn4FB
K9UlRnCREnW56ojdfMtfeDf8Vlidxon6O4Vg+LeD809X+xBvqiJd9Q+3vyz1WC+iL1k+v1zZPXIg
gPP1A//BJ83f+EhnhnWtDyaDHsWY9/KFiW9NzY8aNxOoYf8G0oh/AEGkeb3xlZ2sTjOPhnzTFvtI
vg0PNZ8bOyy4sFyMVbG0ThMrR2GWd2xhDwA0LLWWY9gdu27CGfoOVVjumfp9OzYGOPWj9CMB+ePo
DahzcXsulEU+DBFBorEoL2CYpK6aCTgVwXtTquX+NKjxVLaknacpNZXFI5ceZT+RvrtGNEHGC2V8
ZoqgYeibE2wZonz6wFgF3V2T5aP7AO2XdbtduARfDyOEj/g9kpZdentR9YjNOIDhxfeO3hSpyasJ
XBbsKswcbpq0NKqug1zbZJCYAAM+kdWFnpzmh7AgZ6kuQTR+bEW84sMEI5relpO5AWSzZH5L8iIM
CVJ/yDJbIcz7PSDtVqDepUwjLREHMxApoNCg8HmdrvKOChoXJAcUbJEQ7CXsfflQMPeaMXNxSZSj
77AU1SoSlWGOJ6s5TExSsb1l8b9vF4jB7CdfCvKjBUR33t0BpaPTrt8ulW4Np56+VZ2/nI+0rF4w
c1DNR4tKDsLMD82PVpiA/N9NCzW3yFcQJBWQE8W9W+f/j+bXx6Ei596K3zE+M2/Z9GtwhX57wqKK
byyfKlYyQJ9qmF6UHalFulAeRGDc1D41XnkvIGZ9wyeHEcrliQVDp/3jAfGZfKmQ8hBeQzFb+KYA
4gSpuS6irw74XS8JxHyAY8AdRfx0P3anr8u39t1mCU0Y/nTrCH3By18B/KziYqXlbjXw9IhyoBLp
tWE8I6c5EqzGzoNM+yaNsEjR7u2WzIEJ/LO+Q3z9Xll3vB/Dk249jHbWuA+yKKjxDDIvJNNvXGmB
AHCepcSNN7D9XVn8jlVF77NACYja+dKWxnJPsLJDuL1g0eu0TJt7KUt+IBFV6psIP1ivIzGwQ9xK
RBWriZlkFuqYJac6wP3Sf2GOXDVqbvJu54VStei6DROPaDddkNTS39IUYBNLdMz6Qy6cdr2d8I8d
Bh3gPt2vd0LTYuPfv1NY/fb/dBjHl/n67X8JoqYhjsQ0qIfrkEax+4q4vFkA92gvIfnJnJ0CoTJU
8O7YFxmKayBJvvJZUyd7T7xV5gH9iowS2jQi1SkVYKjgIpSf0kO4dLsWDVTBbcQTL6i0wDNokDpy
IymhSTENd4mVLq1bCXqQUg88KGKyTUQLlEKdftuJlYxQTWEVqeiy/BemI0rVraASgFrpJ3Aj75OZ
QujENbR/jQlg02KnJWuC9Pc5pzHxKAHjRf6izJ/qMhDnJa0y45U7N2BpHEhb7qF7P4CNM9/p5tHW
2Ksx5TL3OOQAvXhuPq8wh+sV3xjkD8c81ECvYFYUpnc1KK7Osg7kA5mFnJWCsWw8rrvOnWYDepkC
5kd+qNw/r9TybL1eNeeC//7ECt+ocAYUwZ8bA/PTgKegjBiS1+xUV76/o0NHrgBoorLhLq8oxPYr
ZqVaQ6LrIFkdLT2GDAU63LGu+7KV+ueWWT06DrR270UokyUskQ5RVZ92betFSH3BK5K1P0bjEJl/
rd0jEo7HaC/XEakz0EMUexW2xHxzxRCe2dQMXxdJcm259qKGYDaFf4D5L45ULxRVllcQ+ShOAUr4
ZfER5ci7dhUTZ9omHV2WQgjfI2i7xLJtbpg/NvvGoGvNc98YvnjlpkvQiewCmqPgtqrtNK07jFGX
eFY8wukbPqaLixCjSuaV8VRRA/yv6gBJ+W1lWEy+3+sW9zQc0Cpiev2hbvGDlv2GZheHTJsRIilT
HAXarTCbO/AMIze0YeBi7oGsm+6wEt4saXeRYIj6wdVNEJknKTufe3pWbCsPcTMfNZAEbLiwekNi
/pQenj3/yof2gMNrAXxdaRZi9bWHzzyyEestER9w5yu2gRL57b41ZX1P/reCPYOtF1P6jMakowHR
1IFy+pnBLnMTK/r3Kry8NlxWpjIJrugQ5koDhuy4I3ngTEhJLVwqYXGBKpGGUOCRwJq5MC7x1/aU
THpwJYWHHCH/yQ35CjaV9JhVVGas6C9GwtAsibQVjgiffRRcRCM+M9Bs+1mQLEtQW8iNHiIxB0S5
OpCR8mcYNvs4Vck6Xf14ghXNIF7aw2p5t4fAY/wlL0U6HPSqR2lEd21OI58AkOT5sIkP3eKEPFSP
F4KElc/zKTnZRoEA1AHAESVm9SU8OgKQx6X8yjBRMtGcLszNzmxNcDEuAAEXCgnVjXI1CaCcYFth
/xajO7uY4ni29BJHot9bRIYWecydB+MGGdkWUFOPNuy4HqxOaKzmYmkAcXD05/93tNDuIvU/q7Sw
4a3kpX9fG4wNpKZ+GL9UeXhxl9BQ5rmDSE2A4RHbCAA2wPKzz6WUaYEymyRg55Gs/3alXhMpn572
+FciehviGwSKke2XXZp1kkR6GX4VzojVrCYIsQemhuN/SjriLB3UUGUWhprh1LDoRJ94NhkxlD3C
dMfFKmbHTVVggaA5iydXDHGzwAKZ7cu2AVMrJdJ1kiFPcbNdR1ELsHhUXnIEEDMtLTbgnSjYOfgW
CP3GL0SNs5zrez5hNBzO618qT4zL3RG93hAOpJqFtaP+BrQrsI1Fnbkin+TG+ySKirlJACEas7x3
wt3toNglTak2wEcK2BIWtaQVQzeyazd9a8SUiPuyISi5tiZE6Kw2GoFSVzISiyxE5CVI/1Ot/Nun
ZtHjEt7Wljy1Txr6M6ZDmZx107aLBTqnIwqWVy5zbo5331V9Y2taRqzLC9IteFxcHJuR0Nb/OOQc
giTK4GxK6fWOHpAA3LGuZXNJjO1ZhGvoMepJ90at7BvP/rPNT1kHo+w+0BKxvf9Xcrd1JCNABsih
EesYwO69eZUZu1m2Q/31bEWPHugJLnot29n41NBzp0UozUs/gpZX7l8Z9ttJ6pRkMYpoh5cvVXBR
xXvk7iXXt9CBZ8kKbfKmjukfixFAdzgA70SQi+jR2YOAqGjFKkGN/rRntMExIaCUaGTXhepjgcsL
hhMZN32/TTPrQvY7IjCjRzSBEJ8MDOfHQRnAbe5CiExtOl+l7Dsu7onFNdAaJlyC/GQppOM28MiJ
5xoLYHSfhkj36Bc206hq6bnU/aPZOYHspcgA1xHSPSRkTMcsTFfz6eoud74h8feN22KhYtqBzB+t
9j2u/BJmX+5nyZn+hCG2zdnbHKA6gVRdd+m5VR8OHG0mUZzhJ12S7uzeDpNbL8TBV3Of0y4ztZYO
TnNSXMJaVNu1dc81GBwvTxgptW6ezTMDjbRUKcn3ajv3Oe4koh/bCopKiM0umQghYRqhTb03Juuv
DA0NbZUIcQj9Wv4XFexq6X9Cj1zEZtjvx5HU/zd7p3/sr8O2VJf1OuBIIXQ0vDPsYSZ459vrNtmA
SQ6up9tp7FNEIwULqtwXqlVNydRBirK9pit6deXt8f0ym7zMiPRd2dLj4oT/SLF62HGGB+AF1mb3
J7nIWnfRmqtiMZfRoM/dt/KXm9DimKilEEBwdAai/nuMI/hmd2cFrqNgDzb3qM/2wGbP0OYjZAh3
rR0D0ClhFJGSvIz9LUbppGCaAcybrxvgZ/i52DUthc4Bm7syxei7RHp1XNMpcAHLwwtErk1UBbhB
TdaKghc6e+K/4UWKbrGUcHVZXOSgG+Zsip6VH/wfNKPgi2r2y8TgX9DzPiDJdRJY5Nq/EZTmf9zV
1pRcEna/a4b7lGuLvEVSipUyXgzgDk/jw/XAMt/Y4g1wLnnoVjxV74422oeLLtHc/eTzKbMpJP6P
u8Hpn0qQOR6fPOEpgNi6GL4hmqwbGfOfWcixGDPIR3KPDMDqqAw66OEeiabUHT6UYE9yKH5Q7c9M
HScSaoCgtHANYp2r5q6Fd1ImVR9jRsLJIr9Q9ZW8RMoGt6KCju0Y3luWcKB7VtPKL9Z5fLWUqINZ
1OChR9iZgzu5OTYdK51UxH9jR8cDLHVo3ZSY94ROHRjt2RhmlUbVOoWstkMBLNE/Tsdy7xgIQPI+
BwawOJLVoTDzIfjFA+HyJBE+2DND8d2IZddFZ21tqYCWw8QkD2CqTUU4QKfArAGtGcAb47yrbn9m
QYztr++u2QesFavnk6pP/y3y/s4T3FIlxQRCG5ceZrcVIeNLBzcteFYKtaSwtWd+sWg87mtKJGav
Cahz9AlcvXEFZvkUI8jYrqxkLbNeCAkl8CkhHWeggWJxyXML8qNggwF6u2jMyo3JpM4/MEJKaHpI
IOIf2kF8Jz30auW+cVBrsFWx7wmrJZsLMmV3hogduX43ZHVkU+nvYmQlDyxv501csOQHc3CklEd9
pZ3+pxqYcmYQqF/RiytWTmOk3YZvznbt6mEwKWqj3akoVhdimS5uJkde+M4WU9AYet2YQwFHxUpU
i5rpZJwU+aS2KMm2pNkR3lmcHrKWbTP2CdaUg6h+21BoH7zfTs+p29VZpQkqiOqCfSFJjDd3llF/
GyV81W61rY1MDNMIvsMGzSPzx+km2Ak/4CHGpHSYL868ofn7acafpiXsfc+6VsufgNwZ6xsERR7g
L87EwpilvtKvvmv4xNvS7e6dueqbm4dZBhEjeu8X5tipjUH+OFLaiWrD//WxvpzQEPjEU+UJ3yZm
CXD+SKq+093um7vQCND6hqEWlmYNsKd31OzfnKCqE2UG/UjWBCCCD/D6ZsC84dB+NDy5tbCv5qeH
OIHqiIs+Tkdm5hVVXN1ysyj24hUle5iHqm3XlEDQ7lUtrTpFJp9zpxxqmCTMF1NqJrGAH+7xC8zQ
gzdSS9ceAIk3I0zs4GrdmIKdDRc4lhQCIvEFN3dpa2nNQCXKlB7EjOsZNWPlepJFYGNReWtCsUVL
06yC0D5orUwv9Jy+l+tYPLiUAb+mMOJPLSDuJcLGIaP/6ygwG4hh6WMtGIsX3jab3iek/H7YInGi
wxepL8Hh9pfrsoVzpUDCsoyQtBv3soiYL5Fvdq7FRwXC6eypTVu7MRyytzPBIedHSN9R+EXnfUXR
jqeSL/tGBJsol1MW3GMxu6Jj9toQC3B+xF9P5ndn9lc72Rkpe+yYj2Y0+23QVvX0iwZk/xMOmhXE
PaIObSxuHTbfjwSy2pVyvJ/LvU2BqCkD1/Mb3jEsenP45bggq6jgdCd2l2j19goeNJkSxg2Rkh0h
6bn1Cn1wtYgbIC0z3+IGqEiDTpaTYSStFFZuY3wUlE0ntZPxvIcYjl5twXbIbKZ/11KyGx9rXlI7
bgym8FH07JbBeBZlG8cPtCBV9vhHY6SVPLK04CAscXlt9x9uUIEjOcrElKJouHWDJSKdrd2J+Uqd
HOZKfpJtXE2Z+cyS/3ywqn5iWEzmoAnN6jKpbG6tDMFGqZXYqsD0LRlvVlhp4QYha6aM1I01Zspe
3T9L6+FG5qJFMJysHWCQvBDbFdiJs/MOqomisAUOwzmo89p6ab/hTwH+57i+x/68/mZ2YuO7SAJX
idiZ9+jcMDtfxsGfQQbvAMi/hzDOOLSieE0Nub2AZB+yZxu/du3uZgZQPsJDSxs0+0sA4cuH1sy8
KXUbwC19mEDBRNrbxEpM9GlDk62GkHfquipF0Weyykv5tKH9EHX7/YnKctNXcMyd0um7FLGLmloU
rPB1sLYZtF7tbYWFxm1vhNQiRlzD/g660f/Pky2XbLKvd9S78/lwCYIKI/rICKybBDvOhLSZwC13
g/LGAYxDsE+0wvbS/OIAC8cu1g90FRfd2NIUvuaKPmp7dP65/YH/k9Tf7SkBzI6Yjbnsa+liR+AN
Pp+sc+s4oRcAI35jA/t1b7RpGO4F2tDAGE3dt6qautQjeoUxbl2SU0GHuhQV3vY2l4gfT7RIt0v2
SAGZxCmfT5NYeX4Qo47182qeIPGTXFgcBJWWJK6lAxDe3QdcqSFcoCv1AlX0nlrs/FBEARHaSq0J
d2U1MNsUzKP7H3MrqOdvo4RJhMZxoRrtYj/u96gxezJi/Ru27nsySIhNG0Aa+hkwrXt9fyuUbxLc
sgRfGJyaF8d6q2cOngZVK1T4nLdct03q6brneIWJUy+Pjj/myKXL6YH53MzrSkVTnCng1JUW0Xpa
cE0hf9Yu+Yj4VWIx9+uheKlta22EceV/pk01iONHeAvy5ifxyXgsXVdYk2iXN26ajK+aSFKXJ0jp
2UHYBkdfbuYfmvRroeFXYID9s5Pco1ZQst4wyM1LeuAlxNJGQf0W4ooaDwxFf6ob4i2SI2ICu4J1
j9Fflq6+Fqptwuc1S26m5T+iv7cBKfNyDCLEQdEfLksFspXxqvrXwuE4fVntV3h0ywNmCR1lEycT
ez+uNRnOeKjWlIlXbxzfmW4z684992fWo1xXk7BygvwhO4xSSQT7MUn2i6qjo0gXSSvPNKhRINTw
vPvpBpfRC2YAdAwZWtNYhH1VUE4+ufXwh0LgblmRzAoMgr8LhENGSfeb3xSl/edV+1oMzmC7zKFd
4MR49slXzfSIQheh/yl5JBWslHy/J/g6jHlDgF/uw69te+VT7WC88BMCVXagGc3w5gSSqZylyvQ2
tB3nsvYojxDCPKy56/bR9ROmbe4Gk0b3QbR2OtFuaXHuvW/ycX74imFvOCeF2SiTEm4bqMUmUhYV
cEALqOFK5dLzgWiY4A46R398t9uNCdXolC8i/0wEopc55zoKAXxmmO+/tBFpJVBKXKDDrrH1X7qI
5VQ6UuS7HW1kfc6qToW+YE4/ycXB7I7spp10SPc54sVc1OKDPiE9rad/hPLhFZOeIXM8bnTOA4aN
Ra/EYC2aXrkUwASqhcKLcR3IeYhBJIBvWvfzqDkqbUiXTB35mmA1nZQdNU3rCsWJRuIskJaT47/r
P8upAMwJvPybPGhqSLCO3Czgkzg8PfqUzyLeTBlyOq6ITFZ2WRpBw32jbi80CuTcfzH7+bibz2E5
QmCOv+HHrtVGtj/iCQhRKSOaSFljitfnp42eqp8HZMT5rv2wIHn0vXytjzO5x5jG8gwy3jKAUTiZ
5uT74jpwpnA+aGrFmj5VLhU0tTHn6XnifT3KpWaARz5yNgGSkN/bCw20F9risHJ8HjbLCNkWA+Uv
07c2DnGVsAMuCh3gwfJ5H2iVnJgfdErcy+GSAjEA27sq9LSkWDSkFjk5D6meRhOi3gx0/p/BlZjm
srKAaRj41NDCuw+xK12YVZwL3Njgm78EydSJBoyy1/bNk2zPefERnGIP2lHb8CYZaHqkGhNfEPr2
6jaa2bfhv7fbE83CExfsjdfC3UedEu7nrzmT1wBuZ+x9D/M4m8xbotGTEQMYeFREwBAyIcEWP/8G
oKPE9gRhxYDRldK3DzUsBBYwA2FRduiwfe2T7ngEEE5e9r0axikwWzndfeG3MXSpE4FKMvhKTX5p
pWFVyj9zl5hUc2rIB1MRsadQKdcfyj1YNu1NdutLNOWJLvb98GKsSYCL//1Gs0ZCKF/ekh4uDPyS
O6NHfmBh5/oGNmcqKRJtnh08NP3qUJLQTzHq10R3tQJFWOkBTERdprIsos8EvqFT8+s4uT7igULu
t9IXwSxoK+NPLVt1XDZtLx2JuyhF6pqI+N5PST2hZ4OP5NmCnhoRgcK7dyUtsG5Kota3JAswisUk
xdpCBtp2O2RKbrDxDoSJDC+q44qPNPnnMs6Q3Rpc+2NImmYr8awuJbaGwHyCTxUWSjhIdOdhB1ec
lE3qek4sGzCq5f5rcfKAKJrk58yZNaz/OqzZWE0DARqt/ewYb4pd2xheDxjgVCzOfTVE8uSIJOue
ieKLARUiz3A8mgp9oe70tUFFPI4NMxg4UQUF+q64qp7ugFLzKZv/+NOJLbsw6oNOgPgOqJFQulLX
C0CHpz+H3f1wxxmXoJ6w9X6eJr/AQ/9J2VS6olfOHJcSa1d5yUEbJM7hdWXjUNPQGPrJ4nd1w2Cl
WsaJe3hPC+gxWpoz9MhfRVsxwrCjlfAre16QWrqlMQy6YJDokKK51d2rb41/NydUNeVRY453zZO2
hJGNiFeCb1zSApUwDAUG4wXXBnOpjKl5x6EERztSW/x4eTHo5Ls0bNCBlwRWR2+Sb2LBL3D6ZuZr
csZBh2s7lhdDGijhyKjcQfn9eV3E84D0+7ye/fGgWw4J+gyPkEzbeX1sxXP/xC4bqAKFejQ7m6CO
70lJXQj3oMjh+J8V/piI06LASTLnpG7ElRp1/2aBvAxr1F4XrgllIZyIPgwuLkDCiH+eKKGkXfEf
HC0lxrE9ov+PtSOBH030Tu7c05LbhNRMeAvMSI64W6+DN3ZIz9v4sQI1CninVbOrux5mzIsIaUhf
10oUqVc449YRVU/xLwECdPgXeB2aHyIx8VTg4NDCcPQXNWgSmwXYmjJVUw6Rbu5TU7bkV1XW4Ytn
rwx4oa7WRd0oraafEgXGwzoxGQ73eGXiz5+xE2gkCvAIIzddPNMxv72gomkdruKc0CoY4CPha3rK
+O7GEEtX3goEldG5lwc8t3YYTEwYTzo6T72NjM1HDMdrqIWVzoeeYlWpYmhiadBos7ygzVdKz31+
D2zdj4nmsM9Fw9/tO3fknjmWZ/AN/WLi+DZHDlKOKXWawY4IIb7DvYFekw+O0vTiQTCBVKZ9nZos
s2LY/ydt4BwNbJTswBgX7+gP73B9lAED6ET3/KMruJZzQcg4DZyGflOZzRX12mCBid/uPVTGpnAV
9huT3mfGIJDa6CCDgXGeiHA6oIhM3/HJxJ6hWpxXcwfEtrhNMK/pwFg09U+U4Oc4vuVj7YvANLDm
TM2hOvMzfKGcZn1JexfftMCyHEoQpIaNVuD/FHEGxCJUjrbCsOvo08a3948WlQZgLLeshJQB9p6U
UvmSfr7G0bNee1e7qN51BuWT9KHhjzSUu8J8KNj8NPIrMVP9dIqIb2Mlh+fGSYAgCzwH6eavU4jK
PVYevxjVvqPu3QQ4juQ2PSmAY4iV1pBmfVFWKY9AkqJ1wbapBm4CCZAdxfqZJRCoHGo09caWzGKd
hMFjMU0XWL14qJAO+6MGOXjXkHHERtqi8YlHg1lxRhKUoZbr3r1OGE5msti0di3M4c3czb/L1Xmr
Nn7MZ0FeCFNlSFAA48N22DB/u4cNqnq5Pd/zyMzJCFM6Ro6g/vS7O26zQOugC7YKEq6RF0TT570G
VDpqr7MbOurl7NfG8KnhFirX4sMvYOTA9PCvHFykRYRo9ZDJgXK8e+qi03DzwTAU5f6ay+bMIRXK
fsTp3N8rMoaq2i2IeKAxUW6awtwucKbiv+/23xAo47ni+HvGnJZEa7fH/DGookXlXpGp36nCucpT
GOi0kWmG/npff/SlsFD00SAIbtJOOWM0NLPP/zm30yiphYz8ROueJc9xPxLDVzSFp/eWJ6iCrFej
xE/ERCZ+MSBHd5WSlrJKj0++i/XyuU4i/rAuzDyAZ6K593irJ7n7dNRWzHhtBQcmlyX6jYIdiWU0
yiruQaoLsr150PGB7L1IPbGeVqTbX9NlC2/5Pj18wLhK6uzJHj0y2GotxiX0vmprbsTppyykTUuK
qu3qkp7aYAaH/1Fjc1AE5g5fwWOqyKDHd6oXQ+Q2weIHjJaXjEXTktTpRUDNStSOt5CpkZgBbThn
MB3v3lsQZxEk6bXVwlnr2gx2VaHfQFexsrH0UXgOhfdY25770j9p/u2y3T+giZtKN1gHIZnk3GNy
pzbOe8mbERYuVA+IBUX7d5rvKQoWOFtHRSvHF4vj6vrvMtYxsQ5Hegyp4hKrbHjxpbm1urn3WMwA
wiFpcjSr2z58v+rVng7TvEFW9lKoAi0lA7x7RDJoLjEVZEbuILGdP6ZNSUMM6A1jYq+UjLNKL8Be
EIUJ+ZV0yHFqXijzLtEDityU0/Nvmlh70IOLtjd2ygEaOcdA46+OCwGiFReQWVai1TuZRekz4mlx
XEWx0iFiCaoQdxFjFTtbTZ4JXrd7+t/YMuhCkL7Fk2DM9TjLCJbrXHyp5aDHKJWgs43bzJdmscMB
caks22Md1HLzP3TDEcHPTt58aFeDskgdhS/XkDzEMkNxr615GLJKwl7qHtNFMVd0CUJY0GGObIpF
hsO9GfOPBRZ1IV5wR7dfil9WzYy+dislxWOxBSIjqM1rFJGwZ5+Kg1nrof1d+7a/h+0i9qI2+qPu
5/nkMVJskzhe7FID1E5obJaSkN+uarIOO5p2yDs7vbjbN3FnGN+XQMyC4dwcGfG8POx9zcH40yp1
LJobGN2Gb0iXvbI5oeyiZ8ptUuZgJzgVZi8pvKjjkm2M8Ga6/Ms/ZpeALdcCsb+vCBZC5ZpCqjxe
HtqNcwuwUvZZaScjcWRzqDlCBXCo2tjRogh1e/b3ekPXtpPzVQ+67Q8tJ/d2FFMlrZ3XGV5LaNCp
RmfSMDAkQpci/ZfO+Y4XH6/hsb2n5z3EbHdQnlZdK2qYShNfkztKn+Qq4VaQTFFYpNzbBIAIa5/L
Y8zZN+y5ikYetL8yImjZAWPF9V+qqQy54y9Xj7cxFm/bth/6KO6G6tGDawsh/RTzK/S0XGXxFbx5
T6SizohsonQwkibLzRXr5hsOwZ8vQpESyKR2MC4N3TLiPX8DEjZ5lLhqRi9KpOgzbaksrQsNpQfg
yGbzcPGColezoYdy8rMQEXe3ckyQTG+WK8SWIdqol3w7/goHXM+d32nYIOWT2pYrkkx8XrjyEzf1
BljJ060YRqfF28yYnWydGyER0DQUj82x8SxJ6Q8CTU0KwxynLFkZIPcQN/6agiAOMv3UjKAgzg0z
XNPK+MfFmovoRqD8v8+Rml4v3IXCzON+FXR9pJiivqP0ukoyDd0MfA53NpkKaTHicisPaJ1I4ifO
yiCCmyieZmTZJftXPq7+7HzMyWqvvyzRFt/ciDvHHJ0uv3GZu0ZvspEHsEfUNK73QC3uTZvZhWqW
d4IeB6mckLNam8bkY4ay06cWNTu2WgMVabiTKLF6a4+NegTtnV4znIvERGTbD116JXmng2HcH96T
KVEcFAwwa3qS2b/XhE6Gp3NCDlbo19F8mlEB0fOdBjEK5n0ySFExXM7DZ5RBbgkqgzOhNaQWqrHj
NqUUjAN0dVw39DA9h6uJtG0Eus8kEvIzdGBaTVA4MuLaw+pEver7LOsDiT7p5qUCS2oNQvmWNW2A
soS6h4Kr3nUkf2YYUsF/JwwUVywMq5H1iBtStEFK5OgsvxMXfhU4r8+CshvZ2O8GN3iA12emZV3V
I2+V5Nqm7lJ7LsAAxQBq5MQtMY/o7mFrUcjhvVSe2B2Flmo8tJmplVaL+Z2CdUtER3bNp5SuYVzn
v3eoqC0JaQZTcQBQ1yCWOy0gPagyTYI4BYvjNZDUjHllloiPHQ7nfvKs9dZSnwyhz2xkvpJDFU8F
JUFRjijOPwSU6oqqT1zLbLO3I59ox33zxveaL16dxB+tfo0kvaZeMoWbmoRheUkPxFb0BF9RtuzW
O5bYJZuxPGkeTwCjWkqxErwhgTrdp8JPopf3bLnlghIKlroTGlgXMM/EmBYI79rpt6RbuqXfmxHT
hjhw8We1ORedgFmp7T3nfxVcx2p49jbyFVZzK1ok8GmHSvTazXu8Tbh0Rlzc/rFnwZuV57O9FZf3
E1Akm3ziYX17KrhRnWluNPxEWksmNq+NSBf2qo7WtIZ74BFca+2vAumezTUGrCaXaHJ6AvElJCfv
eLegnBYWOBbTSKRjRUmxN71VlY6fk5ifaVKA1vJoOjA1DPXmOAHNIOuqpzvb/iqstJORv8+Hdivr
HT1e8REBiBuNJp8RW+QNLeShPQTYKpYGrwuhvN85YgNCCpoh1I+26nD2wBNAzeYJWdSYnlK6ZZ5N
TiOKKz/dzSnREdcjeqPhDL9IfGq0FCAR2wolo8yhTLQCQWdxb+LxKNw/Guw1QtFMTIOaCg4F2PiU
gjLZaoMtfbkV7d34/CU6IQ0BewTRUykohXn8Xl7Ds7UhykaGUMzm0o+uXjHFiq6sT3DagQtm0HGi
vWYOal1SPSGH6gKusVAT0xv2jXwMCHyMecuqa9wSDlVt1PsL2Aq+GXvswJk9B0XQ+RIwW1rn5UoT
lbzjLyPOKLtQufnNENOIqKQYG4HbnnMStdOWqiAomnIGJrojfQDM06c5OGO0wdc7hahXpdsGUTA4
hzjfLOpK8o6neC+qweRKlxMVrBEhUiMLFvZhocmx2sPH/HBHTB47jfvJdshnB1bLKQeVknPfRBZQ
ex+ZXe6/O65mRtTz+XwfpYInbYyc0BiLHICppLmaggrNR+EVpDnpQWU0megIiLrkVvgKZDwi2Jeq
oJzKEquebpRecVKP/pH0kdBDFZIGLppAiGKlGgQ1/4h/8Db9bKu12JgXGqkRX64ioaeOcZkzacrP
WrkosMwq17zjSXQNROzqYHeXRO7+tmTdE25jteyv4BICImgDJxG+KGNDMyQs7ERwaSkiIqht4ADR
wx9Io5kLGqObFqFiHulC+mdXcOawzueJwIwFVQsX0yU7sUfOJiK8G3kZd9qNEYtbXZga2jV3RZ34
fXnY/hvuB8+v1guWAL6P1tWQ5Dcg9BxDKN4Haxxki4Gn1X2pO/Urb1XFtYbEPpkhLouX052dh/06
ymQoD4PJ4UynhgilO4V2JYM8LYC1QKofwU1WpU0bp/SiL6M/GlgqXtSppFkuS/lpQ365AHYFKcrx
j/CXY4aif7TnSu/1nZT9lW7yZg4KQNUpnED6hGw8ncUNDQp0lxA9wYQsAseJm7AHGgLmU7/Be3XA
W8/uGmXPGKAGkYb4K1rx8pWxLoL10FD/JNNVOztjB1MGGuZmb/7mUl4/hsLZDJTPBwZPJ+fPBv/H
Sdby1UFpkqGXzPcTBB3QzGP4WXfivoSobSWWJin+zcpk7xmGsXQ/tLFRNefejO/+QfAIJy2E1pca
ZSsalom8mORcy9CT1D3N7g1V11HubrP3D3q2xKG2+ozGFreR3ANdH3uxTB9+/D+wjU1Bdn9Rh3MT
RgjFuACyswZ/ZIFS8hRMq1xZnTaL0VJV6depVgJiyEBcRb1OUvY/zyycGtSYlB51bVNURBYkQy4+
A45lxO85C1K8/sc1R3dhS6WmnBMcFzhb3agVcFR2f5Bxa+DB+8Xq8KZUzXVA6sz3ersKUkGMg3a5
Y7WnQ+BFb+GdvNkmnBdoKNIv7l+UQPU1qh1QFftesB8oiZiGgCV7e4SQ9grS+ibtJYoz9svlsqQ7
XcSFTfc+ZtJyk1c1EfuL71LUdaE9B92KPhrqSvDyNPMwxDA96chqgmybc5KpyJ8xEkV2dCw8RkuB
6q68SJurVHRtPMg2SXc89vnX7DaDL9LXNxR1nZ3iRqzPKpJup4UhwZ2yKfoL1qt70Um/xAkdfbMU
eHcb8Q15WwtiE3zgx+q10JEUT50CRa9wtQcyLaaAmqQU51CHUaIvHobO2ztfeFYyaPmRtYCmXcwO
+IjSEivmSFFUyGt388+J+K9sSZ8Etj+Sfg17HDoU8JTGhOkuQTlUiKSpwqMcnJkGWpnTbJG3g2G1
OgBCxY2t44foQ59qR4eQuLKwcRHQvIleTsgggQi3zGc7SF1S37p4UIGzFD3bd1JvnsD7N2LyyU1s
zz2navEwt2VLkcHu/tpaaafXaBp6ZSuTli2mpzYQGzZFlbXgRfHdlqx1+090m0/L6ltTy5Sa0k4W
WvjJkXhAmhM81R9+Ib0M/GG87E0HQ7hsNof+ran6JCDleoYYyFugCf7Fd2wCXWZVVnQfMoQTDC4u
EOVzF8n+DqcIijsiBNakuHaS2lGRjrdOsbvj7q1TW1lSfqYPv3uq0TNIpmGbEtXxp5X+VS0LQAZ0
hx2JzNA04pDkxMNgXH2TfCkeoevKhf11lB94FYGvaYnVPg5g7xsTCSfqBD7CekHPnGahfHU5tte9
FtnPuj+PjTDloA0Ih7iDrcYhcECn5JQeR35xU0g4PabIJr4j5UOJd45wjaMtAeVxxESxJdIza7Hi
SE12z8abzs9JWdgspczdfFyXb7fUSGei1FmHiQG7b9hGEh6Cum5eEkx2x0mSBdC6CvQKenYJtW8D
dAKOhPzOJdTbhWJuK1SAghBTp6kZpQw8YETjF9LCrNxWKeDFBHLALJyN6djR4XxLQm+NHBpx58fp
5bQec2Ve1mm1ZJZGmEBWQHB/rnCIgkCfa3e7xEaXRiEU4aRMOkq902fjr8VeDeZfRZGp9gGEWjYZ
wfU0UvNOw7SrZMgng/frUoHyVk3X0RTkbYoipR2ZUpWvE4OcEHVYwZuvTg3vUGFBSZwH984l5Q1e
6bc5DvJH3zGZWU1yWZlBzuELrYrz+qFMq36AOwuIBdhlMCPV6Z8s3h9Zlzc3q2++64nbtEaJoxHR
5T/zD5KJueZ3bu1xwm/3sLGYTXfv5WP01u4qAHVMEzjQKLBrJ11aZtBGIwZaiYRLZPpyq6xGBP/Y
Tea86ggAtxtbvizbVMxyKzrEKNwFbfAm368n47lHSHeIIuvoFmv97k/TaVs1YAFpoz/pNFpAr562
+zJKlqOyw8Dj8ewIYgxpuFJyfqSdFdIYLf/BW0nuaBQUCAoGshvLB6rGxD/hS6xgeDyM+GAmUEBz
uNkp9T+JARyFzhaAhf/Bdry7hen/CFGg51etG5+/Tq9/sbhcwH2o5PZYWafbx825fZ1dpGTJ0oLA
N/W+Tt/eTckJYxq10uyv9blMXVkPjqQPDcEFI61WKN7zj3vGKlrD5jQw2quYyviWMlEKTB9ZW48x
xjTzT6DsrH4wlPqC4pUjuUpBmDB3ed4n4m+JSestgQtxNeZo5gg5wVMBJ3wU3NB7yUKxtDFZeqL6
mAdhvUFyZRXLyxqX4rdj2+dhUP6jtQV602936qoQlXAt2gmubIDPyj6g0OX18inJvOmE9EdOTqJg
NBzmBFlMq6NBUdrUfqZwt2PwKD4KUHGyofmP0Cp67BQMMvq0/eWmHbpSWiJ0QXIhAxC2mwxCrbNf
i8/k6VP1PwsDrxHwEBwFuaXiCeK5WtWsaFRTlBg/b1xQc64j+KwBLsZsocWF47E6Ws6kCveoexz5
odaGVSR+z24lC/8Jjy/bD+kVBuHcajhz0upmoA8bBP/QRi82tprXr+QvIAbeLOt0HR4sUPupphl4
MONkzNUpG1lx1V2rBglBmhuUwJ7cPsjFq6Z2B7ffANhs3pOgUuNJK5EFF3S7rktF8ge6QFzCUkfW
RzHUJvdogwCzOMkd9BwM5j7rRJxLzEFqqmfn4iRgAncgxXDgMBQpTymrJNtQNdUY24W/hAiKlIMv
Krcsb70l9DrkklX6xgV60tnuMlM+N2pX5b6jW0RN3bb6TSBoB9+3b+/0ZZdY3SohjwJLq9QTfdEL
8dwRPTh/UR87NnhfwyQm27NOdlYhifqOHEGBWsfcHqyGFRIELR3ADqkF6HC8mAuS9RZSp+ZDmzHK
0E5TB1J8PuMNDJ4r79Ri+APpgALbZJ8IttslTGh2IbFBPKGz4dqry5oHhf1vXNfuqX6dCbtHC4V7
VnlO23kC36cyP0sqhhZVQ+HqEvQ66FqTOeEol6LeRkXopQvo/Fgi5Z2b5lu5ziUcO+Pm0om93erG
57xBpmPMN32tge0EgExGz13CflGvbwnbbPKu9rmMiidwXtretG+QTaFEx3Icr8vcy2TRTNyPoAMU
FGbG7BT4TDma8X5b5OZXuSgGzUY0WWLQ+GEtVaTthXAhg989njgxnKyRrSNsk59o/MnCJQDiN88/
MSOOU9gQCReP0UU7uwFqv8TTYmdXhI7lkb+ygRDnl9pdLKJUgLAvRHdtWVSOtdwiN+a74CSFECTT
2d6FKTGpkn/l4BDwz8saGI+pQcrC3e7E81FfiKeaeyxLPTzHbZW3oevm3LTkxMOOfAn43IbDKCqt
8d5WKrWEkLN+IzQE4rQZympxk5ZS8ahaEplm6SEnpQy/hfB4HUNRUkUJdAJP9XoCptr/iQ26T4x8
wT+cUUVk7BSzrdAS13mJQlHwa5MdVWrieEnI1bjkIUfHBu6i5QNMUKZBfRlS+FJU2yDsc/RVDBLO
q8AkNrfOtUmURZMbrOzxOQsTOWN/ig11sbYWf7cEBGoCxvcjvAeECwmfiOodGSRdcDqDR7BKZVIP
DkzdAUSYgfMubyebVO2ZyrLvkWugjEWFZOgcdo5pW7TMxUO8qvrifvGgUXD2Scpmg8mr81ixtMnn
1e5nRFjrYaMknF5R+0JgTSJSz72BidZYyJN5D1p15xCbkKHJ9oh2P8sZeclO2fqO8ssj+WRCWjw9
pn8hTrlET9lrJMIFbMnrJbrgbGUw+pU1C+UV+k3lW+b/BRerrJNKUbOom6Efvi5OrwYyrKd93sZG
98kZbrJ0OEODgvqsr/Rp5RYgKF2jgw3aWL9BEu8K0Whd8iMS+ypusnNo2jsafG1NAeLhXE7xAoJH
XlOzsNi22cOjMimzthckYzOq1pA890qpI3n2m3HUDS2DqpjEPBph5rDSEhgj09Nt4H8K/Y4I4KQo
SvximEEKpCGeQMnlqHTlmx/QDJaS2HUw8Eq7Q8Iyi30SdhyiNshjOUK7SYeI0d3NaYKefDKppNOp
dSc6Bjyhd/btvpNoBmTBPjQJkuKo2kQ02Cd6wOKv4drlXO9rWBZHx6UIFobJlitwLd2DmQwlgcdJ
DdEWtM0c3liDbP6oAlQPpeI18G3DBEHDgap+osVO1ejdBpuLjYGIPmzlw+FIor332pS2Qc15PFvC
BqIuPzuXb+/r8E0TjxrhSow8mnAwgZ8NDzS1tGgKSpmT/0DZDH7Vv5BR4R7khl9FxeK9Pxxyddhc
cvRGQ+pHDkQJTgoZ7AtbDlb93Z87CWsNTqehymga1/6i9pvrF3pk/4aJbkSiP7w6Ck9yD63Qj+9m
SQkMh/fzyRnVN/JKriOySUo0YwxY5MmwNbAxtlMTA3qH8KRIY1zxla3O+rweBZ1pa652fbcM/8Ig
d8FbLmXWjzRWLLO5BlEu2G2mziEUYDt3SsYc6njmVOq5YScO4DgUJOLicvaBxLZOGvnbR8ylxNOU
uGAsBD3USyksyEyWAiCPxXXyANX80RTdPqiRPCZQx94gf4jBSOKq2dRdF+DnjxWJFHF4zYWGfFi4
u9ZOqw+vZVdkv/2IlALTDXAnPDcJjbzDqAQqPuJLzzHL7N2s9cVLSvZuKb0HlqUt4RVuK1QnRyok
W37F9unOtXlNfRg2tg3/YT7hzgTDif6DXKp0/Hm4jRnf/1NH6u+1PGy4btQMP9qRFLONqEEwFqXq
BIH99AISGbpag75+bQaveT5PtzJ4oUOwgO17vOLOrdN+ngnnQ7xkm+v5rq9Bw8FCo/fPHxPm4p9J
Mh2cJqg5KARPD0uQLUt/RXDHjyO6Cl6Q5QeI5gScDjCF7f3fUm1yelfMRj61eWt1J/AT+xuyKgi/
St4ZHMw1Kgt3QZodPL7fYw0fRCbYGWhONULFJUSjcSU1vOVUm8n6gDNvR/SMANArP6s5Ogvr9VCI
3Wr41HLVpesAy5wh8z04u9IG1w2WUktSFAXT7hbhYntxEYww5OtG3GHYGW1u812X/IQ69nAAP63A
peEEruLXkYmfVNQbyR0mDnjF+Jqxng3EboY+cVDPErM/iekTA731qwqk2c6AHw8omcNP05QEb44n
DoknFhKKECmjIheV6cE+vkQ1cbQU3wOviDLhZFlPskYPW1R0NyERF+pti4uqtYc5M5j6+xLn9bhc
7Hk1x+0jLRVqfv/tRPMwL6fwyOOOBegU9/y6ZO2rT4anA6EwR+NNTVUg8P+obb45+l/QkGOfaZnQ
iFFNDAL5mzGjYuhsRPQYuGt+teRw1jtMWhsUx+6G0FEIbkFpLYYbbROK7B5IiBIVuiUG/n1auY6K
vzQc3hZLbTJeCfPJZZ5oy5GAeVZFnVPPE3/Wr2U4wEpCFowy7cJNZQ79cAQ3PCG7aRHFx5kXVh5X
AV9qbAS/rvHsn7hWijMYnhdI1ndVLyILd+P8n8uM/EnxT8m0IeECK6A6zsGA7uOnMsatsoR6pGkq
hnk8uRR2DKQTj/Zo2xLknkCFflSz5yiY1G9B1gqlUUni45VmRb97DQ8/7UQQO5vEwPJlpN8h4Tuh
7kQQ27JFm8wC9rCF7U8eiKvJGBZS6c9RKWm8uQaj6WLFq0u90V/So6ai+fZeLGT3gwMuzXlMv3vN
Zk1i8vLLFZLNGhUifN3PbhjsJCIO9gjowpV5IA904fTneQGkPh1y3mQu/5X3qmsj9bDuTXOLE7if
0TQ/GXMSt4z4g97T5wQ/DbMpEmSNpJf+bNYOBcQ8yfh8NlOESfOu9Zk9iLK6LAHsf6XhTD7/Is51
SrYmllyAqXXKuenB30bOg5tjIDGs6L4+XMDjGJa1S2Fr2gvvt4diFBv/VsitmGFARrANGpB+7UCw
ygm3Qh1Lcc3BeEXT7dSaOZsYNb+j8KTo0SwVgCip0xSfmqrz9CQwtX3MCA+AUbGF4ksCJy3y2v7e
x0d8vWa1iN34K6gh2aj86jBv521qnHxAaOnH/6KH4ItOOrtmQX/nB12vx3j78L9Em2fsftMEWLCc
AsuO/v/Uk+4tEYwZxxtOnHGw42DaXfjfS1e1p6ZbTitLOTYZf9nIrROo9Vf2WekXwETfa2eS1sPx
N95aAyIz7kGYzCjcPqqEvMvj4S/klYeSU2B7myHO2QY44HYQXbBnTUYK4jAsxdOmaGYkwoTMZyi7
V1OCxoFjqgTubAz53eIF9jR9n3FN+eBe3YR1+nrtK6NMJp1xuDdrsOqqmA24VSCjcYUQHYuFHP9G
VuHtLzeWXdYWoPEv3MYBMtWse8XkGzj2oodf22fQwndMb8NfLSbWG1dVXdGV5Kv3QGetN60u3iGV
NYhoD+X3bK4q29WWY/wmGlcdJuhG49RaksaIjyDKYBf8hY/KWkgkkbm3vQ8vfSJ+Ig1GrQcRIv5+
ilBkR2BnUu0c4VPygtkmnkaXlpNF/x0ySvH4IGtnwxph4y+CELIyUAuIWiBKumcboctE7bTua9Fz
yj21AsZV4OPsh/qUwGyajKSXqvM6+MMcg06QWzcJYs8+7zEq0O6L1n/WAC+G9Jt9UgoqczSBUtAk
RsbtqoQNls5h0UWqhT+kcloqaPU98HApe83Bmo7kadTy3F4PGbMmiNlvDlbq2lvMfKC302v4Fgfz
2IO3XoNl7DpReyvq4S9MhWNvJKJAN2v0udco8HcC2iX8i1ULY95WZEAVh0Ol8BDE7+O8iI8g9Cz1
9c9I2wioRlID0yPFd+U+mDZVgsMY1oUP5VE4Jv+270+OYF4hr+xDaTE+88z47JYFdy/kGPRloaex
Ph/SkcfEBIyGuzKTiSXdbcasw1gBC4Gds2jDejvKWquYISbhW03dTDeWM2Do3S3yKRDu7SmLgiGK
kxkXbAqvoIrl7iveVJBWktKxzZRup5eU/gRzUKWHmK6Zv7FsvDDGhRgzXsARgoxkP8mapUTla0Dn
sABlAKFDeJarpQvJOhg8lARYeyjff0UJa5sBMIi0VLM+xqN00WtLmBSyEvE7GPFhNgKhNBAEmVg8
x9uIz/TlDFBbwutvGSJ0olDi/W/AKsPHfmiAbnauyLssIeYuAgCpsS/Vfbub4FkgeriqDnP3YZzv
J6FGVcIpkzUTaQlBqokkZBj61azTnuTiNv2Rq5LT/iUv4Y20jTlcbJPjzmp1jsK03YLs1E+ihLl8
o/Hj7JR2rpOUBgimDWlWkrTUzuxsrVXfqok0eu+GSN1roJtj3emluSElf6M02wnc8F5S/ljBpXDs
yTf63QfaaSRpPETLBwRXvHPpmvQkCo6HhqABMe1xewoYwk+9lrl+5A4oRINJm6OEgbgqOCI9kyl2
hCVja1m9h9ZSTZ+MlxzYQRcGt1ESltmpP7pCPvDyVUkg9MxC8Ch2X5NEvH9oI20nKP8Fp43rc9D5
1sEnxXf49BdX/aL0jrmrqTGox54poPZYIfvMyebNc33FnJGHMhkLuV9T+CBczYYpfUsNMxVphKTa
6vcxjM6GjWGV1dTl4LrkPGwX+aLrpYFf2GUHIb6eElmQSapqCvqsOe5nFuyviDoywjj+zlz8Cutq
nRSzBo5SPINP5g6RsQglUYrdVXt40XLXHnkewHG/27h4oW1OduRLv9b2hg+VJxVLIp95jPePhl3i
I/KSc0OzPxLCMKFG5ik1qq4zFHdohCEAWc49icZpjZ7fXkpAoqD3nWbTrIxQtcH2mmjRTBXXSBsu
g3ptLQpRfWbSts6wGB/7hbKFuINtNCBGDW6NxR7nNsRkX1zSSjibCvZSTbssNoYq1/DKugz0g9zo
dcBI9gmobAZphlgh+HTcrOkIZofqDh+hlzXEfFUAazQpE1gH+jMC9dyrQbJWJyl/LLJAVIsm6yR+
55Y3go04pTE1G0A+m2/Nk8bwdJOecoFDXKlKBk7Pv4GVlWQIZzgBy0hB0TLLkFv3iTWY1Ahs9FDc
CaS22qyLGqgjPTPpUBjbGbxQvfaPl+g6gnV8baVyA5tZSvEfxponzOpgERhT4OM7TLSYjGZ9tM7P
gZTp6GCrA873v/OHW6RN225HKQjfoPyt/QetSfA9Oz53LN5qr4MK/tH5TEzk6L7+2cEOap0PRG8d
cDfvBUy9Gc2QbrypVHGG/SqwKECcy889v81XAT3RS5YyXWQ/XGZ07uaD+yo6zgPOsjjAAr7l5Xdk
tERn2TZ5dtA9ACzUsB8ufNh5igIsVWdkVDhHU3+aLumcFqPtqicCW4LYA2KrwGoAIYLKQw9UYpBx
YIzsN9VbPFmykSQpc0rgL5ue1BJLJyu4Z0Vt70oU6WEImBlE3Lzgl9sRD336W8/a/2UD2MEP1WEx
yzJ/2XQ+3Zjdv7ws1yjEpsXO0IabpmTQIOVYRsF2Ai1ys1/zFWfGyBRBpLNgsEL7EWtysMKb0pmr
VfcdipKUBM15Wpa1zrNNPSMBP3JeMF/VnrFmn0eSfa6myDhsjmDTliBqp99FzIVWSpWLaLzei/18
qFhacRyjaxJIrlH1MkOeQ3ucwVle2Ho9lYZitZdJOKIeWE7nN0FwBpAjb4ylZit4+QYj6SDJuiS6
t81FiBo8tEI11c7Icl7nYPy4AzRr7vkWdBaBzhSBGXRp1to0nKn8ZaW77+q2CGY//Qt6QOGdWcqJ
guTjdLlM6GkrLiMuKfSlfpGryqBttVVmV9pvdDbK21kvf3Q8EyzDKDKtCKvkfCzeEUXCuGXwidFg
x1F7YjMbSz+24k+Uz4gsadO8vGEQh+apU0ueXM9oo3zX/uvpIEri9bxbr/be26L3nkCG9fme0C8d
HGea7iCpkYdT6d1ohpnZIdbUDbpD+jvZMtJgs29pbVyr1oEfET9B/506bXyPwFzkLc73Bhs5NZC2
yv9KPxsFWkdLKyW/ezLEXuSKanlNMkr9zRjpSWJiuchL/LMzZ+2+krDD86/93MPOow0S/M9GhID6
gxRW/Za56mYG5LVWZ62lAcVFGCY0AyYJ8txUM3I94Po6qdocoqpxw/tipiparwh9zDbsztuxaAmF
wxMiUpbq4YgJe+7pYrPRHNgwPBpXYu3cY0K84vw3HLWUCjyOSVGGzo60zZMaKqx40e0QTg01pUnq
GqJ2DoNA5h3j2JhtHLkxgNdJU/uH9NqWTR/cLTOULrtRzVRm/V6ac5XvUK9u2UqEtmpRjmLLLPXN
IBI66HEjTd1Wc1W0LwkK/mAp+FuyjIVHfbghTR2p6UOtY5b8xKxwchnga9nDGGm2EKfUgqutcCr8
pVzYqkTX0v/VoJLDMPjteHgaRMY8gWR6JZYGTr7+30EfafaQIjLxwkAf1Tx+Vev8ou36f7Kz/2tW
dZ8o+NzXlUTibh6XU30WVeHOmpzNy6HbOwdEtxH2C/TAr+12xQuuz3KqOU0VoofXDEL3B1Cr4Pm/
bMqurcMIFExWqnfhYK7yz/t56/YriE1DFiQw86/IgsOd3cKSKMoXBiNohBQoKkqOLvotLs57RzbH
Ce50chZf6Vo4/lua23lJ/xMCmnYCvweqZRceCoy702+3FR66ERpYKHsA9EkmW1P07IpHFxs04cAa
miNxa911YzsCDBHF3XZ4YEzQn8PzQFSRAuCsZBnYsFK84ImktD4TY1/H5mWs8O1soNKpzWjLrj/i
SRaVNQMFnYO8ddgwcgVHVC9h/ByS5UHHsZPdGQVN2UA2Zo1mCC3FroJJnW5nsrjlXopHTgqefKNF
OMykCM2cuux5Uyt3pVDI7okVk0pEKRmc9cJGS3TlGO9jv8OrH3tfgl7/ZUWy3+QkZploT48MsGPf
kPqCgcjAVk+f2hzx6MpovInSbnO/HqKnOoNIMvw4/haccL7zbVIlpfFEAjReL5mAJVxu4oKA4CD8
VDisC+6Pui3yl7KhiXsLcVQuYKAJE8D5qmkMu2KFrsC/RaRqQLNmxvhTB/7uAJdXGBWLP3b1KUtm
L0HgxqL5jiDtfkTC7Ki/ieRspyhodLqBLvZdKr1JD1PrqxVGq5NMo40WKcsZhA7LLELT6vjwUWXC
dDflGn6Ve4Qdmuu0k1ydeO970HGk7MDdM70jWATNcirnFuSwy46Cm5az80FJO35beH0rbpD3FWOk
XuDsUmiZV3cqVO+5F+bX8MxPyksnU971ndowuI7uBVP72DVGgrtJExRCrxQ0L6ujbqIIbrVRGL3d
gkiH6MPMl+hVjbfAExGdfwFv4meK40J9xSvBQjEbMnHcxAnxvdcS1lUk7ejiX239eGNS3r0Lj9Hq
V1Jjbu0EtwyCxy7h7yMrRcNhBj1MMTtxtDYriSSG2PSjfb77LAuA7snUQIThyibQMb90AfwUjEqi
fydsv2htloN4YjIs+E3DTohfSiqRZinuDCDinf1012BCtxrJCTuO3euF87dhK4Bey5+jGAWoM2tF
qGcadX623AZkSf4K+OnI4XBPNFJ0VLO4KUtdaWeTtjh4oqJr0fgV9XVKubSsX7fssrbmNg+yBWK3
GN5QaBk8E+5QcUOA/aRsvD4KdwXjA9itFbGvrmRIu+uSNo+1ruhgh+F2JoSp/D/dVIwd6QAmKcnl
y1lmLpG2fgWp8iTZJCM581rb8tW/yfv/+Tj9JpgVZTt2j/ANvbjshukC3yYRYpNhE8oAruxZKEsV
THgTNbhUh3VuwOy98Msa5sWpjb0sSLLEKeGfDLTaobhYtitVow6YxwDkOXxlGWbkqmpDKnKEcHhn
wEThEymOfcCrDzoaegVrgJQRPfH6OkzrSLn+74k585Num2la3m80Vrz1cOSMzm24/ZhrzzJaguZ5
sdo4uE7IQC+ckZmcFEs7rL8LKorXl6XMdnv4cGjLHYWZiB5fbvZrrcu1E2EeNyWXlb/8lTyhNOt0
Xx+5AeKSna3G11GxGn0ORTGP8gOCYOXRA/3wCTt6JGY2SPZYexe70ZXOZbyvhgAcGBCrVBYGkAD+
yYcWGUCq984AfyG1af+sXDcqjAF4FMqx9b25OHudYKjShDjWWrxbNPnSMVWtdgoBK7UncoHidC1T
TMFCoI4ZHMoV+x4PMkYJ/MAwp315Y+ZQ+nnjTcfdc11GjFi1btnxbemge/TGpqTsrGUZekfTH83Z
a2XIbIMcLvUuXO/HsL2Gk+CEhdYGeQ929if18+tsLG0vxB/U4hKZdNkKr/RYeDF3qNR1Jx19YWch
ZM9fR+be28vqGR+rakDIxeVP5XE1UJa431xyXZI/0tvQzQqm0OvI5unPrnHI7+tddAOX3CMNNXnl
I6QhbnXt40tWczh3LSatRaLShqBeQa+jJuu4SyV37diaxai+JSAAmmfLZysnYhpuJdD+VqDgV2X/
Eus2rDYnHgFufUrtkgEi22i0vQDUZvombp6/E4AbF1EdjkXnvRio5oiZEHHRtda1tBjQuRraQzDA
JehgH8+Vrx2Pm6O+pC3Jsxe1dW18b2GAagDXGqzv3tA3wqyMPufq+uqmYTcftTlEpsFzhFBhNKu0
zNEE4/eOn43AaVSEO9XPZfdzomCaBiOPo3gyZQJeGEYrlkGezMPrMSDO2EtWtane0Ce5cK4RDIsM
g5rYaPlVzgKzvOt6Q/OE0VTcjRphLO6cBs7u9ND+hRxoyzrwNkLIsonTEdzVYMJG1VtubJLeRpmC
KOT7EPLT23wG21xZEFrMIOM6k46w6MgocvfWb5tbfQ0k3K12ObyPfsi0BAA8IjCb0dsMCG7rIpw2
xSme4WDO5EE4cC7GyAYfptNrt3pucmARlsM5DdwDk7jb2tET76nsGx/S5YAGCzCCg/kn0AEogT4j
fSFntQjYHioYGV41UCiM0R+X4b1D8fIcgY1HKDj/nrZWXOleLC+eR5gX4pdhLDygmTm9o0VPa1tL
B3hNg/q4JXZhw8YeZvZppc/vQmpSq7U6HIGuh1wjUreslkkqW6ngSro7xd+c/++h62mFDSOftOHH
0A/cX8fcSo4PTQQZeeDv1iAfyQwjRW4G0UIGxAV9d6luy6vAAR2B5DUSrQhwct9YpCUngUJiIvH5
U5tBVV0iw+xatOvZZIrCID87b+XGiW7hKyKi1nRRdeykYb3QmA1UK47S1w6UasP34x2Wl+4yviXP
g6sR//mqunZBScN8hlXSpswglqQtN6VnTpT6Gz8WTb3dxMm2vSRSD7zi1UnaWxDOjRvd+ZRj0GbU
y450xTYRfiEC0MpT/vNof5ku6mPyHe1q/2hp+DEH7RFebFnSCnA2J2MadnWtb3Zf1ggABb5u1N5J
5yWUGI+/45ZJFzG9AXfc2m30JW1F2OyuyKnkE/Vq1PtCTeHZw1PZllXtSyLm/h/YKN6ADodFB4wV
zy1QB7yFAoyID1yOTyRSfSRbHdGwT9dm3vYDx05PFd7Lr8nxCEa/piiBcF9xVEnTdKMrPzaG+LZs
c25lcaC894OZdMZ6+ivicBUlahF/vtF6IFjB8VTVyT0f3ZNQnNPEq9QEJ3Cc9uEDYd4pvwET06/b
+f4ehWUrV4CF7QH6rh53FBiMfrXekOjvTsZ32DdvxU9l+WI+jXzMS2nuwqfpFS+NL3ToAA2VAiwO
vovk/U+5mEdT2fbB/uusVOK3u1VBCky8Et2LL6UFH6HfXVavOM5JlKtew1oxXsuuIiEs80i4KTS1
sXwoqLcFUwjNr/yVtLpuLTR7Bo704F6HtiKXvDRZV4TvSj6pqxqhqhTwuS714YiJ5H+d2Wt6uQxs
6+0N+WKvSBDLVesW8LB2tT/ItyxM/nufZ98NQ9yVp7aMp/sj5UZNO1HIIKGv7xzHwaQB0r7aEFa3
tOH9VeU55njTvlQtRz+rnpKO4txqTyQerO1TGJZIA6smf/V5b0q0z3bVchVGBjyy79vBM3PIldIZ
WVlJMrrfU4YHJIf/GP75RkSVq0oeWWmFnHc+efBCI+KHGPnmK7WgyrVaFgw+r8Ta7fz2PuJd3Bsi
zQ+y86Cwepp/DKVFMkT32mtzyuLqTkTYfxk64Utv7jCcIEWhelRoO8MnQq6TWQpVpOcShFywROqZ
yKPodop49cKrMsRlHVy/pnCd26FZKRmvyWvaGKPFf0jXxO6gd+u4z6v5/x+1gj8ZXV3pVaN2ey+9
MDoxzPsRAeKbo+H3CnsUwxTepSo38po3OqviwBvG7zuyIIxomVesyAuimfhtS7zhKDgOVtnKQE6E
IV5d+TM337QHEznPJZqUimike2rIZwI85Vc2dGBYQxU4Yl83K1JPpo+7/6Ir/4GnvueVSK/JOSmW
n9p7IgEHtQbWEBAUz8HXgOqm1um1qM4JcyNz/c/ynRVoG59rtuVeVfnf8NfFBiydrgwb1uwH1w2a
wMfppkKmczZYka1p3BlDrXZsFwjK74IUc6ROgk+rmTdk4Dd0FBgWUw2LdkBqmA+qqgEIxxFttR7z
zsEag3vDY6F0xiLGfiQourbj4q17tY1VgpcNk6iWSdV+k22asWKhZ8ZnDNKlK7VNz1rsWrONuPdu
v8xFUSMZuTEbqconwynzoPEnjzKymc9PkSuT8vhc88rNtH+/8iv1VQfnEPfbbsjs9vOJgbMQVdBi
RDunAX3URukr2hdX/CIMnpuyyaQQrjvKDKrNUeQGK6cY+qZBY8jk9TDKOUcIRLBXpUmGaqwqO1AW
Y3kH31N3uke43NRnk9n5OqkJlCk/zRxcejYZCM690yqA1laMcQ0ohDkHBKDWocwuurRVKnW9YDLP
P9fEsRaB7FBTT9Stz9o8gge+ST/5MpfpHRX5I+Ac8Oq0pudghMrSj0v0M4petBcQWDehmBFdweUM
Njabi5qVQ8OwPcAAldzULIocn/QNo06izrbdc1gZEUK7X+7GsBb5yzRmvN6aFEF8ZDf9oVUDj2b4
z7PnXseLALfgKHW8bnnepE+yQbQL+feFJfzHbW2iA11szEbjCz5E8IjgBlWWG6/mwuuwsJfX9MDr
cyf+T79N7bzlCUjDLH22fPfgZwpx0jjZruXg+2y2pjTFLTAwJbzwNxVwAokL6D8xyMr6CZbqxgfm
aFHVrS0FeQoi8F9/F19cdfZemme5i1PxOlvlCv1Hs7reDDFctIdtrwO1jPV8HYntRfd67QxwTsXM
5VBzNKKgNQJJ9LXKDLlg4HEpyWk44mbQI6oKgk8p9ewZesJzi+I8Hd+hW+Hl8insxNLR5yOS/skA
6ea3KNuqb9mv+YYPzB6VksXOXY48LSav/RZ7EH6oCvl0U6cYqUgKOfSb+AdoDYERHiE143XLrp1F
dXvlEDSQkOzxnayLDEIXFMNcU+fUifsPQvg4pWCvoRuy9IhtEOq7BnL5FHSm+dzBZoWwJBioBqvW
WUFIzDva7jbypIk+RzDSQhPFAqzn2jN/oxy4JUSKiCdocPBDUZC7b2f4a/AVcd78lyhPCs1MBOcJ
lqFKDFyfDOQ2I+8DY7uwdPSn4RHvef4j49UCp8+7PJDwYwhEBuF/AYkO46qmKLxJQazgzMpiXuW3
wTzySrQFTKgLjbJ6EUiGnw07QYrrMzsib9JvdmjsD8s/KhOHOzdz9G4t9xulfSzX/cdIfgy81QgA
qTr47RcXtNC3x2bqMNN1iF042385LzW8xl3w3CCK8hLScZuYPoe3yNxBa5KixT6bNoJQj5koOZDJ
eQCL+r4CT3TqLNGwEq6vl+JMuJGlKppnReGOhvovU+N0c+1HJI24V7CGBhuaiCfZVKLKrJPSAKuG
X3ybbWZaY5zbesZc8eY/LmZ8yAbrGp7lAjbrEDcU3J5CuEnpT7a359WIpt9vctWUjVpfBuHyWBur
+cEoScV1ReoLxssZ+sSfc246Hrhzu40bzOAN75hLMUBmqMiyBDyRHob7jWDfA4TgIBShg7WkOwLB
SUHsGquE4Ll1+O2l0moKdQmh9AiyWe/wXAztTH1jmSQoZpMYS7kWOYqN8/1Rp/lsCh6ute/6Gqyz
j783+W1AXNGI34bVzKRPoh/wkRRp80I+3IfFLZnBY7EXTbJwrBPfnWvkYFhtTxHT3oKOnDtXJmyp
C/MYBScooXGRlkocauraZ4yVSTF5SRZLP7kGxymAKdIH8J+e/KwESQ9o0pqXdrXAPhoYnCUz3LsY
Qjq/IIGuRzF/AXV2M1r8/6d2sx14QtwOym/md5LJf+jJUcFwv6WAMmzqEmTiJTiWAlFOHZy1Denv
WOW6lE2DQ0aBOthqHDEtt6rjuroHS52prA796B5g0Nd1nP4AsQ50F124X3mNyn0bcddd98AFjiX3
4XV/4MQi7aWcKfvLKuuqU6b1/f573mrhaP5O4fOg3vPNRGX0bsEjurbTS79hVTcm9bnFeZD696lu
3/rT1vgHTP4yTYA0MCtPFGARwKo/unlIlq4mKz31DVY1SXB/TNLtfha0d8NbaqyMBPkRmEFk7qhk
uVXilGzQvH+7lc1wfmkfHv0/MlJSIdzslPcT8ipwCPdYnVf6PGx3xIAtPT6IOjk+JPg0r2+H5x79
oaUfV0J+s4PE+91/qtL35oXNspMX9oufhFUXfaKBU9wptNpXrOFcNlGPwgkPUkVDdE1rBPvUIh2d
SK6mw+KU86kI2oJxNVWKSxXFEzhkysAkrozFnjfs2ZW69hnd4vuc57xzPaoAWZN/L9uNjz1R64rK
wSDrU/uLRTh2exzPRgZs6uItg4frLJlBHLgUnwF9WkbORvXGMrREPwUlqm/GOQ4JxjyS7ufdPsIE
J1FVyWV9nLmBIHr36pOc+F1NlFFNyeNE5ONDs6OwMu12gEdVe0sb5KwGy8kfAm0UjDlfFy1paIrJ
tAM0p1czJc4XihMCXQOTM44vP8KguPnj2a99kxBokuZ48KWkOA23vc0VSHqR30fi7Xl4DePevFMh
Kc8yudfMbLQsJcDVk5570bqI6D+tL/5tdfYAi+2HhqAZRiWYE3fI/+qJWMRgAtljhj97kb5BAOkt
9jPViq+6WABERRKe+xnRPl+TZVypcEAuMdSUiyrosdnyfC4h8wbDmzWZi7AyzB7Kl6CopvC8qF66
w0ElySLbGlonqlOTDZNbYbzZXTcuoehrwo0X4dV3JfklyVXZ4dPpwVjS3j50cK9ejq1NxREbFsEU
NwA/v4dUhhhEnieHzu5wwJ9g54XvC+W2CrGBJDQwas9eqo6JshhsMziU3mz/OXSDujO9ayPfDwTS
Ah3wDybAY1tdhqzwpr9zZQBP5On/F6MDwsNgjXCaRRMcNwolj7GRWxIpukAZRIw7tP9BJWAbdvQK
HJEV3djKFpcjXzwrSPhIL2FdisKu4EaG7+Jc1YPuMgoaKci8aFgwKPpNAM+/v8f4ni9nSSyDkMhT
ktO9yliIFQYsymvk7pgaFdDRxWAZpqA3XLGEjPSyUEG4ZyLxxLbSl7C3DOdG4xsZ0dTUYJCwjVc3
r74IuBfBFhx3sEmkMj/zx5xPRdsdw993lfuT59cggdX2zNqr9g59O59SmKS4PZ3yRCyJUoUj3trR
Udbu2MYTZMFwl3IhQ67Qz7JG7VwzW7sX03Y+ZADN0ElVTPbqP8KheRRfJZ9uyMkDDJrGH4WSjXQT
HaEj/UrDes+W8BIiVnMu07g6E6WQF8wP3/8KHWtWKMMmJLstv1pgA85v6EunkyAHUP7IHR0iia8A
BgEbTEtYVy73FJjr4RJDS1aUsVv7WlpEiN9kgmHH4kLbsSr+qouATru3OnOjc+Jmh0Xab5Bj0gU3
r7zi5NwuXWF1lXzGpDjUYwn+mFosWDo/eJZtZjscVgVDAbod4Wt/8itfajnzuOVIrfKshpO3GPwe
PWU+2ytSuYRU5MfVc/6todB2JTjviVFdr1zD39GFskwsZYXe5toTuKKksFaI3kx4nHxW5Fci+iQv
zN3GHWDqAEU3LyRj/Br8SmO/SzsrZqFGPTvPFjGE4NxoMnomhdyw3NX5+Gyk/KWIaaI1Bozl9G8J
yzNN6pSM5ykSeL9Dg2ZbRGnqCFPP8kme3+Gdr7WtMdbIiTwl1tg5MnS8Qg74N8+JyS6XyV0cvEWE
vqzc1rZslJOGlHj0pASJGil+iK3IMc83aarUdnnX0L173vxKScr66muUzPkOQ0VfjST21rEzI1sz
y5FAf99CJxk8YT/1mOkAcr44ocBjGC/D11wCjpX7Jiy7AAbjb0DFnaa+4KmU/wkbK3ubGf1ATDod
hxLeUfdLiPlE0gpHrywWXsUbK9hK4GSVzocl6XlcmdX02iy669EJ4bvkELGdM+0Mcl2PeZMzoHMp
m1M6KjkIfxYW2AqZ/BCL+UuTY/Cth206u3l3U+bhhL3zCSGzuBWp0PBOzbI8ApdeeVxOThUew4eZ
m8CiN5It/R0L/d1R8DY9A/0zslGuszo9GS5mdMtSKyHg6xVUKV/RoPRbnk+/GE9SzpBqD8KCbxCO
EUVTX+24GsI9xwuJToch9mdTjnoBJVT+AexY2n+8wpgj991zkoruk21dE4jaUfS1poEBzfuR4owd
ZhPzQ8KubVt274QnNj0sBVs2jJRSKLDl5hMxYXAYCedzeXtAijnmuvNtG3x01O/0i8ij2Qzwev0w
yL/cHR2SAzzejIJwNU/J0StiPvCnQKfTlrlwnPKJSjhHP6ZoE0KV+mnEinfa1QRkZN+Ss8h+XaUb
0nN03dEIjjTuzo+AHFvf7UZ6JhaixidMlwpN5iRAcQhLz5KSTs/I7ucysVSzqnLRgX25ddpp83AK
9PtkjfnsBZqK9VN4qluplAfA4ddA8vcIKKp3KUicnPLacSaz2yCpf0VtzHA8bPxEt/TVKQBubkNt
2rKMaTi1AaLkV7TyXhsPqHX71lgetgi1pF6s5eDv2IPXNwx/nmHnOrw6VPDKOqdAP3UIAZhY9lAt
lA/2IBXkToPT46J9yj9g+J0k4httoGaNg8pdwDnCxiikTMJO8aEm1BLwNXxDfjViq1FEFo+SOy35
+OL00Dha+C/DyJuZOEWeqNGc3yXj9rJVo2q7ZZC1rVrr6IBvMWVQgHBYPBxcz9RV9yG8yx0d0lO0
5Q5WEUzcOoplAW4jctenWTXvQny6qliNpcyRLsmWKN18VEFS1DhS3wSX99Hd9R+20oaJNfplOYCu
0AJIJWCL0e7yIJTiOSVF9Zvk4Ji3Qk0xANFC6Ul+w+MFoIIlF2D7xg46YnnCsqPHbsikYUM7HGat
5jTz4bnPy3lKE9Tb41ya0TBZpDeZUPO+k0jaee6Wl5sIX+/Zl++MhLIG7Yxt2casOTN+Z/yoJImQ
gVcRpgNDrOkfSa28xyA2Tg1mEbMKwD+LEhPA9d8xHEAM4NgCOeWtD88m852m6mgP2l4eMoAeNwHs
sbU8d5bH0TZu9y2EYsVYI2vXZcXdmPqyuvty/n0KWmY4sd3BelWBZJfLcZzJ6SOqkIDCk1w6B/E/
EdsNcFg+ZiOAWM4yeCUdOOSJRZAQzxsRNoyENrKB4iar3hygwZxprO8m+ffbeV24+bjJ81M3lCfq
yo8XlbklnlNkU0AMZMjMO7mrVfmISMMqKm9v2n5BxQk2ADY/TL7VgbJcH8iXYqMP8v861aZsuf7W
SBojeD97Qyt/O1u9Msl09dAO3vrksiGfcfRtCFNW8YC/dEuG9dfYbxHlKplz3S2zeVxJ/vb4FmfY
8ZETUip9C2E5GrtAZHgzTgnmT2fm8aikXu96HdQL3B33Pm++PNBBHKRDNKyygmOl8ZvDV/Ss/ty4
zQuPf+P/JsFOVzDlaBeCFPp76i5OJ8vKYY2vDnPOPYlUpJvM2pATjq+Fxa88gWGFvoL19Lo+r91q
p6/vPEv70PrTCsoG7QOeAwySA02sJiTVPlppIugzlIMjK2m76g0vwyeL5JIIb3H9FlRuMf+Vdtvz
txduaGU/W4Hplo3ALYPbmcyPC4ln/ZZMAElJHO5BOVkjdS94a6zRBh0KiUozWfVcVVZqd/OBijpP
A25mqz1nJRDVe06l0yJcBleSxp44KXw8k+ilh8vLQBvaI+GrpNxT5Lj+32p3NOvGTEhXeBh4hj66
crcJGhwFRfuWiA9BYw+c0xhInW0Y51zRstb2Rq8rPgmqTbJ4XZgEvMsfrrDeaN73wTHSjmnfW8i1
tHyUw1dnS+03oa2bgzIFVnT2lKgJCzDJpXpHgVimk2OdkXJHCxrHurQT5hnr9JgV7Rj45PSXInML
MGUWW624Xi8ZpE/Cr21ZZOBLgb42my3xlP5eM+H8CmmF3MrluF45hMGjpTTpBx/I/MtzGwhQBpll
7JFPPJ/0QTZwMqyCYN/CnH/A1mmqGk1DbwaluqRNarqT2l//mBjBJ2e4HJVVqQ4lKi2tG1jCAySz
5C8Qp7Zgyxsd6xf6L4mR1lUwIBB0XJXYJ5YiyFS560C/9oFCH2DLsfa1GhqB1ONoQARZm0S9JZwA
YJl0+8v2Pl4VSwHbtG4abF2UQNe+S1OdXM8MAF4D7r3QtW0nAT9VT2FiAyOsCaSdjBvMU9/0jGVM
wy/PjIYaOe3wRwq29Dh3MrX+2vuJ53L4TTfVA197y57AiIXs58quhBUkzBfiiq+/I9tSJY5MhZ3A
Tzp9Ot53Eix1ZRMrIiMxoAMiyHAF1J/PO7I9KcB/ZGBWdDifSIUhqerG0VKhmTjH7YhQAkEl3ajR
jDdwjqkVWQz6XyfaaKvn7HsVRO1VQcOubRp1b9lbj1NXzwPHY4B9o+63bSrTDtLAPpBP/65K1WRl
yrrCvlSKNgrSYmZmm7d/1oi6sxoN7vvn9NwuIl1Le2q4gHYU/NXZG27nm5lWRkV7kd36ycP+gVio
mQPd0AeUG6fApSJoZHJS1HhZs0kvVfa5bsfWXCWSirGzvGeEJeJ8ySWjyS12uagOh6FYKS0YNwww
WvoqvyXeiUoTLpJSSyE9XCcobB3/forTBirOcqfvC0jFHMYh8FVDtI+J+hNSPxP6ejRJYoxngSM0
lq8aOna3IjDjNzlUquyZ7cKnsyszJAx74klNDxd4YahXbvbomdSr12hiAwffL9rTEA70q44Z7te7
9EyEFF2hQl8BmXa0UgJr3GLGxldRFWQnBdaGW8u6m4C+YP3wtsmgXfHuCUHwRFYq9odZmj08O430
EpWORfJTQwWb995H4UY1pS7G6MB7cwe1Xu31RXRWDfhqQBJw2xxBFvaVgrjHT8+CmVWOddWt8hQY
SToCMw/sAXSnJ9KhM4XPJ/mnj/hRSBHvknShNLpYlxLLBCiDGMHHAWCi2eBoRfgf91EbGeWC8qLa
jMqCG1iUl6iOeS91bgeWsqsbUMcxis+QK7hQM+lysMwGFdLJj4/tI7Om+6kmeGRpGR9ej/UNFkV4
08jN4Dy/QoMdv+5BXOxYrlFtSjugydvPt96Wo3U+4B4bxkoYKus9b3hg0b0TWIVXruZuHFb22sz9
3rkuUYOnRE96i+XN/uoWskQlwYWRskfDaEAdWyCWspEZ00dVlT1EO4DZPg6zBP6eaBNetfo2APiQ
Vg8lAyeJjFb8dvwL2M5hoOGwS34xcmUHoo690mLeniEeaOVX6YWv9DRFsOiHT/Jm4jbL8G0aTry+
uFYj9A/ZictOjhqylCq2bGEiRzQYOAq+VW2O7QPw14ruyrT6PH9gD9mY4Jj9SX4rYELIIu3nRMFK
Oo5ekjF5Oh3R6X+ROZ0oGAxsYlXa1qHk8mG0Ux1feArpjLlKlJU52xpEQyUQOm43avVOAVRDkYvd
n+jrr/V5QaR/W7XPZdV1OB4nVVB3Eyg+cd/NIB5VMBpwBvB37u/VvlmDGykDtn2SOWUFg5f6NLcq
hXMnr6zW4uZl7eyYqu6EWettZM4mES0zXNeUA2Ub2CFovBOH82A8gpjvAP/dUfM3m5j2nHRTSWGI
/oCSWsJ5yGJBnwZQT0sBsSsU3gqF1iLuSSwq8R1XaOc1g8WVr5oQjgLO8YLZIymzgI38gDKPTGGd
gFAWvKqCnaVb7bxMx3vgOwJmLAHs2+WOKiJFYaT+0QZCgAxYN7CyyvIgOkWJe44KppaeZwUMlhZj
jo4GkafOUOIGCMOfXGMPu8AaJQ3qB+Cb/fi1FilEwy13DqCkIAtfz/YUqH1m4sp6dpOOcm7UhrBs
v7RGk+2+9QU2t8TYn1AdUAOi8nz52hSOE8ZfGjWwtvajYQ71kYNggZq+H06J3KN9em5vz8j+GWXr
/Q7t/9WNKVPI9v+UymAdszYjTlW8RqlVU9RyM+h5s5vh6P4c1rBVTfdRVYo05HYer60SOHirg2r2
8Vym2pehKyAGiFreNfhEHrNSd/YHBiLSJyIugZAQT61ViHArdJpVQXSA3UL6qfU4tnXjSqFgOi6Y
53NB/y7QUQ9oK+JMs5N+GksHlyBY5eaQB4AsMbvI2Zi31VoZhKAEUAmqR9yfL4bekO/8BYfFwN4D
+FDSXOipf+sb50eCm/Kp8B/7myooH8eT2vRAAoVB6X38vEwbYJPqN9xmPf6XyGQjFlqTE2lu1RPK
55EwyMSm1H3OFkd5dL7AuoHFixokAfZSwTrOI55QAycHBEZyRLX03q038ePLfRFmbFh0Qenlb+tU
yHuf644NyhOcZhG4kqtZhEqIInHCPvFvqUGNZ/FG9EDp/Rwbh8jW0b/n3KzsF5oOdDWUk2zlibVW
RE2gICpOvZnpc3xym2X2Z1KW5kqW3PjFXKj0T4b3GZ0AKL7vXwwg4LucJN/dRPv6OmP9t4z48JqD
UU8AaG8waJtzQ0/44RQ2QIyLs4qWToVzoNS1jv3z1ROjBiOYlWzDtwidegQcGTMdD14tfmaAWC8v
rs5EWj6/PTrOpin3aBrvEaJ8Xu9dcQM8uG4Xz9lt+7cWBspbe5Ukc96L8xw8p6zpgksnhSvyk0Xb
B0YFpGT7p7GvwYjDYLOOrJ2+7qMqTaS/K4lA9r7Olqr4hWWovorP3WEpeM+JedfxBdLT5wWl6Wrm
6QLyusNy1G10rqmMSGIACnRjwU0zQVL9B10YjOrziEHXQdqPFgG0cedGpx4bJFulx1ElOR73dB89
7j76B13Evhbyn2iRLbgA5NrcNBX6RmOG81PWc5x1a5H9ukdtS5MNf/XA2uYe2ocynuwXne6fwbIv
IDpgVqXRqZK+1a7CuNkgYNNXql9WRXdfY+6w657eGORrwI4xj0mKFTmctHUVROm0qWkRTmmfgxik
L9hEQtVXZs3oozk05L/+lmR2cygemuOUb2S1AcStdEgc4bFaDsORzmb0anRj1ujrX4bfGMSPYjpW
i6aqESRSraXWWtYuaIncEIGIIPp97/41YJvmva87DUVXt5HBk5AsC6wL+e9zZiivwKbix4y/r9iB
2EmL1poRlAR2LxmRli5CyEWMvm7Md0iOEgLoMMwwxGUgTf9Zzucfh3gLGWBuo3kBhDs3vEqp5wsE
ethBjMMPrlUen40YPOVkPiDYYBjSZIU3/3PJemMonrj+nNPRf2gdGP0SWLjoM8D81OhR/SDgFYcA
p+7GOzfGi2lX89kaC3kAnfQQG0TpOjPBAsNoiDw4XCdjsC9qthg3Hx2D2a2CW7SxGMVXPjY7++tV
a2AF77zwc7iGM59VApEK27H+lDhdtarzrvSrRbUkyKm5TjDia/cigAL9yrStWos2EthaPBLKckxG
fV91WQpf2rRYZGZb0pXFazFHkNA3eeJOYhjyqLpKIogGobWBPzrLFNfbiNZtIueWJBXHmyVBSkk2
+5ikJaXwv4dv8SxzOXkh0Xf/CfXwLnkQlDwwCcHbsSs1iyB8/ZlODFFDTR54B7BRaCLfk2kPnfWO
CBWJ1cqcjlZeIkYd9+iTlFqz5UDgeysWkM/NXv/lhuYVc864yNhf5iwUlF7oMfHORtsBRhEmpIdO
3CZqrxfacGcQqcHJWPhhtgNjj7lFrVH1/dC5Z4+swUIn4oFcXOU/U4EJrECp9/4BoqNrDIFf9F5A
Tov5p6BsxBaZsT+f2KHrFd8EE+z00trrsKLzSHEYPbAaxMPBCH+MmLossZhRBTAmGiJg2elqb4Z4
Xat+nG+Ohq5yPusUljfIsz4LTsLhny8Oa7PQ6i/XW6p2e5o5/PEQd47mEGbGSYqdMLZykqb8Cdm7
PTQoeUmJYF0m8KRCVcVEtEcMWVj4jWCBSTFa/tJGRqjg+MP74O9DM3dbAQ2QcTJHJV2r+G2a+dAa
hqWy9WiTKTnLfR1EsiGdGTG+QZC5MEuK6Df5QPvwHdVguSYBhMMBYM7bxYTzIPV9BpOSG5x3UDrh
Xi4F02hb/KGSagb5MQOH64hCQK62JISc//20w1o2AmESURbkZmFzqos5mdwCPaO62mJEov6TdSKq
97e1QRUqqUFbyTD98ThUe2be6SwbTVJEFc0TAMA18aThBiSpjRstKM75F/lFEylI5x1RWicZzrtD
lwCMfRO1Q0VI2PTzu7hj8oYJhBuED94bggq3uwGLuP3awayAplV0wJZaZG3+G4s06aTfj5eNUeN7
+a6OX/tQmZLPuTsfSOpM5L68ON9AIFsU3LLQJVxI1rZw11skgJR5hPWzoDV6ln4fnDAfZiix9Z3f
xHqhWxRuF0YDBjXCcp/7Kx0aEtO/pca3GuGWhlDMo6if7helY4/P+gt6AFAadi5q+W58/vChq/c3
LmNqRtAfmAlzxlcqGmwZPujKhdGh2RuAwpANP/EliRT9fxREF3Y3nWWEwbNCMse8BI7O+tYbsIFn
x9DUsyd4mgtTL2y1VkLFqv0EuM8pykrz9niJSSCz/uCam0AGvkZLLn7+CvKDfsBWqpNlc+3D7zE4
hspX+OT/2D1FnpFNnyqN/Iz68BhdR9k8faGMsyp5GjXosiTdZjZllns92SL97Ixdp/yxXyeQjQk2
Gj7rORBhPMgGyOGPNtZf20UMt2XIg4mYwtVz1NWV//AgKYKtv90g8nsGMeeRSXO4GOYHRyh2zpx8
r+WBoxXqOT1XA24XrBDbkM8qRKTJSa6uMtNiZFdzXMkJddDBNVKA8fOO9RXvRSRi6wqK+nYmaRtA
R0eNLQZZHm001+Vi/tN+XZQFGqtYexmUb9SJpGB3veqew+V/Csna65d17TB9qkKGq2y/sIuS8Hnk
fgjpWXxDFc5Qs6CfBcEK8t7ovkfp8kR+FtZiK/RIcYsZtONi2uD31zNUuMXex2tGmUCencAdenjP
5xaYE2eMS/N08AKlSs5qoFJ58GW+8a8t8NCRy7AB5CURP3DDGwwmfoCiFL0awKFk0FlVVWtAkdpi
C6/vMEka7TAvI9w4jc1GUP+aVDMhWIWckU2B6Wd1QV+c6YWMp0PLFL8Sp7HvsceXn3E7P5EwfZsb
WvxeRRys+SuFATt4IlPGkh5P3AI8Mx7n+TUcDpd0AKk+E8Awl2iie6ihYs1fhUZz4j75wUwyLjMd
ESPu79T87gUvQ/B0BJWoEzT+u7FAiE8OfQj12W1NOJ7ALuEdDD7Jx3tA+cMnNojyZd9/hVmVtRgT
0UuNaxrQWytiQxLnsiFtPlb48xyLsoykIFEgXZpmXblVSeZ+BoR8+JC++0nxZQaIoIo4UhVxXzWk
TtZ5pK74CIjs48vo7x7FvApT3lF/rR7uqw8l5LgHscwOsAJE5ygVgv1ZB+oJ5gejJmiUtViAtbsr
qBYM2tmYlZ1/DJvdxzdikY/34ht+asvGDBmneZN7eRI4b/fxE/JUY+WgyKH5hpBTbueKhOkpBRVQ
aZsxIXFZTUXDXqN6CihRYgBC1ZHn38cSzYo4wcnc7L1lDv+Xn6d/qJjN2dph2DHw0rOqt39BYptQ
Sg27IDsCLRruiDjUl4Wn8n/HI09Vs3brwIypb5kIom9X/x1cUqmtxmLQpe8MOdIdxnPkQ3JzhogF
3PG80RAttLRRenlUzOfYuqVbtAYlJzGcJYfG3tNmOAhHpN1Rz7lUie79ZeF7YDCnQwNoWycpoxsV
RnDGBPmEAJw3Ft+hiNOQwWecSeMEeY0ynfOCVWbWNfDjOzd29E2bhxXn9uiTn8Tk8tNGbDeFeFOa
9szkXY1x0fJeN2Z7CUpfthG0A7TgNn6wtuILjOMavafCCXW768rI2HMy3qqN9nn07OwuzGMaeqvQ
iZ9tb9yyaahYqdSKd3joV8i/++Dy+IeOsYYhFm6BqvvuZX6AkS2fD5h+FHgEGv+/uoGHkgUIxvq0
5BQso/PsIOBARERNvKzYMW7g2z0Pr0CTFSq3odUBbun4GoFphpAw5tpxzJThpn9ibgfctyisRfSC
cE0fQoDWkW4/1GQag4JudLxGuHeugah1HO+uqHfpFV2VeBlSwtnLcUJFNdvUHKx42qQ3DEKs3OX5
sMLjgw3fiifJtLwMs2Xyy+t0r/2RqI6n6VGdhpW28R9HtyxNaKk9/9pvSHX7T8AF4WSFzm9FeVBY
HTgSsQXUMEdQNdsXw5kSgwo6JBGCS3SleKOfAuHtjtE2muUKHFlz+O2evKUuUKkHybLmuqpGlbX8
u7crcRVxPrPdYOKYDE3F1fNf2IOZg5RdnAOvdAcDdLGTVry2kCR8YwyNjUyvzEoG3PfX5DR0WGuz
xJJMrLocoySXlfR8O4f/qgYK5Uu1FCYMD4eOqOJMAw0qdEkLoVE1B13oNXKd0Nk1YDLkht9k6tvF
yPHwn2Ej7bxegGEaYdTRO7kjdPP0SbZUXtxiqfZpLDbBI4xokz5ARu1Nk8u07e+tWET+1+UF9OUr
VoImj6G4fTQfsmk4OsJ2GlHMzvvcmafy/u9u2cels7E/W7uJxYIeLADNU7YfCRPlopz2dxxe8eZS
RfuYAuzM9xLnr3rVuZiBYzpN7KbQFqlJ38X3+K0iSj/JCZ+wVPFN5heJfQFrzKWCvnvT7utYcLL8
xULITdoFBA8GNXOq9jIwIN9lFMU4VpqCULZ0oOqRCoNXrwpIN3EqSmG+HPaQ/tJpVOmBIX+DfOnW
JnpQO+otrP9ImdYK401Jy4IpTxxD4yLF0EaescxXWktpXM/0SLbQBZO3IwUs7ZhwvpS6KHEzaBsB
oCZLshvjNdMHG+/MfKaJ511FvAYU6ngKeVI6OvT7qAiP9gb/TNumtP7Q4uDYl0Z+zhfqdmbPF+MI
nvBmsLXYJITS7XDuwHQoKHi34r8cCH7FE6TTFCmv8tWm3oHs9sIAGYgWCcZS2OFxlNufv1pp8u6B
vzBY9ECfXBhVJ9px6Gm4XQzuGbfN9f4tydIDronVyoZ0c78NdT11R7gV0RBXo1J5VvgXVdvnXA1N
D0zvaLQSKcskVctbKANXGq2Gi8i4k4CycW3T4O64U1CweIVp+gIRm6FdDE/vQyl1O3n0+t/PnH4D
+XlxZ0soK1gc/5vQhDbXiWBw52u4LY9Hp4+WVlkjGCNr6LYVnJqKrJzKxsOON4ljQiA40qCSZfE1
cx8mBjQsgN0+W9OEAgRKWrnlTr6L07CWCxtuZ9kHn7X4HAH7gtEFFWbyDPbRXev4NVIBmE2HMQ+f
nYqx9T7QIdt7mRquV6agqBjb2EC5veYSn/VsJpUqW7NKcxRrb4K0VLN7ZMVGXoqtIVaLxvKT4e0S
D5tEnYU4W/rWWXMpOAC9UL+685l17xN57VNoE+h/8y+zoqmwqEQyjpNl0irjz073YAb7KKBYQZKV
NWOqdNu9s90xSWBmVGnz+FKsz+3rGFoU0NfGhv2Zk9QDpcInrLaKzyOUAWUHqZiF/JXdbA36MsWg
77aDL5/NpraWkbe5FqI0KwuOeHBZrpO3JOp0iimLk/cL+Hmz9Ea3InaX8LYFPUiG9YuT08/ii4wt
A4yUQLfaGhiDZGyRsVZ9kOVyK7QUoIk4WgW/Npp0nDkLnU4KBFvr/r8JH/pJQt2QGHdjj4drGI/O
PdT8oqXNePQNez7Cl0seLyjk+KkyVQzMcOYwZwtian+wScZveZrLtLUH+/6riWpwEd5U4Ds2kEni
QygnGDC1B0hM8fKLnyk8heo+YO6bBlLOpVxY78LMW0UNoqHb2WijEkCd2DdKid/Omj2XhLqzoDD3
MC8n4GyVdM+ShTX7X4ICR7qbfHgd5YpnpyIxEO4YGI7U2ekoarfYUTYR7jOSKzlfN2j91rGIBeGZ
q4d33fQ7Rm2Vx8XsmIEuI8yto++Hj6QAzo+uJObfT/qCcZykoGJFsSUM3W/WKBvFhpPX5QLtxPok
D5e4Hi0EtRd6u/MCMGSHB6uIvJsZVJSOLk8XEf8E5IYWtS8+b3EICETNj7aguSlsI4GK7nB4TgXE
lSd3XF15QEQraJslCvewPk6qNWZ0+wFC6K5E2zsDCkaxSFyVwr404OUNZEwJzLiTeMfTg3RfoOzY
PwkGuAf8FvKdcfYuDXeLnXV7/LkPXCGHajOGVm0OYZBRv9kIkysTWniMPuWZbpCYsF2NngsUf7bI
g/uWvixXww5LhcD1SturEqv1NR/6OHfNvACwhOULIqtcSbBrhmqY9liAQMOC7BaG4qKverrVyfD9
GwAP6Dyhx+eGO2PxJoUwYRAwxB8b2y3YP5qoqBH/iQ39FqgUCm3i339HnxntQiw/cFPw723Rth5k
I7hpj8J+il8PmsO6xXhrnCb4cDUaUbFvgzzWnweGN+CCH9SeHwWNnuZrJsv/MzLEaKyXl2lYWVBt
bIpcTY08avkWDIGo40DmgADLM/4J4cij0Yhr4JYxhjY17j0JqXAv2hwSc7z2VdSUS2Nj4y96C2cK
qPFMzgsgaqkEbVG+PzKNbRn4rRj1ltyA8hn3O/o2aTGFJHpkz1jxcsICv68FFERTk9OPCeVN/dRr
FVHMRjHT33M3pri+81sluBw6FWC9kIJehUZb5bgyuqotIOwCM6FSoTA4sS4p5CX9zao8kntdOhxr
RRfSroOluYfsE3ALxX2MmyEiRhPuZ6cb5udybjnCZ4ZUSTFtbWwuxlHFgSQhM/Gn5YSmwZj1VMn8
u5XpbSE074JzoeIoIrrp7DB7f1OcAFAEybNk/Y6cyOQx8gpBhiGOlQxHF/SOU3OPx1UEoyErhE9D
tahSYPD8ucBJqu9ymCEv8qC6QbstR3v2lIzVcXiY1K5Xpb1q3THOkyDnRSRqvhGOmiSRvDI6slut
1I6mDopAS2QHWeSYmZgZP9uWu6SyltyiUEdfFA7rxve6PyPZVyX215fPLHp57px0ZPCAozGOnRy4
n2pwIs3Fa8Kx4y2bvl5wSv+4XXrAkSLZB9wHOo2D/o8EvIomluJKlbsQdV+s6g2YbHxbZ5RaXQiX
ScePQdoCn3PY8x0O1ITjGi/uzyNcmmevSn0rgGK8YSMwQHvgF98WdQNhl2h/iOPPx2GtHxe3F+Ui
XIakwW4PSoR0YZcTxxYc2C5pvyerrVa9Y1mRNgEBOmKtbAa/g6244d2+A8tsTdvaeStIGunGmOHV
VZFt0vAqkwshAMceIC9BYg3ZpCyp7xyIvAQ4xQpW91FRXs9z/Bn3K1UO0A482BBAGAj6cL9NkLpT
xIvm1omyzNSOcnJB8pbIFitX41x2xHAuFwuS3Aw43zttF3TeNOi1U4G7BfOYI0yQ4t8aVBl7NXhc
8ncNJR5YsyTWOBF+RFbTtRCjraUTTvpyfEj9eZ1epoj8VX915eUbVODcAJFm0bvX8EDeKhtEvSK7
gzOR/2q4gjH95Ws5E7zSyWU4vtcLiTC6heB8EInLjjjEXId7MbmVyJF4tyZ6zPrIfROKkBd6VR29
20EdQMQ7vHLnVV/gWypu9RGJhbDSbpWXI2A9+xoa76O+jfyHlr2TlkxAeB7588VVykmf6TOaKkFY
hK4FHupLSgkOJjLZXwAUWS9y5wqLNlxJhAW5VL9NkHqhUhmePdOQr8Yr1fyxqno//yC+BX+v5E/Z
nj7NfjPg12Nc2d5M+03qU5dO7lMwfg8EMx9Re6q33Gdy55m7xSU+FQPDhyKfm6Qf4r/K8M3is2d/
ng3qPdkoqXeI8qNL/B5N16Y2G48ufYlSZVM2nNgbBSKidm46yHlJ7IxKa9nL+E0GoM9xsDlNHOKZ
S6RrO3Aq1W6pRYmqKLIrDEMY4AY/FiBFBXdxDMRyI/ZMx5Q1/jlrxgVf2qUIEK21z31ipQwIHUfb
d9lCDlzBVTowpjeXkbR9lEzYrrnxNm4Rli+IyC2kCeLm7feOM9KIqc1UBz4SkNpS71lFFa6fAN4h
ptmtJaYi2SWCCU5DG1Ov7JPBuwPhVZKo1MfSAYi1bWbX7Ij8d2Sk4gioSA7cQQSuHJyIgxUqZOgo
XN2VSIQk/4lXknRqpDkCrIjU3gDixdlX7KKKizup1xx7jkX7vzuFRr6lAPYmibTLM/tJzvD2gf0W
dkgdhAYT1cQre46UgLyfGdbumpLDsdlfpoL4nQzTxDSsCPa78bQW5jImJ9hgynfTFpBs+lqYarzm
ZUWA4vA+9Nr+rWU0OsnArZtt0UoFolcZ2RZ1Ks+bNxFFlwcQZJGsY90ilBSTHEj+AvUcgJCXRqTM
EFXy6r9WdtGOS4rXinfIOnMnXtLpN/isrMnFYY8UtKkzPeZVV2SHE8QGoBo5ogdJcxF0gl0bFz/2
ogP7j1+/115aLh9ODJj8DzEQB7OkQwgYjrGeEYeTvGOrL/ei7wgEIlt7ztrpOFcIsqwSdWve/QVo
Z0IdORuvn8V9DEVPTjfOD8JQ/S4LyJlL34NhVwePpAZflpcmzOMw6h90j3VdBW8vDzNzOmOkCzg2
bIe8y8YCqS5fm9JPy9+d9pkwfPg/fwsszwzw8ZEM5kh5sjSDgwv3voEGGWSQczAfT5WxEe9Sa+ph
KWqIbnXjN3HYuZsUMMGs/lsXosesHYaGiDH6d3nQZ/BhvD8QNWtAoxNpcJxQwOS8ntZQOc5F43tW
mwKYghmf9rk2bJ7DkPrRgOEu1tH9cSndV2/3FGO+kddwjlXjp2XxWcbx9v6nrGZFgRjplalApGay
BDPjcFCnUoXsBQwq+vbc8gKPs4cZuL1FNOHcOb5M02vKzRtiAWPwgxPG10z++blUg0QTzn7m2qfV
VxSmSFPlLk7S6cXPPCRpOKzPd/jueK2kJ96zujV3ZtEHRnSGQpjZwab90KcPIGtAhfJnmJDLJugy
VJc3pwvJtNQWHxkEr0e4K0ar8bwTPuHCsVHs3sJ+vTd6kBy6qzSHbRN8bOpqy//5LKleE6tGEdAs
9sL3nO/y9h8h+s7KMIQqQP6PBLfBVV0RHACWEHtookKb82w+iPWwmF+AF1sO/tv1FOxKHEh+gIcc
LF9bvGxh/7U11+Dgfi2IFyF6WvhzGCkU+PvJIkRRIagFPhzRt/LTE5ofj02k6hjINQsqYsg+7ch1
WRLrIoymMl7HIfwPyXdlOLC0o+7Ga0hqhnGKoF4Sz+bYl/PvL8G+e+J8JWFdK+aflRhgr11aD5L3
w/Jal83xKkbpA7ZgOcIuJY5uGw1Kz6gZRskhiXVZcIjo6UWgfFQtVIm+pnAkRdyOvReQIn4QUjg6
JXdUwuzT4ZaUIecjYzdwJkRKhwnMy0hfHgQR+UbbTHrBNjXW3SlVQ3kt3elzVjwgqBCgFmaHvNYB
YSeMHfU5JJk7483FvhR+QYfrpSLs0Cc9tNDoHsuZFEytz3yuEGqUIKW9cES3FZNFr1I83N+M1SyD
ySEBUGay2QXqLUqO9WIiZiJ9LEtoL9sUZlwYqOMoseUVZVF1BLMoTvudi+dSxo9ptXM5KjHDFpyr
VU1/t3SxD1Epx8dNrUnrDkX4rvwi0EhA/NI+DGxZFPu7yeVWRb1eUCcgX4QYTA9wZZwt35KUZYb/
hZjrL6N/vfqYscVjCJ92Dt/ioyje6HXiYIxKKwgs1YEEBKzpaNiMnjkG9ugHehtGS0HtkTcFW04J
ujZpAbe6zhVzr14UgXZeCy5/rRmu6wVYGt66YIhI3A5PhmTi5Xz1WQjO0OdVncwQU0xz9CWx0o77
FtGZ+rF8UwNoKw3SEzL3lvb9qrWrwX9qFKdTGQG0utPxdlFd+nE1EbgSAcmC7e0KLSQwZTc1sl6a
OUA57d2IIxmnTAceQPegwet1/UpEtGO5IYhpyFiGrRDEWUKedEK9pjXJcr4w0CJwTITqYhLOEDvH
gR5pJZWjiX54bocYWV6N9w3HSPxLime5IpbLvC7vRZam05ZCGqyeflmbt/m0rbVufKCmh10WW/ko
t8wh2Ks7R+D9OTKwD/ank2C4mCW9oowSYafvMRzW067F9YWQt+vnDUH8OYXsY/GHrm67GqVT2Dxb
G1RkOfXrJexLv0HazY2Dt8264QworOv6c1ypnhjLPZoIYrPLZ90xNtxsp0Arm8JEotDXUE3sBbb/
AW5cErQlFtzcSr9VsmynABlelOQbHCJ7kbJn2dsAJzuqCye6ItHy9jZ6La6qO8L4zaSvu+vpEIGZ
IvQ3kgY39YLFHqLztyZ4u6rDIVQWHqPSUQ16zOdmQX3DRmNpwC/hB8ROpKsSZUvtiHUIClZ01Zji
ZCaKl8t3KK9E4Sjq3ubsruiB9s3ktOJTK2+u9bEmhYwSzfIzWKY51tQbSEpYziF62ml5nZQSfAR2
cHH8m8tYeki+KxnC9FELq9V01dgJ1hvt5N/macoadL3sEr0cgnPbsGqXQugvewmOtR8buQfkatho
xU8YXG3n/pYBh/FffOpO8MsBqGcZIro1mOrprGXEOhaxdUKe+aCwkcwOIgz78XfawV9M28SluHy/
HnES6zzX2htWIIdtiDW3OecdKwIcmWgM04ywfp1gosoRpWwumNX75eQDeNvwMny2R9tzPMz6/XgA
Bx3Zr7H3OfrCPa0q/1oDIKNDq2Qu30rDOv7tJkopmi9F/8gWxJ42ekBcZJ84fwTEfmBJuxFj/N5S
2/f8og55QyFItzjAtOr4qo/fU4RnWuyLmZF39JEuYdNusjXy3RmoQikEPQRUBCmoafa26Coi9XeZ
bFLsuL9DaxwBCzQlNJQjUR9LXo/UM/sImZCqyHpIzwf3b4vOxpiYxPFXbLUUcwUY+MV+BROI9cSJ
UXvGxohKBi4N77SKk+AydPnwfuP3EWctKD3uq+AchVnF/EjXRA9wN6fgCcn5chMCjiFEIJZ15U8b
ONjOPq5ida/hc+OQAt/SKiHJkb868gMptFo1SwRUIwY+C4Mz5qhydp3Z/rW/JdSEHG20VwvA+92q
F5hMnfKI6LsOcxSGQwYj5IlC+Iw68EEK80GP5PqR1wwgOkPUk3M1Y4OtVKBYpw4YlvCN7+4x6TYC
PfDAditQTzyQqRzkGiA51eH42gV0SMS3v/GzVWnJ5y/1gDEW47Z7D8Rc9wwYgsqXvNtnfd09rwCe
L3eLRE0vgyYs6Qo9e4h+eq3WZqp2lv38zBJj2hcshZ+RUrkoAmdbE39AT1Bb1alpz/d8WFTZsBbS
6vmR/YTHc2XhC/rVEJBHE9x6ZKDKXeXmFuM7oBJ/M4vBJVkRJxcvRjAywma/eT0qqjnZPNSvke4G
OvvIra8HPwOL8l3dXVrB3CwtI3LdyqWqjhGvqLwamEWv4PiEkH0R6D7sB8gUaYJ98M1dPEPVHikp
wAYo3YL4am3I5OlReWJyiGTzrGkEyaWlmKOmKac6fE7fTdqQtaX/jp6hO5NQz6B+bQruJkxfhQQF
Dx62Rm8qKQ4z8w5T7zWBGTLIeVVRPI4/Y5bodz+798zAWu7CrwANo1ZgTJ99lPIRc48WegtV4Oly
hU6uQiALpJUczn7z09OmU0j/44pNuaWOEGDAWSx2qDHN+bSmAygIC5g4fDjSc9bTLV8KynTdH//7
jkaOg2Slne4GsvYAo17Kf5BkRA/mWVmabBmdpmf7qry15Dv77mNGP3/bKNZcjzmeZAV3kyRTJv4x
yrdKkv0s7gPJ2xEgf/3xhm9gkUO6hwUf2OhUdJsGI+ql98Y1UinCx85irg3Yq/NOjDINdWXiPVXj
/kUPs9nf6eub/OA2KJe3zIMy2ofnB7BpP5ECjl/DbvzVML9gsCrUYri4SHFISVOVdOY+q7IyyYpG
ASIw8BDY3umTuv5EofESaqhGAwp4VJXqFWqAZdEwXfyFij2o6AgavAOvb3Qpin4FIclLtuFGwGxK
de11x+b2fLNHlh/qiAVPny7ZeNd8zNBCTsmkK0y3MIaLuss3huq8pg3O0ObL0xTah332+49b+acZ
3JsorX5+H9NrQJgeytRB5d/zFMCBD1s8litk6wBKhiqrWFavJhGnq4HFcRuToABfLOJkuFU18P3a
IKqAFUvcelNKJ9WvlFqkaF/jQEykQ28dn6wSy0XUdzCkgCTjdhDQHawKdfXrI6niwXPWHls6vkHb
HT0gKPPMk3UoJkB9/if+MAEuwg5yD00y46Bm9ofwTjOjRuB2TZnQe1O+zlV04dtVhvGlpjdsl/Py
TIG/0tv+R5hFE7VnXPUgwxBKp2EPmpObiVWRYFsCmLDOUzMznrdw80gdEphFY2lyRx3GPCNVWkPK
CCo58IbR/kk+wDtlMiQUqvrsl7fW/Bj780S/cAetO6vq99n3q3OyGJefcT9CLCXOKRWs4nQcwun4
WMrjD0i6mnC/9akqMvlGr4UMSFIE61+0YCm2HI3vW5Ng0HUMluqfFA4ZSitLkY3Z86DnbzBzVrM0
T4zsM4eIgQ4+jE9oO5MIwR8wTqPYZSZlnO/AzGabwad5ZDYqiJrzgzTPj2fNQFLLfjjD0S7MJD4S
nUxohNhl1dnX2vpcNjZ757X3n7q83dstRJkbIdU3A2rjNgX3AKHXz2VGkVYYZ5RrlFyAINiyPX+m
vJe2BaZS8cLbGmX/+LDbOKWYoqBFqJF0w2wVa0oGJuP9Zq7B9f65k+zvCOpKiYZQReSuQ7HvQq8Q
WrKnmtNmOp9RpjZY2DTlYr/qsXPWjHRvoPXDM7i1XQ1ZtDDpNkwRfi0zCK2ashmRF/1pGdzqX0CG
xViAtu0EmorTXcjpOE+5IFapyBnZLQ7iEP4/ALo4c1MXHYani9Ky9rPoS7UxTeLZXuE8aTYV5ws8
NoI4kcNjrfe1+iM7elfaSXzoZ1mMlb6nSOEkE1ibWU96dGRCwitxAZRC1e0Rym65Le6Odh9D1A38
N4OhubBAUGfJtqi3ot0Bi+IrwXRgffJc+osX1iRYkElUA5o432LTjl5QxatD9eIK6B6LGrgB+5wh
ZIXcLODGorAZclWcTUWZEYLG+wFQRfNgImq023ZWK2syfgivgG6gX8OFuPzvbtvUPJTEv3bfnZFe
wZIrUv0H/ApwghUUclZGJ8D6bHOD2cM7jDKmkQwSGClyuBaYgA13Dp4ogulhB3XWaPxRKyADCP2s
Q7ZS93MW+3DM8yFKKedvz7Z19bFdUgkiDUgHe++r+Tim9TAMpNFlRDlLlB4z7UKVvdLPkWMvhY2P
IMjvfncqi498cxfLhGfK2kgk/8iILTRLUaVjUQDQ4qmAQjJQSqYSGXMHcQsU4xw4Q2oumuUl8+u4
se4fPLUY4c3k9f5blGT9qXr9VF9eEtyLPbc5alvaFK68zGw+Ia9Ib02ZN8ETm4uM6DhNBLVsmwip
Bat28HN2DrlHlFr644ESDeEQq1tnBRGqdEKD/4b3OeeJ2NbDIqrzQ50IfW2h+xR92Q2W6l0m2ubi
gHrVk64FWVTbqiVT/SX0tSWmFD5xe0ZmNm5ECX8AkWU8t9BIylCO22khzSAg6dNGOfuPxxDGo3ho
ch3ujopSJ7UIyfjyL69iLpeDxIhSjzPC5B0y5Hs8bnqGBtyqolpNQkgpLdZbZgapzFhjr9hk62td
qZ5Xx8/3a3yrj4uzRYI7OnLDky13g0sFuUysd9h5kRh7I7USi5v7DP346S1CJaMWslVTpARJfmyw
w6DUs/h5L8hmSj7R9mLIhrGDZdhXBR8pi8gbbAoaRBRmLKLoCr7T8CzWAuvcAQO/qsirEATOkEQq
J6rRFkmBz1NN0UFlPSirRZR3DGHW59M6m9qyvC+Klzlx0AIfMGF7sjSNx3yAUQNK0zXyIzEHczds
XD/OdlgBDXH+Gauhn7NMFiuN6FoUMUTudJ2Or4mksRTFcc0++pnG7hrrGZSgwxNNsGoWYQcrMSCV
L6xOD541iec+2lZAmR8RPmPw5/+GIoaToCr4FfnbQti+6xMPri/OPQTG1Tbwbvw5u2DrT2z13o3/
DQCWqp+e9bKS25VCXAcuWH9hc7AGMnGPR0jnCvsDNnza04FOnQ+vbTFlXibl1ABQlWMekaWCY/8V
Xr+AegFY1Dpx89nUqEjoxYNvqFs68Nury1GdQyQPXTRpE5wPLApJczFss+Y+IvoZz1bvsMSazewk
IxRAx+ZD8p4jUbeCnbboWfY82IRHJ82YLKWEJcQ8fuBVQGV+uFrK3c1ab14cjnGP/FjDeobB/VBy
XivDkWJ1EQCXFgpixv8ogpNVbwPfL7zkeGs0bQqJbhoTc8nGBVpE9YhyIOOS59b5e/RGl1awtStP
xRZzPafFpaytNtlge8JK+bvKH+T1losIW4WR6Tj6qL3PBIggbV7m9b8ePMKP2NCQ+T3bPPnFBmbq
RyBVOARuADNYDkXUkkaOn0fGU/QSTYWNAUyxanHEl8IxHnv3nE/Qb0N3WuZ7askJU5qs0V4jeEQk
9ibDY5W4FznBAtj76yh6cNxSbe51bj4qnxhRuyalAG3/I8/a2c+99Bpe1GNjQRhk0odR3dMvyzrA
2Rga1fupIQuF/l7Qc3mP87lQ+/lBA8fmvrraI5nnuGIVIjzFM+EApccpmDErdJ/RYNxRhvJPdMF5
HQcsxcak6A3VA2/1tRJmSUdUCL2yq4oMGE9+unmsFv4o/x8owE1rui2N/9lccXMQHc4j2SAfcotL
ABNoJUxkts6Y2IRlaAHmc/RUduLp2cpewGf7IBCfv9xr++kvgW2krwzQ4n1zigIRJvDOEpF/oq87
Dz14D5mE8onAWBBFyj4yRDtQxCtPQ6/RQc3HnsmrK+2udRf/1zusp+OqaZeBPtie4iudsXSqReLX
A06P/BjD9g7IeKlYh21e4pLdgLyU/H4pQ9W8Q/4QFmoN/qOEZCYxcwErYsuORmW1KmiJ/tn+WVtP
IwZynWdNympiIubw1DKlw1QlLqhotoYU3g94dAGGrp44r+xYiwHxzSBt/d78Nbi6ze6ZVCubbQJJ
W++cengN+lzMLLrrPgQrN01/IhQmKr8jV85IzwOMIEjeiInP0/gpRAHVa8Tm8y17Q6Zx6XNqKv0i
hwM7iHuUOAk9IPiPfsVTzHbsmKxW9DRAp4/YrnQqjLi3elzkvaqNLz6Xuoqy1dh94KAWA57vC1YT
kIGd1hkwuiHIYQ0PJV5UThnM0KlG0jlPGntqW10M0/jcVQq3ab0DK2o2TN3+B7WxCf/Qr6sQfJZ1
dWH+4ubpSA0DuUv/hKHtxLHOzsWAd7uiWqlcTSjNsrl7CSsrPi2CTqaQlwRGSlDDHMb/BcEaRBGq
pbes3DXt9LMhurexlrLmbCt+5MawbXTTY5AGvxnf6QBZm32JCp3kfGHAU175+MnAEyA4Y19w8dB+
LIsK2xksqXu0Gp1bIhLMIYK7ESALXGx0Ko95ewE13dpbmK45KI7Z3gbIB24opc9//l7hQ7/pjcJg
0h2k322DhlqEwYkNIJF5ayyEOLiW/6sXj5a8ItndqwyhypHdVgDD/myquahcpGdtgV9JsH1R78Uz
hz5q+4pwSV+0yiWQVJ2pq81uEaKt12J0x+fl5SUkddtU34h4/6cy+gohgVGmVvYDH3/e3yImQevY
tO5Z6cpMoGqzvq0VLdi0Eo4pbXxx0fPAVL0eY3/VATjSad+2NdM2W5tc8gHBv3TNzl05td5bODKV
7jJ/3qud6lY12j3b5q6swJ6/bw6QbA4LRZ1QRereZVxKbva/LIQ6rYab9gYwvtVaYY2QhfJzx4FA
NzoiitXmF80/nAZENf3FUcIO8Wa9tN7ErqHsrE3p3Nvh1SFQZp4AzclKYuR1LvhMzoGbWZl/Icyq
USZoeT3kxojUZtuT3mLOvNy9fTkOA57lvMlWyeP1s9LSXFzdT61qlz2+go8MLR/LL2/YucmWYpme
6tp31Hy3AHPlaRW9ryZ6eeLHazalLsYHlw583NktevRHEiznsfgW8JqCnlNuK8gmT6MYDh+Il4Rw
r/WloWprGCmKy73Sp2lKKDzJ016fNYxmAYgmwMNUWg0rPenCqsiI8lJ3JSw0Wn3nVvvYBD1jBYU5
1BwmRJ2WS3PPAIpMeMoRsal9QxbG4navSk+8vGejpqqenaBBQCo6PZEik8V0nN1bmZIjEXLUGATX
IX7bfxr+kQnmCHFAk8Yv+zqzahdMuV/hIdfXZUd92ZqcJIYIBuuMKd0sqBiXLsIdvhg15KNykzlq
iLm8JoC90fRcHRxP8FBDvogX7jvFV0AUtyZ4jXZ1j7kpIYpOd3ynRavDvRjS8LNAKDXEwzaRRZXl
k2Ghnjsv+kAj8+H9O5ZD1MbBgTUFajWwCua6VkngH8v1uq7AY6RXFW3RyfH+pyGDNfVRFZrsvFgl
xXUj7B7/WV6EXSXUFIKlMXvDeQzAxz1T57SM73Tsy7OzZBUjnBkPdpJIYLxYxraoWt6q8fWGX+PE
7V1uRXQWMnBV9bDIEsY9PewZzSRWU1sx8S4QSAVrghkRULRTDHDgY1jTjZKjHUsLHYxwds18oryD
z/0Q3NCUM8sJaLivnAzi3RUrT/e3GVkxYMdmVZLMjYQQx8i4nYRsxDt4qWwHybdKCRQs/B4j9C+2
6JAHdoRNA7yJ3qkEnEhWEB4osxZJ7+kZm1Kiss3dbsEwpus4yHqbFylve9rUOtWCDpdlkQb9jDSm
wcMY+JQKblNEwm7b33MPgIM1wrfXgAoXvgL3tb6aGBnTX1ykwkND96joPql7htBm6EKKreXiSjtm
qRLbQoXTdr/7V2fp93P20muKBToEZivFOWVcJysuSGoDd5/EcQmz4kpQqVI6HZkQJQZ+6gXpbLk3
Cgcq7MdjWr1ObwRHucJOV5/4j4c23ueGHs4kEGh4DfmVD4Jhxyj1oR7bvsJi6JOhQZMR8Obzi5TI
+/8PRKCaX6fR/gCjuH4ImzrCnMhS67iIJDV6t7GiHqkDhEyp6eggL/Ov1/zxCkK80VAcyNGrf3FG
qUSLUGuNGklp4sPkO1wYZ2rG01nJjKZyZHNdnz8SICuUh8rPxJmF7vFT3TbXVRHQZEOGVhFTRp0Q
pk8AgYBQiAALfS6nVyN3fZzY3CoQzpdETQbW6RnnVDe4bRBTFtnTITuinFGNyv+hXvpVFwVsQ2av
1eQPfDabNgVIPvwZK0TkjWqomhps+0OCKsycTu/Juzvm4XIkKbFNACrqz/mG6z0Uvw8Iu5e1vIe6
787IeTE1N4tdCPodhlk+ofeYcmopipWqespMGEx2PR9A9+Sz3GuEHijRkKSG/3Oxe1FnM1NYGvmw
cuahlQUSGNV9dVAaaNVI9JWthdiGmeP7BmiDMDT3kWNWN34zScubMf7PriM/N2SbZzDrKRhrRLyG
uVT865vvGpc+iVxdEDyy+HpCDQIelDIAqe9AGS8E8lNjpXZKBE2DB5B7G02hoAhScI7sGBy1vn4T
jyGhDnzGOQfNRpYlJmG8MOA0xtSuS8sjs7P6PWyUjaASTeDcW+g1j32nlPrx6VuY7fr37SPoRFg8
UAQTyiVntOaIvNunLQqxZNcR2SBypEcPFVpWJkHS6APgbpjl3UWTb3KNWpU6I4yWET/11NAVm9At
B3B6jAIAnSFeA70MBl/Vld0QMygww0oE45cxKBwXUCyfbjkhacHLwL7+LKSlkZ+8RNFVyGCPuGqj
JLunx1Iw9MyMsL7oTYnuzIbVXtKf8OzUWSszrr2pwiRomfB2wUWJawrmnTBCr5FPh67NKvUQqF8G
73S7NxD9h+ncJqIDq0C6lAzOtBXAK9o+L0Z2R+oFUj6gFBbQ4ScD1KS5ZP8wDH2CvhW/jyVl83do
iA2HDmKUtkvmwKFpbbaFEQs0MFOS+xvIyylPEST20X+ZTcMquZEpgMuI735reAylQXpfXVmgVdWk
R0L+MwoOCiTJLPK+o7+Er2rpbZO/14E3PId5NleURI6DuXK+jVJfvwtfgnD0AizsYDCchlDFSArJ
5BebdiB1+7RjflaA9uCkCP/T7t4JrkVIH+R/E4EK0fb5VGHA2nQog6s0szgQipKAybhvR4aE6xyu
Qp2QDruX9QKTPDdulVHR4Rb1WyVTAFHGf3T/XPdG6gNslEkjybv12w0bYhjE1kZe7tPtFfIBXF/1
Hb8veCkhSyzWHUeBzIUJoc+Mwbdn2MwmzB83n2SL0zrXgIDZfULvacbb839bYsNPe+tdEgvX/dQF
nO0YO6Tw2G61IOfsOYg/go1ewpIIybGVUDCqWaOcxq7bpxvkZ0MBDAb2Gyp48JCzS52sZuUQgxgA
cPwiJH0k4fSs6Yl5h1sdOgLLubETSSpf+detUrIIQKKTXPno7Ih15e064copqnIR7vpQNGKZYaW5
Q6dCbVpCvx1GLHSKjuo6MWg5FajY4HIzUaDXJG+R7Nprb4iy94K3i05WdSUp8Uguy0UFUNiq+uQ2
i2f1cbX5swwFvMKoLxugMyFxcoFizhnsiZC/YLdP7bGliA/KEqCV2B10TtOTQsnqJTFPJYQxMXUo
bjUpN2uemmempAKVf2MOg/U4ldlFhPuhDaLZAkdHK4PjlhbEH7nsQE/v60yVoes+1NChrCmwJIn2
pXbx3+nbjDPQZeBwC7m9PI051K0ELcmhS4agIQG+MQ9WMopYOZ9YZnVh069u5V7ZLLjW9zBsYl2V
D1mErPyReT5NCL+49H6HW2D7yQVSGppKiSyP+V+CLsHCsp4WfUA8k6RLt4UjWrsH0p8O2mVUEnAY
ojn2UirYbUxP9CTAAqzeuL0kV7HQRA66GGuC3Y8p30XlFjvS2ZUafoDMwq/HegJodJk0hYVuG2mJ
wYhIyVCX1nAS/zGitwTQBxchQ/t3jpqieAusz50M5p5c1VSvBSpeq3zLwpKLxDdjAxs27vVheMb+
lii9FpaTB/cYCnL0rtWWPczEHagQL9OuCUkD0BjOLG5P3M1ql+v9MvPeWfdkXRO07+Kl1w56bvbq
eqUbzZTEPTWapCo0KX7gjo25ew4OwoVmmA4F3cWTUgIyEupnQB76YEGCRx4g38T6qd3f6XhNkmj+
3BeSEa+Py6WWLlitFWESiaP4iYjo6jy1JA3g8lagnL+O8DK4lmSetKPBNX3gJFku69LRGWd1zChd
VR5NR7Qrng9nRgMg1QN4FBvyTRMJKB+D/hS4794lNZaaoFB23SIz/5ywXjenAlIv9zLMeKtaYf4r
ryJEGV0RIFIQ4qc4vI7wRxj5wcnwXcBqcd+T1sbUiYVw6tGpUM0ZtKHaJJSOoO29DQ8HqLIDx45z
I2l1O95tPw4GWq4Uk5E6E/B9xXsYuOGdec/iYOXVmfc2dt52qOmD3Cho8lJ/MZmLxPchCQXzOvKG
5BhP10r0seVaxXxbP4inJ/xjcx4MEmrY22UzBM9UbueIRRL7Ixz5WnO88fHiNApQfgA/g3azeYth
eTxROUyvSovcZyD5N5JDM4SNjqlIvmPcDMUQu8vEcRGE6BwV7wPyra0YFLEG/3QNiReAxAQEFuHd
F5VH+uKuHxUCi13Ug82XE1uzmMGEGTllS+ZnHxL48FO9OBuSKVy8BKibaEYeJ5/7jF7iCJEOdEu6
4EeJUCl6/ygeKs77Jvl+d4yD0tXlZPIJI9rLhruWIpFMFvSpJ04Uq/uIFEpEj0mW4shV8zRLFP4W
CpuaDRWLmFSy03/FJSE+BxC4rdrsqGNLj8GqLXYgKd/Vu6yCEEd2g8iKriccYDGwnce4Lv18v6c2
PN0/AvhsD3luyFfHrrfIO7UO1LRAFifA0CDcFA7DILz4EKO2Zn8I26KxpU2vX0foB3DIosa4TkXH
6dAvvfLwnWk943LKz7UH+9ih2ESc7WuOkNIQ91hR6y5S/oRwTF1iZXqKamtBOfQ2fgflUBTDFySj
5kip/8dqYclxGUEFBxG8PXyNsqfUo12rYEBxMKM8iyRb9SO02Ec8aqlJy00ntfGC0xDps6HBp09m
CEc9ndvz/DIHRjwe7DD94l9REBprheoIBnoKFeX/d5GdHc8JTi7EPH8UERw0/D9y7yJ0QNIJBKI/
t90qYp/tUtc8/GRQuNHDZXO1MebotXlr+/t7sASZOxCA9KmWS+rBpb/ZEWFAGSZ9QsWZjbaZBkC9
pQpN/SyfcSR0PoELaXXRs1KUZNDOs69EWfs1ROTmp+S0Z4Kn+kLztisrpa2Suw7ENMs9V4HC6Dq2
TVN6nmxS3zxGEaCxyMushNFn/+p3fm9J30J6qUP9+hoNScB7WN6gST3zLLHlSSccMgdhjv/z2i1+
UHwuGSCAB/wm4BwRhpACwo58zuqpa3hwYoj2bNnf5PohStywsG06IjpVK+SkTt0eue/koaR58rsr
xGcVUzyQR2B7mFEQ+5p7lT7xqPGXajIcNAs0co/6qUzEbUt8wKYKipqIo9dx5z9dgVQSQmiOs32N
eLG5JzkbCv1zsN2UtnzFDU4bM0Wif9ka+vOPiUEJDdNLqelpRoo+Fkl2D1DcCaNWZGmJ/630PX7u
UjwWbUi42L0GlOFcBbuxZiajottg5251hH319DQdVF7KWxYaCZsZMEnc5axFQEduVsyzTpEZhqb4
qicxJpiAdQn6h5VAsu8GwL7bQU8N5EEnJBR4A0DtYtqYpMp2SnnDGcajKIH7qHxFhr+1byJBKuxh
qnXwf261oFQ+4cfAPasz8imTkcKQnLjD5ZJdJD4Z27mBHTh8EzqwyfgiaJx11FfwoZboCSBJuhm8
WgXi41WW6n2trZT5tw755sCSwIb5NbVwM7y9fmfLMSTSObbwFSU+LYJaikIx+8OWydRPJt7OKN4Z
bc/kbMfR5ls0MyukS81wz8/hSSUKgppa5BKNdYE9pzxvFLHyWNlXw2hlavrg3oKMNUms9PLqm2fd
37C1WWoC0QeMxZyrRqpJXw92Ue5V6bL2p2RmlwaXQR1brCVuszyNzh/llnhbHF1ctMy6Cw9E6Nur
XSVQhdSyY34WqN+OJ0B8YEPX4RVjc8O3bi9U5wbEpgHbBjiaEQv76ARFfiL5NE9Zvad6dIazS1ak
omusIMTp9U6Aee+ylG5+fnaI/ZiXcFSTZVstvi9FVLSdBBtVEREKCLclIfF4w+Tjvqr5mXlInJ7g
rEwD8PXb3njWU1foUW+0/GMLjIZuIx2ofrBtpMMjl9PGzQaIXLiFeCA1ncoeZ0/dlqolvg1AxGij
811G7QG2fVlbaoFu+ZBieHE7GCZivWAA24O1Ct0htNSQ68tEbWwCKua76/XNrWxNbfGnsVcDuRfN
ud5Pof/zKrK5vhJs3rBs7E9QY9+TWvRZwrdjI5fLAxMVqlx35Uvm18T8xoW9V5+SrxANpp1PaWKn
3PAs4s4N1L9ZhfG2OCZN7mYRNw4iwZLf3dVGuD7/Avw/Wv/0XE6Zr3OOCEzXtdAn20KvreMKCaFA
A+y0RDg3qa7jSECCJ2lj/7hUGRlEVl+iGeYVYhaJ09wWpd7fX7hC1yK601Z8W0zfdIvi1wRJxySh
xRGWISqUaJoXB4F1XXFGZUninUkF/3rVEJm/2I/o7Tt9e2hA6VyxXr/+4R03qo2AApUKATHUMcj8
ejfAMPML+YO2HoON61wvpnpmbTBCl2hGGUU5OWiTypGPAdot5BA1HE1mGC8+1LAX6SkhhH6pw7se
qVuhq/i6LlzzilX2Ga7xg0R0hL2SKqudPcSf4BbjrwFlHSC2Qlj8jm+FcnxBXiCpIs4JIXI+aoh7
TiZeaFTRd8lzadAK32fj3tUm1ltHi22F3C14V2l16mYIzaiM+lHBGng3+SRTdm58jvQ7Yc+oZbSW
9mF6DPYEF2psG9L3wNBkK8TPmxc/TEJJ+rdZAW04HUMb6MKrUbZb8v4SQL+OOuwBl+yWJ4h8W905
46lykgLCzBKvqN1i+VNzsiUSaNCPILCD9iQVNj1mOE9r6Usa1a2Qw9TOQ9B+6HFpZsP7sOpDVAc+
Bc6guJeCGChuYB91i3EPCsOdk5tnQhUJCs3+WblpWiS3aDsaaoYkSBcqUo6aKSR0NGejnFITP0dB
YaIiZc5x6C3wxUsCa94/I8VRP/Qv7D9c4Sdc2DB1uEy/KlYTEgEBcG3Bffc9e5aKInBauX+4Nmaf
nGQNJSMvgFdzwaKvHfMRcWBlI9+R29LMSFhO/neV6f5nR3/i6xwP2w0/8M4d6T6UaPIXNmITc+WR
KAKMOmJKyhVSLz57EajmZ/vvR9Y+xguPZpCPPumdIZdZHqkhQ3L2NLemsGdxhbpLRBBOja5oGwUf
GiR5u52osyMDPUIKAvmYUyqHj2+0uAoOZhjdW4LnDaHNFsLhWi/Nn8y5NmjVdCIdIX+y8uwX61Jb
d1oASQGFjXbYjgfPpopNq7DBe5P7txiHWLVfX6pgLKE10Ltdyqlc2h7vsuTlflj/1XEAnjwQB7DO
o1vz7OWeaMx4chbrbyRWVandrzcTp4ZatF+3lbLYbY10Ea53YeQ7L8/W6l8hbxlWf9UMmXlBtggV
Ldrt0O3k2VTNiJlrCS+LNpIAm9+0l9y8J764eb2MzrapIa802zBRxMfPqvHmt9s0Q3Ly7DtYzd15
GxwGqDfNRuiprv/72gsyf7dWlyGlwzJWK/r0WK4GgaM4QzRfqpaG1YVDEWgI+zL20vLneuGCoSzd
iHRcEWXmuzXuTXctH/xwP8Li9Z/L2CiPYevKqwkTzpobFQz62mUtuRF/fRYo/nGY7nbwY3rQq8+1
2A29YKwl23YCWHIUgxoOl9/xLqrqMuonTn1fN4aF/tY/LRac5lntGfB+AKE9CpyJa30pCM4kvVfn
Y8YA/H/LSQptmZF2iL18WOcerccgmHZ91x07TXKY2RvKtLLLMLB8XiOyvt0C+9GooAPB4X1uyTK4
h7Q1MHiBnCb2n4A8Qm+6q8Z6n8yACgBb9HvTEHJZmMrulo6yIOhNz9fXPHd9XMYDP9nTjTi25jUV
qXNvEXJNN4mOTxc9nyFEazeWFuNSFP42X3iBDiAvCtYlQbkphc3qA/kXf7zLUfVoIpyII7XouSKx
eMbdkcZ9Jk/oc7zKSKzJ8UoR2K5LRRYHIQYgd1HLBW+vp2KSz/e/zSpUpkxrCh+OvtrdO3sGopNM
ycnElczuL90UxHb8iBlRo/pvQaZz4tSmP/Q3Qi/VgO1Wt/X2MWwwP8INBGRxu9G3Ypc3VA3WWO7h
4miVqXP9nonbe/Jnj3AHqiu+q9OdtEVjHHeW+sw0Ndh/ZsOJOuDan5+4lt2TOMAlPfLGYjksmFQ+
uU6XKQ8Rg8+BlU2ICLjtqdNuvWfnZAaxRKnYjhUwZJ2l3NleoIochxzxPCmsfHTdajaGhJacR0gv
DfziRxlrl9K3NK3uumbhoKlfVQKaT81cMov3E2lMVozBlEKMJ+7ctQwNPa3eAQf+8exTXnT5qFqx
dpmaoLSfwvcC+jl8KkD9EMIl1o1Ii+FuRVPStK1SafLaxFqVhQEwbT6VVPXsDiSErkHUgaRXeiB/
LM0rci8tPDTGYs3BaCvg5jDxH5HsOnZOuJSHTZpgtDE5VTxjkiV/NSnDHTU3WwH19d4dG3kTV4Kx
nQUcoecX9ZxeOTcfSm/Di4SxHKewOd4hZACqJghtv1excD33sGucnkETCawR66m8kIneOr1TGwYA
dT3F/8kyx7Zd1uvmMG8HQWJwXviGlrAe4CWQ8o5cRSvTgtvITXIqJ5AaqO0nO6oa2vJtRbfcN4J/
q2sOyH+M2z7wU8LWbt6s8ZtjxKuJo8J2ztZLcbiYxJ35nreQVFwXAgY1yQpFGhe4GcYsfJd0EUQv
pjhCu/qUrcRrNfkk0ZuQjXZpMfW4z6JzInzODo9d9hf2HGp+Al2Hi4nH9pgUdStqVZNYgj313n4+
cAZ7TSM+IG7hJcKcfQVrlo+lW5WLpu2URyxWtw/LB6q/9i5RkHIVe7D7Ii0+luVRQcscE219pTLc
BrXnZ0AA50bZNXJXa7NiwGw366IDOhbbID61veUMYbKFtU5YGrBgXfAfPCDoTKpDC1xe18ECSaD6
OKmXIu8Nu1+Xw11cBSlbM/gULyS0n9wglZ+77/dSDHxTw5NK+aN35ErXNl2EKjaJCEF0do1WFmRG
3Nn4fSq8JZcLhnE5MRg3F8oNEvFSx0ysgerzGZCk68H73cr4/wX4CuJG9TLaFbGDIoQI9yIfTUHf
cJCip97hv7tt4NdJxnMVG+ILu6WDylFiy+9tsEOFaZWuRJ+rVHdOmIq0kbVQVLAnE4Ogp25tSwv1
4lOmTXAk3DnjmJeXBhnr1e4yL94YpTbHZOBRTa2MpcOgTKyzeCO3b3X+UQAL3sdQsbxBqAT3IcNy
BQmIdqouuhLxFSxzjjh3VVFz669VsdXnH5rUlWZj+vVHToB0+smFrPyHlAEyJpVcUUM7WI8O4ACD
OdxW/boFADEGN10m8tbpKa2XRXqiVBKj2bUOuDxSf7PKbtcXb4DIzCwJ2/z00cpCtbGXVPy7EIYj
n+nFOvjEPK9ubwpFASrGsJagVv+MlVTGJoB3pKWaB9DiCFNEHnng7v9MLw/xJm4NVjt8BWKR2mHM
If1AZi/sf1+Hc54ugu6vkzw6Ra3ij3J0cEhepn62pYoVvs/C196iqMDU3FG9CezsdoBMcbjjgxTw
a2JswfPLE6yWlBVvIijTroQbASO9wTTdbz8y1bdvruMY5q3hHpyBbILgcZ74VgJW5sm9yfhguJc6
Y/jSWukL2GMFUAAZWEsoSxAePck4cNlE+sP/HpDpasZkr1/orUbk9FS7fC2ezQeDjD1Xv3YjQqVj
WXDp2llL9nHfC/iK6hYGasKo0yWff3iSUEKGPkmxal3no3X3jKgW9ezolSlFLhd7J58I/1Fn0dAG
IbS5D6acLGdqItyd4wlbvwV52W57qGEPd0S/KOlq3GTXttVihDYc/cPbhcQh7r8eCHeQdyEk4yef
mrs+A52GihloYG28kOvvY3g8c+6fU7/qfGCNFiHgTfd/GxWulUm7PyLv22HK2eg7yPZ+EuO9LXUF
3Q7nHbD9QXOpNFULOzHmom5QzCwMPd85Ue/W2tNNd2CQpt0WCLETmLx2Hk0a/S/Pj888gzkPfaRm
OaOGAXfxwjRMERK9R/P/hYXS2xE6+V02lpuK2YtCkOW4VutrGYXb16HMFTDtWc97AjUU0rGgtogD
Bo9opPxXBcwmH/rzbqN99pmCzWU4chWoeeJHcqWmU2G8IyuyzvWgBKx6PjWjroimjiISZ6FC+IZb
+abdJvlmoQyCEaIH5dJfWI9LP5xpArRE0W+V7Ymu0Gar263DVGgYE4AYnHIdDU9IOfNpLtMtRUWK
xUNDwdrAiITf/xMdmucNUA8IdKJ90hEoyzXoWuMiUuK2CUunNKm6+nCj0/Hk1JPEZq8xR/D8pOxv
BApVgELzLiuEub/o5oWe6y5ffudE99EIimAY0mUk5klFK/2l5Ur6c+V3Hxn77zqca0aea6D2iW8s
yvIbKMfQfFkZe1Y+3ARAqV+jk6pcJ74orxonsoQpZWoSuLnrFCWMfrxfXU10V9qPapypX+Vm27Kk
H1OhXQFLARv/V0fZ7ZQlPn1sm2kcsxUB1WRB/41AmEgBe3Ed/70XHWWL5Vu+PAmZlKpUac/9lgSz
wqnv48C6u3BSWlDAq3T3YjRpHPqfPx26d4NkuU/JWBG/cO7EN1Pzc9XMCrMTTvbv3f919crJzJch
mw1aiY3vyU62DLXN/JF93ARvwv5dghittF9+3C0YiuF7KCRa/1dKZVC5Q6BUVERxZbpxDDGwvpYO
oKz5QLyy/Jk7vprx/U3b3MQ/JqpbxKtCf9b5dqkaDEXimeUKglIg5A75vC5XCcQMIGW8djWZVRLv
q17TMwdnmeQBhub2nkFqmQcZgq9UP7Ibxku9f9ykX+IpAIjmx9lIbO+8mNpjymqzetDjwBeMR9mD
pqS9J66oAX3ZgW7LYwY2xLmS2ptbZDYHNJz3PBVGm9k14Vw8DlpZmLn5guWd8OBtEAmoVgOoWET9
EYfTh2khgpf6IM7kqO6uwHGf1IcQWmkY8RNkUDZOErbTg56c8RhfQ9ZhptXKS0Qf/x81QfAgv+Rk
dNvySK+Cl+9IbwfOkubMjwQwgc9tK/m2VnTwGGEx68XD2VruGpo+nh2r1w18Dr20lL7pTu4+vrDe
gai7bu0Y6mkHulDivaPXv+CIdpO77WiOpwEEpH8O9laQuGJ37dEpZY/nAG0hJc/JGc41mymHC4cR
6ViMghPOVnCp3SIjAgN/1wpcn7idche4uCSZM+d+QaPOXq5+/CZ1P0E4UdstmEv2iLp1CQreCLRD
gl5RXEZ0o1ECN5F/6cvm3ZWVT8er6R1WFjztIPMDs8pbhXlJDwgIK8baT6q5sHHqSeK2g3pgPRn1
edJReO+IE3Q0Az2od1xS/ruzU0qFJwjuHV+ZNxZPMvQUYBoO/15S4Kq+i+iC2Yq8C0grKmot1/AS
Qwssl4tcB4wn7FyKam/Mb1JhxQOQX6cuXRRWOZJyTVC9zVCQCDLjG87x9nJYnnNcnhVn+GcdoPU+
zf8umyM6mBqH5YeHFHfHZ8fUoRnxoIeDYGZJJlOcRHB+JkIGjmjbtTJufk1FbTs0VYCncq+PdSQl
LHM79AfYjzNfmJe12fcNXy0fNPSZHTv5j3LGjHmy46OSIbeaSPCT7/8ueYkaiw3hc+sE5dzdP2t9
Pm5y+yN63C4ynrxJEVYKCNYnIoameEbtKs5n5BXDJ4/U60hKPQSFOGBNKH7F6Sh7FPQyalT9Zrnn
askUuzzoMvszF9nlmHZvKyS8J81cspfoLpAW1CB/bpJ4CHPRvUSLOKknZTk6sT1IkCTu+LadE8st
o7V5fko5zhMYg9DJ35UkiiaU4iR1pgqB/FbjO5FK6RN3Z+5+liw/TuDgLzD0rAYG0ww8PGvyNdZJ
lpwzxLJiBn/W2jk3c1OpgEDYpaTa9Y7kw8P54GEFhWaDeUd89am37VO9S8UuHy4c/appNnxYuoEv
lM/KvIkSrYrFoVyt5RDS89jra0Ltd0RFjP264T9eG25D/W653aBqbiTJNRZtZ7SCUSbxYXBc+b6V
2WOsZ4N9VcLi4W+X07pgogBWb1LFqMaM3S0GWgE62nkmGf66rx7SCuxM9PyPqFcNCYQM7zb19+3d
hSaNks2nJXeOIWbay8K/NzY4vSKQ6/DCHbN3KOw+D9Q5fymHGcbr9c8/xQFJWVQDEOmM9tXUGNV6
Piv0UcOyuTDGO2BPiouJSxNmwAz5SCkwwJmKUDazl1oOr8/aKVNI3prL5n/tMsVRV0uLilaGUS5g
PBxomgHnYkCpzX198CY45qrHEfuG0Gn+JpdqoATYry0PLlMieAV8lQjj8MdFxGEHh6LC00vDhUiK
yKekNxexSfQFM1KUM+cNsJgZBTYoW0EDAER7o+Jdqq4ZGRKvazX5wOrUN87Tz6jiV6ndtfpyX83H
8xSPBPBppUCuKwhdUCujswhjTEsPmcI8N+YPDZPvuEsvbNhiw2Eeug6a3pqBL1QKta25/bblLREe
Zx0Q9nWziZbDrVdCqVRb9IF8nOjH+8dSuxTLUQfO9nqnLMyaNuDDvG5lJ4QjY0w2dOCvcXaHa7mK
eXy2azQCwYKgqMkq2iVAR9qPZihMbMJyB6Z0QQ3PLEeboy/t/CXYo/PdhWz8VDTcdqwTReJFy8l8
W9b5/kJN89ecYrV2HvMH43ATzEnjySlzbaLJF6SIe9YMkVvVY2iRuKSj/Xjwj6dgLBT/XJxw2Ovd
C9ZQv4J9FPKVLVnEmHKD6EZSdVmQxyFE8lc4mVmjEfG3dAuFyyzhVGgFg5h+kN6ZI9ZVfTuUpPug
UOSDgVTVWNwFxLzsqZT00GJftgPm7D3xzOVYowEZ0qOH2EtB5ZgnU7JOjfsRD22v6jqOOPYkzkVe
XqG0yq7lagxWu3lWeymofcZJbtg16vZNJ2IXwZM3c7rtGZeHxgH92awND7O4e63fm9y1pbe0tzF3
lZ6ONoBHU+fo9kgG3Jty8LgPufROAnw1+Jz2N5zu4sfcI+5pLC85icPMcNgra9qK17BGWwOzN/9h
R4HAR+m6gc6byeSMt7+sCl4It55hGllbJ8B2mPQIRIBaSvAhsDdK9Aqam7VHVgF0EVQTlO4PoACH
1gSq3di/1ljMvUnZvkK2rfFqhhPu8DrUwepAFbZgavILib9/DzSLfzRjTcESx4P12sAjm2/TYkyq
lvfzcm091m6Wgh9v+Ql29HGIKMfPFBFkPK6sLYAGI+5fjyo8vn7Ufyl49JZ85T+B12IflVGkeuw9
k4jQPaHwRIHOB7khc/2CF9PrmGVguAp629ILSYrmIONoGSqtEVdWgF1GNc8tB4M7MpG13bHQMlex
3VYe031p0OPfoA+8bghdhadSgvlI0ofdkY9KTP35ZIK4eCKXTUku1+T7f+UwP0v857hg9eWbzAFr
pYRh4U0ZcXFUl4mrTxuaVGuyR3OMlXIBBCYSGsVBL+mbrskilAn4AwFXjvdhO7oEuYUI32MpN+2I
8tofHuLgSKdGJBpKH09WAy0OzvkLvrSExuMBvVX+pgLJsk3N1IRzFBBVQ6h7wzZGWs7FWDQT0c1G
lGyr0YbBh32ioYpNHGPXNo4H5a7AYpuG9YvA4MkCY9ImZeJrbMf0FLaUrLzzoU0Hmnl8UDM55d0H
L9IiuA9ppIHEc5TCjUa7d5n+7/daHWgrfeDTHfPzJDnw09cX9rcwnVExFpHg+GJlZ2kO53+3UFPL
ySgJc3DglIaqhX9qAJlBylLVE9rstAPaElXBCa9us7Q35xQfPcnkF1vaQjiKLxzQiTpjrVds3hhc
+b1LhbLX36JOPdGp06oilk3hR1yF7r/O6AoOFgY8BJufP/dQO5XDfrU2uztIm4mAgKdvhjd49HHb
/GnLTp46Oz559eIP2y4ZU/TTj961ozBGZtLCTKy6QvljqV11w067u84VILKAp6z93+sx44npRZFf
qcLm4KZw+5a990WfXS8QFb+MzsFnnNxGVKISF4guSpJUVDuQL9g+vnBtSuzALApTKZU4dmpiP8pY
glD0NtgCl3UgPwvxuwtuWssbwUJ+XmLtWkvBKQ6SWXltZHaKeRUMsiJMaPThvL18ZFMMrJ+Vjpmj
xSdz8ynRfGwuT0Lek//LXmMReFquWiw9L/rTyRmT9hBnJChAn89YpmeT8Mj1VPB/+GaiBx5pjgie
oF0/p7zXm+BsKHfyx+HfzKjFilw25SwqBepkjTumoSbSfPsE3DFY4UTyBbao5O1zrSqnjcZflbhw
pKSf9rFwkrxTSOw+bLU39zNuqB43oORTVc1nUNgRmOnca9YqkeLfW17i1NR1PpMrelojMb7U3J9J
VkKEge8nj332m95lBOXvR2qvjeaCRPV2L41Ubue3q5O94rXQV2N97Tl8SwU9OSpdig/oOEEA/bY+
O6JjoKVCFnd3n26ayQzqRS2Pu8Pgx8uhPNbcY1MWfU0yC7rer2duBpuRTKQpbZ1SN/6MZUV/zP51
IAW0fKYqwQIER+o+bL2SoFcocW+Pn+FA3SYh8qjUG6u5ql/gjdnnVt3M8I/m/VRkzTb01cYG01cK
pSSexTY5PhWSCdk2A7QJ2rOrFqkmv94o6AZBSVmQLUnkgPKmxZWBgeDse0xw77E5G3PT7k6lIxJ6
dK0anPE83Fc/UzCR/kJ9UdBB5lmgD61VQ6X2BN3Pd2kyapACkBc8LrLuEmfSZ1ZOPeT/QM3PGkXF
yvi2G76lqC+u04YT3HBQl8hygqMV1bNNG4rdD079N7BBxtY+hN81rtxmtavmtdoBjanVaMZTn+I7
oiaIBiflf+w31xmrzKwgF26yUqVlGxBgWZHbp/tISatN7vK95en32pyGo+QBOcAwBN8RFIgJLjbl
ioZAQ8Ms61kiP0SMQuP+eTkkZ9l4ZjDxLI0dVdXNOOdHmgk6SNeic4XoSQJ7z916keEJidm2qP/D
ocLKwagySnwF7qa7dc1m4jmfYpBmug0kWph/AIqOd5sEFcsZ+QUKaiWjvBOr+N+Ioa/psjuc8CRc
vHAOSuJIFc2xtJTz90DfMPKNzdVaqr+5r4Es23ISC6pjppgVPmIEv7rtrkmh7MunOpa23JVhfkBi
WQEuaPcKl46Ga+jpawnpcZPOXL46V1Ww1Gq7HBDsRtfgktTYOJGfx+8bty4BZ7GuklxCeU7GvPO1
483zJ+mNrg1IW80LBlgGnLPeIypz9u/B6QxF3MXucNtd3bA7miLGdw3CJwP4Q7uW6YyiLT91n9uv
K33LBIFGOGN3D1MvIXlGaZ4SPE5B+IRCwzv6yWsN/tKUcxw14nBa5iqQZ27DQETyxwTebAO7Ve1r
Vmn7OxsKUSdqYiQw7WmsNFfSC2C8sVgS2UBFD+37toIIfbZwKxSmLY7sthQ2ZeJQnUEOZzlZ+zrB
NyEKgtisfGoErCliR0KxKL9XBx+NNu2WslzbVJTbwkDrJvg1rCvJkieOJqG+EOSB3RkBcG18HHFl
LlDIcLJ2cEGpR55q2AdnWQ+E8hx89ssxseLCysCAq4IUbg7PFJ/qBuZxb9hRocnokYO3zXzDfdkN
rJ+EB2sIOfiUhLFm+aiFNmJKwoM7PbSqnyE8rYYQebr+OZ9EDvFfGNGhFslzIdxRI+oFylC5vu/M
KLfnT0iznYFxc+bAUQ4ukNX74ZoMrXFYI1AGr9+c1isIckHzIUTIz+2MtVxapvq0Vsg50WNZb5LS
TzPF4zPWQyK5Pv9l7xiWUqeO9tzc9WxpP4AzlJwNQC1wG+HSgo6g7IHtnp2a91hAh5UFr9TK/oNU
1Z+wXO24iOX1BjloIbBb0xp1tvHSqeh7LERL0FeAvFuJqWa8NOX+1oc+WsMG5ftwdZV1XBqLAGY0
1qKOAmifdzVSkQe5ZMNiqZSltV6k5DJkVXE3Sa5Ct6jjDS3SuTb1thI8S/gDwExqu+RACtq1bBnk
6aVeQkHRSdpfz2nF858wSaWUOliFt53bsL3MerogBOYG56eo89jGGWQd+3lvYwxq5M9ygTjqc3IH
zZcO5eO1kJKPIjiMaXTiFhe4JiL4vsPh16K34A0NIuXxU0cKQ+r+YwZ3qClibrr9yOcUlZz2rQlN
Rsni4dgSbgxcFSLn4lIyE+WQTtqVQZn6Kuq2PnUAkdCStdit+Kk6E2bMvlapqUvwMdUeAnfDLWJH
QG0wty7YixuhCm7820BZujxeLBXmmRDQF+98M0SG0Acj0JiVDYrOOjXR8QxFCMpINylltyJbVg45
L9KFd03AC4iCq1spuPc3xyIorMJl3+tvCqJVFH3LfhxaHmGvF+UtHcaSL0tWsPao1yBx4iyTJ6oX
csK33GaEt29MCf8EplUBz9B9ev6vX482/ndzGDACsqiIl1WBnCo0E40FY1SuE/w7xw3EkzoY8BMy
CfWvtIWNBFekzfE7K8ga4Es1nLhixe0p744LEhIXcfSVveJDngeo5ZDHryGIL3Nd2r3JGVeCL7s7
W+l2Slam1od+Qlpc+K/FuqVzt+OoOKAXvkeWGzpVE/ii324V3cOHD0QJTIu5bCcxpxXjPesIqWw9
ojzo/9CS/czESa931rUdcuqQfttX4BDItg2BxpZRK0gX0aSr5aT2e9xP2gCHalI8/z39QTHJKYSW
5SW48DoLM0MuMiBDR58ZmOnfOkvc+tJ9Pu7Q/iU55S1yn6OTguRGFqFlepdqwaXng4jBrCWVX3kw
9OiPdORXWTo4uZ9tasU3ekgJSSznXu/uPJkKNXQt4Cw5ysrRbdSQLZk/yg2KIc4czw3l8q6VUl34
t1Q0xETic6YTnDAvSmSPcmzj8sI40s0duyNf3dvhcJ4h0oK4res2LAwn4MpKnYnvruqfEGCecJWL
QUry36IAnjND2k0gB3FYjf0kuGtUg9+t7juysKLjs6+JRcmyt74xQvz6hkOkHVAj/kNZdEzL62Jf
jyAnNnuNsE+QElC8HC4T1C0UGb76e9YgY7E/iBO4p9aQ1LKL+KYBA+Bp1B5G3OPlGcSDTc6NdCYC
+9R3SKUemfeERerKMIXLV1hXbIaY5yvlmy4r6gb7C1wjCJrWmyhv+bOdh00RyVuOH+WrquaNLBoS
ZpIuGTlPi5kF7ak+Xh+RKLWUFdjPaGGVGk3jDKrmh81XY1z+T9jGQ1KeZmMSzXUQF5zyJLN5PbJF
GZiOTSr3Jy0uz7W5sd3fIdYA1Bw1QXPf7LCIkqvOgO6GZt8kqNmTx6h7f0WsvXGXPZpefzv7bLlM
zW51R6IRQhcUTp+pKQ2sciK0KDD5h0WtMvVT/jxW17XCexdwqSN+6YrcCegcr+h7fKQluTSyx//n
7VuaZpwBCeL/Vut9G6pYmQDm4k5g8vCxwecg9SCbBH91EYBoeguQt3G97V6xpi63Q93Jc662H2yM
mBH7xN0R83+CKvTj3/ydIO6Kcm91WGtAXHjcD+lL0zZHnFipBouYAbumb3ihwyfqFyI+3yEhSA+j
A2Y0vjyppG3zPLFH6y3Q5S3+mUX+78s/HmZMlCeEgeV/G3Ii/6PcBSK6ct4pB2xnfurS1EMHmMpB
2NOWvld5smhtdmQ6WMLtjq1zoJTss0vM56Vd1AWLkQowkkaTQvQm9jsdsXi/ehYhagGru1vGUn79
bPPXLPHLbWmvhmETYaDSUikPH6vqDr7TpU/okIyBz4Bky0+8z2QPKw93vMadZ6HXD/vHgnvggBKX
FG5Sidbl2qMS/XwHCmx0/ymCDbxjh2//t29li1b73FhnKQtuI+iN7eYv7WYgVrIKVOYMbZHqFMvz
nTcHf2ZtT2kmLLimxnOX4e7h1bDZHI3nTxzXmoZrQAtCAU7Vts41O7ePhHX6fHMNXeyNgBsV7nA0
ShlX9KVnIx5TCiI2INgQKrjlchjn3ReH/qBRQ3LAKj6PGsChuvkRIqY4zaRj2gkdSgPdB+JMZFcd
W6VEElKytsUuqrzxV9nPWeYCrWtiz0uzT+9cl2KrFv87CfzXCvG+oZk3ibb/Fnzxbljx/VIEj3kK
rSMECH9Pf+gjV149+ERccqm3WnWe0/uJHmNlbUHtjJa8lK9JPGcMNHngLMwWkwWxGW4Z2UnYhQTA
K5hiUiLGgjKg0OQrwbazruh8PRvIVZBGuJHsU1oii0NMLnDyHCa7JJNRtpxdagQ6zYSjIy+SvA//
BVlKmZKJ71UgHCMU9ZYHBnRn1gtrKs7MHveioMlRtcKnkvRtaBegyheWnSE7XvHd1WrlS3jQvf6U
tk6emwoncoXh6BaVYblnFRs5YNqR30tRwgtqphe970AW8lHKe/Ao0IWtQkdTlx2TmjqqZvQBjDfV
yTTvQoh3/DK/vRUMxlBOiyGZgcJ7e+9uPgfEbM3Ucg2whlTZaVaednY8n9qXWN19fDLBxyw3Ij6u
xqwdttya2XmzRWY3HlHslQlG98TmKNp2nmULSRdtUASZfUzm9qbbwns5qYDr6Ng6DnsFf1SfGWnT
LnPRczE3MvhR0EzX9adHs3bNEcK35MXHeqbsVuyWqyg34zAIeDz1v3Xq3Ri8dR1tLjKqv7BltDlD
smkiNTNWAPE0V7amjOZDi9M8GzD5k+t3aT5hpaphO/dqrFtcDWAmQf1q59JXJ2RDoz1nZ6wREkKd
aMnD/7IiiUf+g8PcHLopgIOAU7fFrRlv1yJzM5+uJDw/ILqtZhtxaZEVFNUe8QWkWjyoQYTo5ydM
vm+oFmC0TCphCzPHkM42xfnyJuBpJELXf5zanm2ttVXjshgVYTEtBSdWygDu1k1KeJyaU0TEqhQs
/5Gsgg6Wt+5YaAkHK18FSBijycWH46IPngrUimHPdk8b3dM8cY6OzjidqYc//Y7g7pZz+DwvbC8r
kGyb1wAz/BOg+qUOLiaqLqMfevhMi30qrPc9xYz0pXyeaOjyACI0JXTKAx0IlzVkF7bIMoQGm3/E
P/xtHZAcLUDFwimpYOevqLmTHIunxMmKGoy4gxFm7MqTOnkPjDvdp6jb3PG9k4TTFchSiOi8myAI
w455yC2m+zppNpWDidZq7aN8P/e5ftaEL3H/bxBjdM+vtymAVQWmVCOlKI/M1oFvHvY5jNv8152l
jKMftqHvY1Tu7T+GbjbKMoA+EhqxrfRZqix7OW88jDMIJ7/1RPLllDaONKZRf+cvdfFmn05pA60r
1SVuhLl5I1dkNavpSvcXrptXjEVCXTu+ovJv/cvRLmvRRGfBas0vEAsQiBJLa8T1uHv8M5aevqEi
xV2SyohRAuwJcNdoNQfHop1pi88G/GZRFVGpjI3fIZLigV4i2FGaH2juyqne8AjbQUwXwk5Fp/jL
2olGrA2fIM/KaPfFDXcgImKcGcQv+ZiPHYy+G9I91s5IPs9VzJaR89cjzHV3zY+GaMOdB0B21MQ2
f13Y3oEV/dH94u4s2egOMz/VYkM9mCWok4PtKDET8BQRAIvb1gcsXhnY65BzCvt4BViTSWyLZLyX
qFSkhx3TOsSKcakJiBBNWWicbq+aM6vkyvOfhW5IHfGpdg6EjVlIDSUeBHz6tRWpK0UtrXhtRGvL
jmZSgc3ZKpC54JQFXlSo9/49wNxqevDi+nmG4lT/BpG5Np95lJa8UGnOWzH7QynEULKp9Y1BCrpF
3eygo/tAwwIu8v+e6aamUb4SXJbPiN4BE7+TUIPGxzInmqXYlrn2MSfB00PdLe2LjBR1X3xcEHSH
HgI6DgtWrryxo0xmwq8OLAwIEI8LBHeqWB5dHsYdaFFctkDaQcJXOeMEqutxN6THSvmxC81NUFMI
8frDPjnKvhvTUud8mI6EHF1hcJkbsbeAiPHnxDRNtPB8Nd77m92/l0PriFNH6dzprSx+xrgwGWUm
l6oGl1HC6pB2/rEwvqDkbcdDCA+BKjudV6c3jkYpEB3cJuPhbMl95Bk6q52jLJG5UoQZdcjmzxyw
KuvL/3PyzLgP5IbiJRvYECSmjW3KIRAcrYaI2hXKhPJ65ihLy4KvoF9m67hMEMpFpG5KbaY+s7NK
yz3lDvH7blR/Tev96oXe7HA2nc/ByZoVJjUvsqR60TjwiU0M1bpLgRJnkK7sLi9qPAJzHqdPVJVQ
MuD/yKG9KjJjwh8dwbjdyHl93fIphgKmQqLOi3OqVOR9kTZlRRfaS2Cd5EDHBaaNXfi+ekOT7cBf
DQHjOibqU3NH8dpqSYulkgFLOPjzFHialzdc9S8fN4SgIjgJ4NY3myR/JDhBnr/gUlKYPcZt+pP8
M9Mz+oNpMxjDP6MfXhwx+dL4vQC68wIdcfTbM5XwPoRMPab5SQYgAIr1Gb2A00noRHdSFgXwF4k/
9LDtwH4B9olasg9jbyFf7/YMmV5c2Fn6xyaCPBtaGU0YTvwkasp8RjC1yNP0VUMnpOT+5zyjFgas
uSv+ICQAWW8ptdTBmcskurtnDBWpL9DcoPMifLZjqi5nYSdyWOHfuJVe5Lrw4H7ZxCtjXnzk33IU
tjjhcxaazd4xRRv22gedVA3XQeF5ykRIaNP0jYYRR6VZynwM2pRCzMRfWPtwVmBmUJi60ncyXhS7
BZVyzNxFSZnK3tuu+Wbx8WKfAhc/cju1FAHz7WeWPc1hO9760vt1+J7p6BjPzyaoUTpdX7MgU6k/
eWgfrQsfHWMc70VkerjnVS6WDB71/oOxyIq4ZVsGtDEf+BSAWZGP1iy5i2dSnHQVnxnQMAit3JjI
p12/0raHE9JMq9FRInp+EKVTejC5koA9BfgccfLTZ8E07wWguP6A4wWVbKqkWwN5vC5KyG+QeKUa
up8L27i824oP8Lq4kF0oWKUVttlmH9wwp9GzORpwlb8SqOfTkqqrhkrjeKP0LUoSDn8XAGZ9W8HI
ifhl9AFJFSFxYVOMXI3Y+DwMYOOSEWARCMOgovkrB+KpGjhkC9iC3OEWRSfOZuHEq8cDpnRHgK91
rPELlYb5/yRfHvgrZR4LEzus9z5Ec8zHou5coEMjZK2N/jhrxqoP5ugGH0HeGIbQt9sBp1ojUsni
WC9Q3ucpfXHNu+tLyH6k+JS1/EpbPZzaldHOdWenohrb8bpASxsfvsQxr5xFgX9n78njNiWF9OZE
iJKxWsc0q5NfIu9LwdwDiRxJUbsMEq5lZfuOn3xStHpQMot1j3xqLmdsV5QNnXzbYAA71B/ZQ8AR
cziiseULgVpmQXcYa68fyOdSgC99MTmk9xwKA/KN2Rg9v7dLq7FQBoI4ltaZL9z/w7ITO76ugARJ
4KkISQfDWi/gLJWzkS0vmfPULx1HZx6YcUb/OtcHiX8oygr2xkVKj5zYYQqhXTLLYP/ftO/8Bfx/
TioDryVFDhk35sfjU1+1yM7vq06DWmB2QqBlh3xMzMoPc8biJc7nFYe4pktdTpqe16EaG0Wl3DGQ
Ef03M4esLZO9IZQ7NRfhX0QHFCmbnTOvDzHfwKwuzuzGIZGUpWKrzAjBGmZbqytS5mO4AnWDefSZ
Bbg6uBVxTO1d+4eza58Mmr5amqF5TKTyiPpMgUHZCYpcomWmsognMSsRThSfJYuP9IAyG6fFiSBw
48SsS/hXOgygzKx7+J1Mm45XUq6M06Iub8D32kKJ6+iE4d4sRWK4ZyF8IvpvT55rTRBWS83ozVbe
bdH2xTxOQ5aC5FxkMkxdp1dli0UVaYQ6zcVEUJtpwCzcUo1Q0yOt/V6UozBmNTv+1WWrXVQo8XAr
g+7kVrljI/QFXeb2+B6nO0BsubhlRQ9w2gZXh/aqWgBu7kt/zvDFxYBGBnuGud9Vomy6K78dw+A+
nX6za3OsbvA52fJZY0fY3gAnngm+aKX3kb2FjLvuqxDj0MkOH1l1q1342eGdNKIRS2CbtdsrVswX
EBdQx0qlR5mbZpO49Z3uQZFQnQ3A9gZbVSmvLosxsLPc1YTIg6wuQ+Qv4Q4YagqpknVLZrkoTqZR
2LLsyPfxtsVXWhlgYY3p9Q7uIkAu/SZ1WuBIeKyLIwIONLk8DweK4MNAKyOHZ8NVQus/jJJxboJd
dMNK9y+Af8bTlr3ZzWwvZcxzNnjYWEJr4RFWAMW99VtpCfQmYcOD2+U/7k3mBSUbViTWUBWitW6i
xm7I2c01TgT0v7IVTAeR2eigVm2jEJyMiz5C1qbrP8cs4sEP+LZM2SLXmc9C8thcESKnNeMumvyQ
z/dUKj6E8De+p3hd4z5VhJ+WxflPVrkS1kJbR2VULXELRuL19bOtBRtDthtrToAtsMYZdHmLN5aX
bCEw/wtEJQpBF5BARYhUAa3UGVpOJvDJyh9NT3RdvxgMkpFd3vfruA2WCzx6o433VtXtKrIE6aRO
CWyXt7iRo3S23AkIgOueOwygtUMs0IY8RRXCc2TL+VDyDDFl0M/TwUBdmsV+BsxjqW7gDIKZy5wK
1w8JE78xnbhb11a+eztGzPn3qk2TwxY4gabL0SLBU+AvXComx5daSsn0S3ZtceJ7bU7DeZRKeUnF
CTOtEyQ6QoVWKMm8zjSN4wjtlGyaSqHpCc4awflL+clQSepsf5v40cV52ro6ozeUv70EGbBwdXpx
OSPo1dVQhnfBVt/aMklRJqmAzFQ6Ob0OUzQiHTA06Xp3Ki/jGsElxJvG7HTPEHkHPsroJVDu0uXM
w2wUw2lOlyRBypuAhvEMDHycmn5L5zGAXFv9TJio5/KVgAe3YHGIFmnckn/BcZES1PvFnx331KMj
ixIKBHNL2dFlF+0kDr0CLkn7YZdNsd4FCrJAXH0rA/8tctXTiJB3V/WAKyKWUjuKYhYGSjiD2UZq
WEClJEi9KpWW4S88Yn6p/Y2CXSu3XOf/NNFVqE6Uz/LTmtlNFgI9BPyG4OpoJ5UUBHyC+S0ZLXxI
5glrhZNHeKEGxpWr4cbRYZoTZsuWY8ADemyA30QNdv/vXGyODeknS50NhOlnI9kBqPA8WaGYS21u
DRgAgZQpdOahu2wORJCNod24T7jHe7g5SXhoBQXUIaMf+CbsfRe1F/h0yD0dnQfLKf+FglurMsmt
pnuzBwwgKsCkBAGt+2RHTQeTX68nfccZVu3ZviEQU4KFWazj78W6Xn8wUu9bv9YRnXHNPRFa2XIx
VjdiVeUQDkpYvuAJjt4e4kIVz3BPOm4PpvYwfy5TBkyOcymhNvKcN9tSlUMk64hYqyoGoZfWpDcB
ic9e79lYYOskhK3vx2h6BD4QOUA1nuRTjHVfsyGn8rmkyTKLZZlxy8qreny6oDeN5WWjF0jwx/T9
mgBIWXRa2YZxZ3Eb4I8cDps3LL2o9cOtIvzpxmcAZgJhXQwxKJ1r8x7ImUBlyjUXqC/srgGT+7tl
eg3ARdz+IdC6TGMurg0ROpCSx+fpmH++LJt658/2qebTl0dvJQjjclu3Wrpr8U3nT9cvIwM+otu/
UAhq+Me8FYoWR9kr6aG2nsDGbM/q39JcPzLtKdoVSY5P0P262a/dAVYZeUQBZBj2EmWzZhsN99s8
pEGVrSKA6KOsNhMQrIqYlxTDWXCBCCqmeDwHPJ7qUvcqUo6d9SyPAVebAZFuqNcTIO0mP7bK+eZP
IjFvf0OMSazyhyo+Wg/CXEP8m2A6412XOvvfbYz345bM/YsXAW91f680y/9vvpfIPYt/+L59uyEs
x+fDd4QPYK3UDbW2CtALAsZ/FoQcRDXBOHeR/8cd/az0A8H3BNr/dmae3oErI6DqsLyqfhpRE+iB
XpyuQ6Is9BM7vHtvtvMdT7hGlabP1n8fb2/zQ8mi+xtv/2UGs1uqYkY4QsN2oA/13ejNJdi/BlRr
9oIQckjCtoeXyW1HfMrTSw+BcQdLSl2FdW2iJTD75lhdRQcPHkahPh56rUHmziOnQleNQ6A6do4E
qZovbhaSapE2oBxA9igSdTVVuSYNtXX7LNr9isQ0KQEVgEHHKF+7lRzJRHLKtHJ7ECd/gpK68+1l
jtyht3OjxoQ4MSqprSRX5QoNFX8SpvtaplVRW7+SsMMjUkgje2qXyaKeOrQGi1fv93ur4T4hNPyp
Z0KMoH18PWw6OaZt794clkjrl7vow2vPIWiOx+dsGshljcIpiBdla5P02y2tlPCxweUo5CxlYJTw
drqcfrEIFNPFx4onqUIwTexxXW3TPYahMIPLtORQfRynBZ0wx/+gm03kgEEym0L9XhuDyUzOxv0B
6VSQ8QDiQFn0GbOJs6Iu0AQFNebIFHLqXn1yvOj0xpNcig+zfnP1IDLdFVfKa/5Y3YC9atOTFU9O
xYcMDPq5D8MJm40eIoDD4JO98iplkbAnP67GkIjVwA+YWWhtUB64x965MCVkqijtJ1NxBd+t1vwT
aOTZHxVvwbH0hXj0AIzP3To5G1r9XhkVYp5DNigHEQ3v11eT8agHVIN0NH6TrC8om/z6ABuy1H+0
zy6JaP7qoPjt7/uZthn9jAepKnALb1XH7l0S29vZn3Io7966J3RvYnknWshqjlyiI7DyRITGjJQT
3diT9IZToKZYf8q3qRR12Cvfoe2AkUfCUeId0fsNVt4sl91WK/o+Q8fP51uVbJjNlJnF7zANS65d
TkduPVLCqIwVV4tzf6lmjcwVlrcHUox1rIjYzBS753zCDpEyY6sVaa3gi3Zc63cgElAUah6ck9W0
nryMW0IcwuDiYMhOLkpBajbHbnyUVot7xd01XZVMn/b4FBEQIIFkytWY1cEUNlz+L6at6prS92Wb
jNevxOxiE1x9yRft2KaPi8QjzjxbhZFi0LqLpKQzb9ibKl9aB8DrXOO8B0FPAHgXIjm8DOJn3gCE
9R05n7ubJYCYzgW2i0rVowibgbGwM/u28TlAOtNBBXHvy10gmCHlR4CunCcBypUaSbEJCvgrpFgO
tfevyo66Zbiy42ytSCtrGw1bkKFAYEjtNMuDJ3XsEKu6ZH9jncNgqzSfHlSN7WgBtxrUWve1R1K/
2EsERuYfR+AjD27df0RePHh6EW2/3eOAr6ZgxgLNQKJgeg8PbmPvT1/LfbA4O49X6Ru1dZ52Fbjn
VhTPO8aeHZnSig93iZMuWm6/EZjoC8K2m7MPSyJ3tnLy15v7TyM9/sN/5J7xx5WKeHRKUEuu4yQj
cM7m+n2+BRXyCSY37cNk421yRB9sK6MUltLkWRQzUGE7g7/y0ofjoIsvy1y1YJh3Fenp1WO/dU3P
CMdwmjUEA14l6XtPWN79GfY9C+ygifGJTXvuy+2w5L5e/eBPs8WjeY9WMkuYBEb7mcosscJDuedq
8t/mY1FqLqjoRa56KTCo9KfwcMrAjAqkrYUH2aEcTcGtiG8igv/Lg0S4MovqDBLq1J2aGGeAbCuo
39PDFEIaLa7onZ+ADJUjQVfhan1D333ehHfgXkRvARonruviADmv/gPJ+ltr+bi2Asu9j8nu+2FA
M5yuzAtuNDWcHlbxcoGSOchLFY7m3jaurCpxc17cM5WaJeuE4y6KZrxHZix1bqpqUmEsQaZi+5jv
vXPoG07Ygaub1L7Wg/lV2gsplOsZ9xKSIdA7bPR38BAnE7J4z+xI/VIW2IpgjXmlN9zSgpg+jFpj
VbgnZ/b47xP7DJeaK701cLmznqz2t+eBH6k/l9m7G005CevkRg/6ee4aGaX3QLrxD9WV6XgGkAeD
xKy85c55PjP2Jeir+ZCVEq9c/BbSnugGrAQ/f+mRghkPQXhPKfezX44ZPo5EKFPiLskfRS63w/4U
NguGqZQ7cev5XrDWgFNUKTxoOM3hJHohFic7J2dJaXkrxIoSvrI6Y8neCGSLTNBXMojpw0h3UEsy
inbSbYVcnR4tGbxotPfnW/O+9ppcgFbbnadmujOgZRVHw0aWnjNKITduJ22V7ACVWAhs3LowBGvQ
UoCyY8wVvx93R8oNH6x2SnTLFawLyhYQpW6p/3FADo2dO63n0CAlUbG8VtffbL2yoRQFsU0cXJLz
vyeREkfQYBYEpnlyacOX4cmhemGlsyhtN8arEjNKKpUZZ6c0k1MY+RgFTz2k5g8cnJhOhJKyh9V8
6ap5ewqjf4BhPeenm2OJo1/RFwO5lIO+dIoAfmesmw0b5fkdsb3gfaeQ+8KmJDYJ4gJiczYqdpRI
DRoQlO+P7WIreuJCro5RCT4DEefZRwdThHL+VNugg21O0fArhohH0wpGuW8gG8D9/Wm7sZvRa0Bg
eK1MyqX2UaTTSeIXWxKdqTHCiu7NS1Uo1SWfaIVe8cJkpjgsaTSEYi0SO8KpjizhZIBaatgokRmI
ZvQOJjiFACXMMsE135Nd3ORtTLyauhCe//GKDtr4nu04L+8Wdn7oYHrcf+/cJ/JrL/5C/jPzczA5
tXCc0wnueEOfdCjfgfEduCe23GEqiv26c/nk6KzPhyOwKayIGNEqrswkWxbF2myj/KX9ZMkTHSVp
td217htHoXaLVLkML8Dxsiap8+Mv6HumerPiWkZkxw3kSuU7+ziren2kfE4OsNnHrQd2HmXsS5xz
mErcfCRgUravEqw0nZAg9uYMxQDR3S4g7X+vOG+PG/uvshXRbckdZef1WR9EOCstzuAlRxgOsITD
ueNCuuHbFDZ8exv7w6jpNHcl4RylGgpcj9VnzCbFD80cNWlOfPgRIVnPkqovlUT00zmpiGu5rOPl
TLZDkDm8tikPwP/gGj1v74r7O3mp0WODd8AnUKwzhOVY2kn372/YC5Q0W/FktgV+KHHGfJOVm58b
fzbwLYCruBnKSjL73XvhWZwDbFm9sqPHA3ft24lEyAMl1iDTVNSfRSuqPICIZ2LV/HVbxhbbVwIz
HPp2TTj9CFa4baMGnOWFHu66MXdSPxAUALsVfMC7R86wHSFqdud2gau27xAgiM6uBYZhJFKHqiZM
fHkTdMt1TrwIpFNK1LlBqIbkXEReGakh/D3943niIVis2hpQfCISZ6n2VnY5IE7zstwnxk2sqEkF
ckqKJjZJ8SwkO45ehkwXgo1HSGb3jSwyxTratb+4FPo5ROR2cGJ5J0If5bAUhENpd0By95os4Nax
mzepOtknAKQ3ZwoOcZ6bcHLMh7fs292t/Xm8U+yIZSN7QJ5HSw6zM3BBv3fap1cIHyah3/ly6DZt
HioaglP0YJsOVqAfq94FMidYHWyA3kw+dbuW3NZqxx1jkLg3eZKJ5+KxpFrkOcmeGijFcRobBuzm
pk/1FtE4Q+eyQTPGn0DZrc07bluwT3edpYM+9UvXWED+hypMQ57jB63nW8RmeXSWPgTrcjDjdl60
ImbxrzMssmuAnmPRqkBROJPsFDb6ZOKnzKacbArFDcv1E0xIBFlSldWsWvYEMj9oIyZbgIRr+OKM
Ri6G3jPPunqJ+FEh7MkQoBE+kTeHQJlchZn7VounXkjyIVANTLiD8pksGDAM8u+wiVZjPV297ei9
fmpQjzHXuYnD0qyJ1cHikCFgBvrVFXfEsh82LB6iM2XWDr/skScZBHp5RL58NYC9Vi9uELFQLYuH
53WDFo1xY0C2NgJsOJIVpqQ9/BW2U37rf7tM/DbmjveaOTH87lSxZtAugLva+S1Mlc+s4zaMKnvn
T+jzg35X4eS4AWbGyQ2ueJXINCJXoanmOaIBtbdI1s3C/9IFviYHfarXcvKOR16g0iLjbkJscWaU
J2ztFPyTkIZRsZuEaV6AFkPHr4nXBrvJXTp5eA18i1Ea/WrJWqpDvbeRXZu6Yggnrya3pXFlLe0U
nIFBjv2Ix3zpoycJ6j34lw+QcmNRFm1ZfBdocfEg6juqV3YmDu8HlCHO2Dy50hM/GkGtnGMRtoLK
8R1MPgZr/NU1m9gOjUaL2lxy/RQTWqMO6gIUXuuhashaCtXlD/V1THUJ+ho0IC2cxwCKHxdFOm/J
uXnXcUuGBQAbDWutCRunA2ge0TuTtxlfCa46FNprwRuOMdunS5RAbKX6A1DnjhYKxbgybrOmmuSu
JQZV0Wj0/FwqIjNq4JKIZH3mV7M4dWoJBzdV9D7B3A8Uk/InEXbfB0kJ+kc0Z9m6WFN6lenSGKba
OldYcGuY1/G4nbPjI6x2iefUQrYh01ZonwOujKoV/pynOIXyZbGaBApVPwft9SqJKv7g8UYwP4sw
Zc8M/07CvDmAIoQS7np660SG7pE01Lt6BuoP0aFaVheW5xPSBPtr+tYfBkO9V6vUNkiCdGW58O7p
p24IKIOt6ehfl0yRQjerkmYFAbI38IJEd48ILa8CVyAwTKsubLze1kVWTcMW3I30T7TcwXTeAkwa
1YwD9yQnqYXo534240SkYMZaH9WFp/2l1yx/rj4dQCrvUbgfagpL2ZCDMWci6CX3+hL6IkSRSiND
YnKya79y7VmeoiEbnbIYBF6jjOxoB/4eAMkAdGrHwWMHplKRZWE8nPp9+Zr7AVs41zm8lw0ZCHP+
s+ZkmtKteA6mcVOJ9MsUMkZ6hmjlzweAmyp7a4IbrlFF4WxmWrFY4/xPZzV2ZuZQEkm8AUtwaNXU
GuxYw3AukObrjVWRRdZCzQ+rqmxIXvpwHOd639jnJrBcTUUYH8ksQ7MsDTmUYIlqfxSYbF1HbpVM
g4W5aGAS4YZsRoQ2BovgE58HIIoCsWyiAlN9BgBvHsbO+VuwmhyMWUTH2vyL7VG/OwU5Azs0O9Qy
ht/LY5MzI7lFqScrfdVj8QvToMY/lOKeerYnM77dRF0gHPf0+pIswsKAaMZA5+KpyPh09UPf1pTK
m2IfKxwc2OmBhQ5Z1pHhVFVAqwXm2on9Ntnh+G6rBWAQDRBKfwILjCAykxUcSGAq2AKVgGvG5NbC
ccawjkkT1kt4b8nzgR/SFApa5WiPJnGTbdsFR7DUdNdIF+U5CXFUmNM3CtcwJeGxbEtRpfiQtrRr
+QxXTOHB9l4cwopjNNajiGrCPV7WKcV/cWPcvPj1ycrQTf3135FdrvYMccPzjHtBg/Hpf8ZX3iqZ
9ZUqGiLvOYCEqMlTNFF/o9gQOChumKnK1WLjFDtRm4V/RdlXr65h+IcKJeyJEYJS8C+F2izchBZd
e9pJ75pSDpWD117/C51+XJYvEWx9I3ccwYAETjAv2lqqRRKUrHdjIAz2T514m3gNHn9UA+A4/8tc
AB3CBSlv9z2kM5cgl6Ivvf+H+HUxzkcUvF9YBQzlmclTTsO25CPH4MQgg5bOrDMZfsw569LIHnnm
gE27rMkJ38WmRANiKQojfIpdkpVwEWQSySHLdSyoYfKfsbcQbNPCYyhzyMvYgZEXSl7GB7lNAGRY
a9WTyE4YZCf7RxHqgwUGGZ618kq/xx9C32ef79MtUGIXb0ldZb8QTBFYZate5Gqt2soISTZIwCdQ
NWpnpfujgnTpw152brskHKngG8w1Uhbyad61ar27POkcEXU09NuSjAYiMsrxOpRYmvLP2VUCx0M1
H6UCLMXAxrVLs5EoG62tHRDjQp42udM70Bp+8Gd66iyFZ/lBynf2syWTk/p456AjGmU6QTovq0Un
1fl1vjLIVIvdAnKw7/v1e6ClMueYDM3tjNvpJYaaB+bwExyi7Mpr8OC4+ZaiJjdQg+ec1fHywCeR
tBvQ8Apy/9GCIdMIYt3qKTzsGU3+G/GjZlaC5nMHiKLneCoKsU7AhbY16lmtl3vJgAEgpiekC5ZO
8AyJ47s4wCnyVPjik4egdqpVjDsKNWzktthQYMoaJr+3XC2SEZUFE24MeWrs4EcH5G7pVf+3Tv+i
ZbG4Tfa1IBgo06PT0liaQIObDc05DmMQt+2LA33nILV2YRJTnUYQnpjA8SWUClSzxrj60C31viI2
lENrExz+gIATkgD8ixRHJy7wBqlocjFO1eKrHBawq/QO3f+jQQhnN6KMqmhRgcKRo9hB+4iM1pkf
PBpu14WzXMiTsNFwwQysA8wFguBj2ZiIa77fTgqXl6wc/mA20OS8/fhyb7KAPA++/VyvvYYZcEWk
AROdQpG2MkoBs2cURrifLEmRM26IjFpXHd7bO+g7qbZDuQ0rwKQer7YqAbWGI7AALYuV6QoLEF4n
gTC0gqfRrxkaxJXojEsPCggCnHj2ka7hAlshR00aVunImNnoBou5OTE+5Sv2wUILdguY9UcB/fsm
XR3OU/o0kwz5A7oMDA8bM/4zny7Hqw1k3ZBFeIKQCIdkopob+J0TJypPlGlgD8iZi+zFcCgtQGmX
TkVp2ex8q+o6yesFIR4nloGmOMzNED9JbCfTbo7mWmV+VWdPq797y6k9PypTnfZuNB/aWgkwAyz+
Hzb1XsaP0sl3tVpDcS/Q2tHcvM7IUaMglCNwPnlSwLuOi7q99m4g1yF4u4RNOwZcotJ1aY0OQb1E
7pTg1ygUow557CblrZrJox8LF/4Smj663/kPJOY7sHzBaTF7DH2T28TC51pVgipKN6dIO9rRuxHR
u35FNo+UOe8HfX9JhzeQ53k0vH7fBw3Hpc0GLC7GYxN28Bl/ktY4v/oFOrwKBu/FDBWSyTVE3YxQ
6kKUSO3UvKzqbnh7TxJ5bZ/nRZvdnr89W+HCalX6lVAPEwsplKEzuBNvA0r7vT56GVlfdv545xkJ
EomYoKGAxzsaPGHwe/+BmgZVz1JJ7UafmAm3VtF754LTFsIbaeTz2u6s/tDVi5MgFhIIgFnbDWjd
eY4Ew6f2GKCwRjsOYwEJZ5OPavqkK1IdzK/poni4ho/sukUpKIUgIUgCYV1AIOHwrFhct1UpQ3gI
tjBxgH3w7uma86tOH563rpmTm/Ktnuq4dS+0hWA6gTa5i86Tb6hcyCSvE5Yg0r7FTL5YRF5L7wqj
adwEpQx1KIqSt8dbiVmB/FS2HvW5g6Fa+pq1mwH/dJeJDFJXsHoBwSEZ+7eO0GhiMD6yVQs+VXba
6DLeaCmP0T/uDQsb4QkgMMoBSeSQzSYUOwIKVixSGxrds+EUIt2RX4SFXJAGDzicw+IlH8gu9tA0
3UQRcMAp1Zf8EbVCyRhtqumbdOnHoNNFdHyBreFzEoBXjErSv2oDasNVBG5ZonW2clMaTN6sOGiA
itZA205d/jXOeJ4Mnv+Sk3TBKLWOueGctgKa3rspz4XhnmPqzTaMZXq6vHyyC15sB7Na/hEQ2h0P
AL6FYGiFXemqNkgrAjruPjkhraeJjfH6PKGxHlde+2RQLlRymqeQpQ1HA5/ZHSkXbV6r1Vc9Z6nH
HAhEqTuG7pcMdiMjKj+Pdl5EFZ4kiN6OXCY0y+o/ysqAq44HQQLIpf1OBmuQBSXYvshQnfJZ4Tmj
YcynWgcr0OiFqaLyHN1UWC4j3IZ2pQhZxgVvdxHwP8s0EhfpA2C1SRO5qCR0Kj+qpyKSJtodlloq
MmtktsTXYrKNLeZKbpDooyhH9dMJ3uajtag/LgnBNFUa5QH0yiG3xNBkdYHvtDqfviKphoEXPUn1
y3edgq9He75MtcSxvMjSX0lKQ8mtRIoRcrgy1XHWAWyb4BGgWfT86rwheQrWlhWz6EL8ritsuUhY
BrBJfWEdBo0heSqmpUVkGC7puSWsLSAsHxwvTF48OR7FNAIqG21zXXrOxMAx4Hh1NMnZ6xlQy1Os
BJa7wCpNhQB61AWd+TxdTtPCdzXh3G+okm4P9zQ05dwiI0613h4cuGLVAN6f/V+qNva2co8WiAFN
955fY4E3PSthxHo6AV93Iu91LXGPwUnzWInlg4dmYSYYZ3uXdXa5MNccE7jnN9Hxgt9jZE+PYoAs
YVOBbRLCcPyTJiGeKN8rR5w/eHSvNW5IX9fD6LWiRQXJQ/DwCSR3Q49UNFnhi07GPe5mWBQbwtlf
rW9sQtgTOKN/uix+Y20d67jEHiLfn3iC5/53gtbXjyjd7/e7XfENrzPtI17vvs9ff8E+DztZooN5
G1l96xwOLibsm9nvOIrhAsf8DxBT2Q3EinITZIogZh4a+8IyndBRVm4tToY4Arhnkj+7KcAumazL
hhdc6FfOP1M/MAoNA32LHieql6gCvnEx5fiQyoZnT1H7cp39XncmJsbdgoPOMLE5saUdu3TeH0kj
Aex7ziaCH6SoL8lUe/o46MCB6Alh5807NMBmg1pWOHW26Hayww5xQ0n8jTTYNlUQQS+vlGN8YHug
VMpNdioUAVyRxkqDxpddiXuKl2oS/u+UTvKW4FfkBgrUKDoqdhnDGOZbsGQ6X0Lm4RPpRRQf8kzb
xTJOCiuCdkRLo3FGNeaXNhoxiwPuiFomi1Dt9Z+9PE/ZdKYBLs0DNBYFgRALLHp4MQMxKMGFLeoB
7kjTlAKUoqa8TBKscgbdZ+E9auZl6fgQJmxchPZHt0XpbEi2e8SmPbUUKcChKqgySpM1SV2zPGdk
tKgOaFuXbMBQ1hM+WkS8ZZ9L7b/DHVEhu59P39Ieq0xDiTfiWd0HNHMvq56VldGWChX5pZeB0xi1
rUcDfhlHCi59xOZ3Ax+A5Evm25GUJQ+yYxIPag/NoJX3oJxCCzmIF0dr7n+o8RiS4LhKJOl4cFBn
xlWdjB9rL1v76TGjawj7H2dcs3/pFTXfvSdBVLJTi5/YqpHmYluZHV1qtaS3wNNkB2ONmlAIGvSQ
gWPhUZL/d34vP8z4ckVcvtATOakPXnJwVOldg5XcpODugFi8lWdGihko35eQrgMKBTndd7SzHTnx
duGbfQ4GZC44mqWZ2HEQqxQUL7SPtm4hYvBeCpOKOgvxKealo7/A829eQjrxsumpBhZEz7KqGp/K
JpRtk0n2X/XVtSLKBPk8EU0UHm57EEe5sP/38oFYaF0/8b/yLiCPEkeSg8kL+1igG54L0WOfeoz+
mMK1OQjrAptwODk8RxY4bS5gFwLJxDnZnNKyIVzf9z9YZc9qp6IpEyD4X/V/7OabTwUwLa23HboK
pW/np+GF3nWIEGzxUzURv0BtnhuPMuV5nKQfIaNaqwboFdIFFPls7lbT8ZU1ftnAYiGWvUvZsvN2
eDXusFwF7Skv6BWNzO6nh9tp74yVFF2zY+uOAxDtuAMn7ZelBxScM2U4p1lsx6qqBTT5Grjaswjp
4BGU62jXTVccd92LiP28zrJYGdKK4900bHNjnZ97R1n9rmLk5GRzGjQ2YGd5xbWOiC2MRG2wGZKv
E2F2nZiwHotb+6kgGpzcMIgVrZLYO2Zx3QCBw3PG3WtUPACcQz9F48nFkbwFLtUguhJmwdwfwFxJ
QEE5iGgxUVdmMyQidj+DzImxpspLQSAziESP3k9pXh88dcfWCC3cNGqKUPeQgKVoHjfIjRfxXWNm
BRgKQYKVwAw6pmkYIjK+6GMVntPsCUbs3lCynastxYdau0HQQ/pMbds8qrfFVwwnTXGh1G5xCt7r
dcr7rqBdHONw0ZaJ8KWf09TSlSG8pxInVtIXcl/JJdTDouSWBShefxNVhdlNgejFY7YgVFHV26VO
QmG/NY7ePMYcYjU2w7IN45dOxInZl1TIjEQ6zwF/TpL1S6hbt2htxWbziNu+gcblRwa7O2kGCMRH
3wkrC59i4DpOiB0tmg17VnL6qOILyPmUc4+Ec6bXwW3V3HOv+oyxzqSZPpgtF3mPqsiR/Hzo2zNS
AsXI+W+w3od9CPbK7dvFJ4YiJJ0sjIfhko2IjPzY9lj/5XfRbxkemRJffZWG1cY2ASl4OR3X3l8Y
9TH5gwc5I7MSnlgFi8T8Os9NDElmwHhIzMgfgpPQ3FeOr7fMO61r8HfrEVCce841zYMK12Aburmd
MTbNFxhqRhZl+WWIa/ks878ZermDhR8X4SMYJOF2bvh3oMxKLvW5T+yqcVkRdAC1SmtQHB+VYpjv
h20GWeIrVkNYu1HqiAnMNwJ4sijZPrQSDR3dwpS8OhENO/DJ1nIKILsT74llWGuDE4CVJgcTVKlc
y5z8RIvHIE0FiW5T0diuZkBgqHdtg5+xoV3q9oOAhLfhkAIUjk1C7ZKYamvQMtfEYL0mSbVDfGvM
TP7uBBzVluz1eicT2Crqcb1whAU7vrOSKSEKFAXmzN9UwlaVtmSdQe1SPZJWwSemlMX4qqgvzWe4
llUjXhavcqRQ9IrNHvZK+yh8/oOT1RgbVOt3oor9Zpe5KDybweRLHKIoN9HzFn9Pqdj5V2LWym/8
0td2QVwxKnKXiHzZIGwFJA4CS51sECA4FQcicmLuxHzStU5AF/MoLesUkZmpz74xjr5vzn9Fv6uX
nbqSEYwXjKsOGFXMuWDCH+LDiWbHfdcsrzdSoxAmMD8Un7VnQZtFBK/raQd6thFk6UsW6IypvCkf
Bu/O+nLJ0yecpERXvR9+POmgH9vDCAGajmmwDk15OAfbhQ+sKCKf4tVjjQgev9TkCO8j8KpxlHgV
satT5E3EcvAzLqbvd16sCbZWEGojifceQDLfz/wj9+uWvzM6V4LcrVxwK1iQCb72j9nh5YvF3tpJ
0mpDPGwaWcu+bBQNnKAARQEoYlbjdaAWwxGQxB3ohwAJJzDca5kqvvQxgcQEEMMfBO5deIy/qUAK
3Asc6RN8N4LJvveysANRj5oD47aK1ix3KCaSr+F47a6Dibykn+vKK4ugql03yjB5aiJjuSJvDqII
RcS7Mkz29x7CyY1oRDo72ducaSY6S+5HTBLXZdjbDvLFXXKRel9nhvRQygOlJrN/SMZya+pm2uEA
E6OTaDcOzm8Qzvcb4KTMxvw+C28Jmxu2cycRYnVLqUGy9KRJ3qqGLiXjMgL3Bp7AtOa4p0g1i+zS
Ef+GgoC1WvdoRvhMIah2aGNDqIxZLxvUQRJ2xUDfyv5hVtm606n6zWdp7ezciUXilMsYPtDy9HGT
VFuczRJx1BRt/wuj0rKeeNMKRir3pbdyCdBP9mo7O7fUCO6DB3mE9c48n/5Bs1WQuRyf5Lt4VA2P
kv21cErDNZXpEgZutJHn/E7QiQJnizq0k2fEt65YCU12rjYQlo3UVhfgiE2e3Vi5Vu8y65VolIJt
O4obKILg3OyNqgZIYo+FZ6/tAwjXLU02s6IDRPd/M8UqcC/jam4LAIuHqMbP1A2H9IusA+DyxeDe
qEiBRcBXYoyEOvMiwFKOdGeUEh38wjS5nBRo/jCbQ2D6wMsgjPbhHGBcWBjb27+NGtf2raglL9LJ
Khz+H2U6xg9QBOAOJOTwhmbPZud4ufGvpaxwKoe/arLeJrcB3cF9kF21zVZiSldlV5253lKlf9fR
e9cr1Sn9DcUhjb697V3F4PIpc05s8WNbcVjPOJt7WolrOVWIN0i5CdNjbioMhq2zN/YHB41wkr8+
FZIIRUtJCzH9uHbFtKuZssGihhT+JB3zpSnyF/L8o5m9uWNgR/qg6JbHeO0xUCWTBF1PTh9fRxXQ
geX+6xH8YOOUQO7kQzj3BR2Qxi1L4tekbzCl5MEcy0WabHMsvXHqc1A+/pvZQNhj0jGXzCdjpU4v
DdkgKj5/AqdeIcTul25IlrwMYm96TR93rFdeSDcV73xpr4E89N7rv8KaFUnSrU3VZ6fJgm9TxfJD
XB1jdlnpUz1eX88yKwPra3p39oAxnHwRJXZjQPnpmzcZfkB/fk3sC52MrsQDuGSNdxA6QQNY2dvb
GYjTRfgopnOwllHcrWD6VCgT9tZpRs5ZCqX3N/go+UjU24JH6bcJvHt1qc7+YCwR3RYwV8Mp5gQR
Z0P110uc69o6PkrsOUnkgeocnIlPv/noM5y93z+MDaavzZmtqWhbL/bI+nRDbjzeLeeJ2ZXwS3tZ
QDe4lIa/wa8X7Xz9QwaWCpVtc6h7ApLReTngCVb9J/q33ED5MaskxyjOulZTypIH48h7CJB9LQqp
THTsqcQKydDqAqTBJSlrLHGpuBvuqt38lFnCMUeR8Lq0xVifhqltaWVdpDQUlihH4KJEBZgykReU
NGDiebbiKf0JXil4ogPxsl/GowpkjB9jOijbPpGJ5pyaWgDJ9EvzapLEwFkUIoI7NQqx9DvEGIyH
5zMBImVK0WSuhlgLmh/H+f1gKO+XyvPrQYUz6OSRzErovjZOTvKYWONREuZzwYE7LfOfAcQHDTGi
v7NBHarReAicrfDo6f4/2Fb0zQR2lb67m5o7qVHE6b/u7oxgbysWhof4eEuSkeDnmSLUxGsZsqn/
bE+tFitSLySvBWwW0FZL6YmJ5KJmANN3kcYi51Eaome7ekt3eh5e4qQtUBbJWsG5Qg1xpfYOepfT
G1sUQlgtr+J5SB7GT1nN+VuPFYvn2vaPu9WfgaQy98dpVcrzyi+XZmivKY8+7egMDv6CkvKE/ZVS
YSmkosy1YdOcrWV9gXRzwCmwcKsRSOa4tzw3qTVEU5yEHR6gnrIKcrtzfFosDXfhAXbwz4Zku0W7
RF0WOavntKK5Iij7rtx0wvj45TPhi4Oe+5HlmLflubEBi7Le4ric10WJvSFtPUMUeuO+oYnTUNSI
Slo0EHfvwWtDyZQIiHdjBCH0P0X0W//uR++niq2naZAngFCJ0HIeIHH6VXvssdQNoWlBgLxvwntU
Rt5pwQH/HqHqomzhLW+0rz61K3WqKMKC7qz+wdEOk7WMwfiyGA+yDDh53PahxEQThCknpN8U6C4a
DwIT6cD8MOU/q7ysplsJfbaouB0LrVpxvkrNBaMyk0RdfFqjoWZ4GgKSq0HLkOuJHz0U73v06g7b
M9+Fm4VgFbv2OUW2tbFroRx7s0bNRjXpiOpz3Ni9DAna3pPwVDbqAclO7ExGg52jHSaPFzr92U6o
HWEcizI6+gx7egpMZfNUR8Y0q7Fp+LxpJ7k3cG+AVdjI0KFjV3yDf7lQsWxHOm6ESz2h0v4r8kde
mHXV58n0L+dBNLKkhmE4/1ZDsvSRdj+Kpn7sCWu37ZOawe82SX3a8zeht3d2yJ4vcyeSo1h9/EWA
gecWTmWXPe9o4SImm86qtS3g9OO9n70TeZXAIu3cB5vVeUmMpT7DeFzpqCjlRzZAWwTtd3gjsRlU
gcS7pGF9hIeoFT5IsI6n9tGfyK2Zg2xB2ZbtXjkS3Yo+aubeZSDlMKdiw3FAShYgnyMac5BlJ/HS
24ARA0eaJs3f0sJ7ReEq68xAinD69xqctxrvy+ccXkDLimB5VDy4egsJtBbQSsPH/PDqJvYDOwmV
DqKdObyTf2fe8BwwEDm3t68x/CsJeDd9eI74V+MV/kliPQIfFZfifWsQ1NPzT2aXuCmZU1RXkPct
xxmTRRrwtnJ/Xam6V92pYxrkrhBx4cpNpGp4qjy9GxPE87EVuAg/yvHlQOCyNJp+X8oUKpTOvl2W
sywZxrW+LjJ5Y2tGEinVvF1TjFRhBSZA3HWcDvq7vIpw85RMrQIsUF552taHaMqeLh78FbuR8Typ
pI+GcW4f38TKlz7i9hsgwXEPILvb/kXHJDzlFSJ3yPHgO6TE9toknxfKA0bl7VjTsjLShXb/OITN
PrCxCxkIZsINS2pHsQhxTycqTTG+kMHB63KI1KnKnW2jjc3Ip2v7kOgYKasVCYLL2fZJy+vamhCA
eQ3HTN8QZicl+uIiqqUk1+MmmAAif5TD0rbYvY4XyPL32S8Em0cwdFXnD7BVIFihSOKZRqX1SsN6
qDAs/N0FY45T6TXafC+cMtBeTPMBzaRO2/Bo1YmJwYe5ptCmi2ZGM6g7mQ6SFlJSQs5Fe5DryRVc
QeWbmPkuv3ksaS8rAFPaZ9DmR6YuF8Vm36536bPOcEOt0mfvtJmLtSNtbj+9FqssJTQQp/K4Zkyf
j17QD6D/YCIalH6Q3inCE6X0eJb2msfiU2holvhoB3AHt9gtl/EUbQdzt45LeBFUh2kVE2p07YJh
0ZEzxZGjBLPpWU/YGqoVgfsZSwusgLcW4wrBjz1WDyaBaU5S1Ju0ogCy8ijURKijzkttqXL0rjJm
nW8BM7gDO8HcP3/0NgnS5yt/zfiL7THwh+R0K09lUa7wrygz8Z2JHbUbdXSqjyWphCO3pO+GUyJ7
rFXZsDS+vXTOTPtlC+mC5NkbFQaz2STBmWsMmAKfLBvMrmQ7aJ7UE4Zk18XMKM4JtNOD6rBeB8MA
zwaY12XXh2lrdZIUhVwHTR4AtwwdwfuSRobp9ezSWHQID+jX0OG1KRJloDNGZjEGUPBvqvlqP5mV
UogXl6fN44cN2Z/IhU5nYLhdHsugIhCcVzzRybRjvvTWn97JV5veQvNemTQ2vaXA7MqQZuK+d6Ii
cxaCq0BHOKIAinphuIvax1B0eayoFeoXhU8PaASAAU4h4pHr6I1WvY9LmXbHzlXTkjLhNqQX40Fk
MIGcQ7oxciXrVVgFxB8sRizQCO4Ej/Pz7WCL/m2JGS5yPSL2+vNOjtq/saMlbYSXuwyozi7jnwcF
WOmu1EjEKoF5/OZyQnf7EM/dwE86IQ68+tdIMB+QsU4F1MfgBEHbnhY/wtbAk/q8FNMTqYqwBqMv
bg9qV7LGmOjoH7RE1Zk3MorpeQuKmPTUFJGghGnm4jN4kSS6a/JIVzhm4j3gpGMOQIUcZUL9aqxl
CW3J4gUW+6Tbe6xMEkP831RBV+GXIC7ONOg7gUS3ahdmC0zBHnkaM5aEJDXTiNmVWzypO6ANTMK/
7/6HBG6rnYIpmrV26N1hV3GN3dVABmcZBO67FO06oXMPAoB00umgCTQxRA/gTlzOdkjuV64OV40u
6WgCnolxSZW1T4C2St0Fvc5WLyLc+o9ujZvf/0tMfG1wrNEUb26XjSgDPqe5jO9rZMV+aU2WCEkv
3Rn4qsP6d6sN51rQKX31r6OUyQa0ccFso1S8mCnHXCCKi3ppAOAUcz/7gJRuzcZ0bLXYbeiFlBGc
+VfuWPCEeSLk23kGcgdJKeZQNHp/xrrwzO0yOK/UVkek+H5kn3rVm3iKr8MBpnQYjONfE5HrqFmW
nFh+VaTr3lXWO7SZj57oRSlTS4Ji+vIK8BX9Krh9KYGhqWqIuj6Xu2XMdZat6MCH0siCnvlabxMS
82FfsVUtHNRomQWq1xwP942b7xbm6bK1swOetY0Z1lnsWrF6mn6tqfCVVHRFR6EHVsavCIbuzrDo
WG7gFxHTyP55piDWg9MIw3sMqomsFSF33woqwBiwu0id4X0uDylv9oX/pLNgeVbn7864GvHkhFDH
XB84XuiJjMkArp7rsoL7UYhGIEitYQneVCLGh9XhQmqU3RROs8lg72wkcxYpyVUYlh0q7sEXmSLL
F7wx7kPZ/VQr5mKLcWzxE/KPBDImdJumrg+0rVhlIIf71yolPWN2G/m7SqpvHpsSkM0wAb+ON3QG
YqTd780j4YqeVP7cU35ZHSJ1EKJYyBdUBaoBwrAASSgWGwHlWKZT1RNEMWKzo5pR0c+1LMyzq1Gv
bpqO8Xv2TLarQ8SPIMxEE5x92xsYFJYwrWsKSr76rYrUDYqs4E1RIZFDJiD37RC9Nd4zclsT948e
hVdE8ZX7d87qL/7Zrz4XQ3C/t1LUvySt6jD/utbyBIeumiydgfI5HJ9JJYes8Rj8WyS2eQtr6+IV
nt0fkXti7gbLRzZqSSIiZBefGETfM9F2SzE38DX5vdk+17rbrOYbg0Tp8zjzSYUNKKGzaImePeo2
+ConQnIkJVj/E7+dlEcUU6d9hsUj17aaXt2FEnhp+AQyDBn0xcI/eqUtagOQmTXpKPVRJ+WmIYLa
+4oJmA/NoBnTzTMNcMiBEd47bFMu2kf75+/q6csQyFbQqUVb5yC/kskQR978HPTI6e4FC7lOJHeT
ElD6STzMRSW4uFYfD68LfTqpd7pvZBtkULuFPfQOUfZxq/wJqxdxDZaiEnF3O8RKUkpfhFGhZWyi
8p1Z1D+a98ebDImxoMf1nnXw/HxKKIWRlTqwzuYGwPf1bUlQaDeQ5ePjjZpZ4JdgLWIczLH/hJhT
Q6i3d6JLWDm79kQ4HdTjlIuVhd9LQTUgiZ9eiS8zsgihpeQaqLJjSLOMi7E8tD+kS3py+HVN2SY+
IV+95TpL49C3BRjFlHZVCqJAL3n01lLyeb1dwNYpasGL55Qofp5BDLIJSGfLWQ8fgcolMxVNPifl
qWspZEP1C4sfm6fFN78xBtjxuJE9KpGtzWVT5hpc82bTliYpS+rd5lPyKEpF92BKUulhhUID34MN
m3RoWp4ERpGDLO4I/ZCjUkVVFpkOU1RFoita5cIFxc4EMQRXVh0JLEHkq6aZ4CgOgp22jdHP1iqg
BkzMYw1QcHTzeG6sOY7EEmQFoyfpWLQE3KzjnvheoOfBLRmA1B8bROx0pB7LVdkwOODnrgV85X9+
LZOMoSeqdct3E5+OlFOVi+o7iWhRfadrNILWYFo5lKQes3CXbqWd2O6JbaF/11uuLJ5YfMR6s2RT
Re8e3oAr3ChH+0Ffrsc6t2WZhxzUiXh7CUlIu9h57N9P1AtyYXd0StAYz9C8P0Ekyx0TsAlOFDhG
XBufMpM5C3BwXulZT6VkxATAKRkQG23MOEKTdmbS/kzu8qc1EUKU0XK4sxOguoqJcDT8CGKnMaw/
2smMq8aUnGxRhScqafyIjfbinUiX+NJOy/T46DTEgAcc5yvhBSprPvSAjCz0EKdnXuDGinJOIPYI
ejZ8Y7jcZixlqKUPC6kVIwO1nZWXwo7Mt0oR8Yqcu8N9RPZsD7wyoqdsIbFcJ4rU1jagux5UOruv
77DjLtOPrW+EQ3jdmqvEbDtSJzypw7e0ax7qGnAhSiL4th04BLr2Um6bx7bqu2iM1u8I8gJtCEzO
GWgoQ6uXaaf4XtFtxtLY4yNS4ve0r3Ep2kmgrHi+50xCXLknPdk5P56IrpCD8UUuP8dIH2wilyaH
/lOZBJ6y5qPKzbhPx+Xu1fmGO9d2Xcg3yRqePlcRAgC2quFNGcWA4bMvWrYA4VTeNZPuYzPOrICw
B9g/tfNFz6EyhmUTp7nR7IMffR0/5GxzuHlNLCbWzlw3dvgeqZk1jterqfwvMz4bit+U6C/tQ+4e
zMwNKrRWbAHArUAda5pw6L9CCClhxToUfRWIdZa+SQC7yAQG3wDeUTbcJUBedvXmGJR2m2toLHdm
iyWSUs8m8pviU4pekDayRupBmAg8wFWxJydJMlrMQJPmFL4rwS5YbTIBxSd9XF78zy7VYT5xpr9s
pnOLTawFMX5J/3UZL/RAoQmqN4/0mhHkHUXh/3aCMCZ37WqzFxq0GxPGCuXXHVRRXpZs+thSAd/M
BSqQWXgsHvtcKVvzoDucXpb7C6Fxl9O91KlSn8hHkq7xJP1cu/1yJp/yGKZBd9WNx184ZiCvpf7B
MBSaOu/eI/Is1j/uFy7+5pWRbY7zGxs3hxj7+aKWT3iLFnm+Q8AtOFd/oli3MD/6RLrRjCvsGlLW
apHXvmRd7jO5RqL70qStH1787/Kt6uEwBKbYraHzaoT/OOUxJnBRjdM1E4rlHUypvVkjyDoyAB0r
i95454kTai7fufd4BVAfSZps+HslEwBWL60h6nU1O/YOV66ypIyB+P5Uo1B2dCVa9yYXvFZgu93W
cTOcN05IkibirMenzvfWhD95/hWnqTEs3Ope7tQv+gfac50BS0AE/aLQkSWG088dunlZhwU+Ahuj
h7mIXNS3rurzH38R7opXHzQz+lr06x1LyRkyZYdgLcYBnlc2Ofmatt7hBPYsw5zCJx6UsJDHPqf2
kDXy9DWJzVsisZ2UplObkG+OVvf21A047dpyrDW8Rz7ss5yfeGN6bxAm8v5VcLbu/iLCmt7UMdsQ
a2RlHGG57QhYqYaLzHV2kFE1RyEc2+WQfttDOhUclXmCRrkZluiLVT+g/rojvD3cL4rvQm1x5fra
6dTPJ8PRStnfNu2s4en/m8YaocS+PbSyklF51Baw5F0CY7npxVMJByrRv7z3yqKBrZFlIe9DAIvm
45mVZNMS8cCIPx/x2LLfp+ILhI9EUB9B4+CZJSyFUdQTgdAOUo1UWnL8TyonmaYT9yWhiK/cAR5h
y6sZjQTbIXUkUv0FQKE1B7TruC11gcl5SBD7CotHvFjyJYGQRggvBhHv8VRCUkuS00BEBacDNWWO
6U46HcS7V99JLUdl/lBI4vZb9Cpd5nQdEeAMh5xMWMFEY3QdMsQPYkmJzmHnLnuipd/imVjHwrBN
Co4Jy9QQ0GaxJozJEGqwjS5vqvDqefd9FqON5AZUwDT+Sen78BNk7aaRSP/IrbCDyTK9HDkzrRL4
yn9WBJVAa3aLqgeUSIrVXUutFRggFzP2fqmE3Li5zUrG3CwcxNPyrbYjq4/+eRIG8TdDsr468nMl
T9UJiLWzG7gA8nSi1aD2aAav/PmL/DplDWFFJSYB1LkFCelWPTNMcnsAdr0Kd71C401UuftrZkQE
GCglbnLRRr+7Zz8a5ezl4hFCYLKJ0j5iPymZlngiAUMe8Q9kBmnlaio/TviGJ5Jm+Zrh5QupJQMB
zeunV255uC10vZiXu1ag31W3TxAwGryZsYfCm0qPE5GkeQwn+NBz+HH1op9+gipQhuTrKYA/0QiM
sKGdAkHRJAfq+SeAUy1bctYCTDXsNQZNqAkWVmIfuGErzy0kporfkL1/JG2GE/3i/5ei7COuW0pi
TpQILPcyw/+QqUs8R4obzcAqq8Z+c/ObNey5ZcAeG2rn8lvsXMehyH/JD7+4jgb1Y/hrX/t2R+VC
OvQPFkZfJKnIiiPxzSQQiDVg9986KQvKzEGsg29lZEsuVDmEu5xMmzRS6CJEwAb15xeFxBCYH1M+
u0s02+VlcoopK1o9CU4fgi+gafOYrq3j/Ew5ThmD+ZpkToGDZkd/Ci7jSRKJT1+8DGOKtak2tpSV
0nUyBqzf1+bfYTDh8Eeyu7kjUUNEtfO0MwTelk8KCfcW3tBhmgpEjND5SM+PDhFp2IjbHkkmoEDl
mUNeawXtQMHwyDvijy5Hlji65ki3YKnUvXs1Mvc8W14XIiUQpcE17uNkN6RQc4BcJB+o+++ODy4r
rczqDWMgVOZ8WIgPdYgxYksLN2IV0KJmNaDpxcWfFCbiI1sG/ukf5IQ83L95jMnFlono08d2UgDL
2gtb0WaV9C/jvAOMkGI/sgLPwYQV3FNxF7SNlpLQq/soOWIK6lxCrZw42MpLSxkcTopCLJLRqdwB
BI8mvjzLefft8QqqsYhj5FACMPBRl8hhZkw5pOLPbFhl3gBtDXlCdQRPgUDsYnTvXOMel14xr3bj
HoTe09cGPZggCQZnntUruFd+3IfVsoJf/ThOLFRAYIZQBCnFq/u4t/WqR3HiiknS4/8/ncz58rnB
9HLDdFxDIw7/9htzikadYBSswlOrqDNLiW16PFul6EvbD8rTaxMOhAslLfw7A4lehGlIsZ3hdxSP
IybQTKQLg2ARkhn7518Q5xAEDqENxkcGlSi2Uff8RunvchSXv+1nqyd3b6fXDuKYEbvDuQ5vK7wf
PuZscq5ELF2xtA18CKOz/axx1uZdlMU/j//Lc6UH1NKlQyYwHE8zkuCokoSsMu5TVagHvp+PwwO2
WBpfsS9kYLHSZnB62FsZn7rsWw1NHL4ar4io76AqNGNr2u+OisMsHfvoEXsv1vrNmXg5qmxKRbKa
tFq2QatWzkKXxiposnj45UANnvbSWc4XzPO7gCK7FPvo8PGFoR8jHvHZBks2rtQlsmBEzx+qw8/w
8UeWOWw+ToOVpJg+8lJMseXZ6f04vLtyxHRWD43d4Ga6Dub0hjUrxixYhk29el9jYy1zKMsFnHG+
QxkoAxqLrTCN0FdjBr6XJEoB/X4lDk1KgnKFKoLHQV6PLUYT9KWvqaiufFJw7hzmQVs7e9cCjkyA
y0txn6OLhaRHrwsrKT2VmagrYdK9pfnjdkVwW1fZc8GxTfnPu3Ep2Cl4OkaB1hN6nlRX/kxSp7E3
mdlyrrRwAtZfQaFqAK/+MUPKR/Twqr5YLVNqUMC7a7KAwIauX74wc+o7L334RmJFDj7TEcHuchvx
e+K52cfVcbS35KJAs43MOJ32FC97aZd+If48E4QspjE7Pbl/YnRbdIYJof1ZcY4f7Egwbvi/rP23
UZvLjtGD2O6FiTxcyBf8tm+c4YQC0fzmky0atjxlnpWqlBA7PrxvZZA6guf7BU96X7AyW8SfD3rp
oYd6Q2PAbzpBnDTuuKwUdiAO889ohuiqc+uROuBwSA2ecf+ND0u+lKgoKtj/uxoOTn1MzzzikVKC
2HNrH8MfF+Ua359gXDsDDOT8wZr+z4DMccdbMneQ6o3PI0lFqdbOg1hk3vXLttBQZJzT10qUmGs/
lmekrnPfkqJw2bZZXmsuzHVaKUQkm2yHVH4Su6CARBIvnL8F0LOnMqNwPENR1P66v33bS/neeEJV
FRyFp0qG9g2HeNIxgSQqSoxgeXrzrTxJeFX0zfmutWLQ8QlIF9rd8QFDLeYj4MyEe8JP2908Ib2v
s3mQRNzTxBFeCzqoLJDADOkkdt+rV+mjqVdlQSR5oTRVhprDUWO/OU+rSicAhJJCYxTXi7fJCIhY
JrNyv1sZyca8eZzHFtEw3mUzOesanVnzw10dtWalPdMA4eoWuPFwh2d4Qvs6ND60PBaZquYijkdm
9WItzmDr4ghnv8ldpbIeN4uX3sOYSW8cwtpbJHxvmugmWHabs5Xp5VHDyKOSFbQCr5YfOx4RUBFA
ibv2XyMfCEnWuiZlw+cRr37OeFfitXGWsr3a296KtK6rekYrMH8kLqS4McKYKeJ7BlMlWrFYEAG4
a8wxjgi1QTcFr2wFgKZyecTpVsXk/BjZsbasiY7XnNvvHDOv6IZfLE43lbIPkzb0z7DKtYD+drxw
cqpL093HmQ9UXL1whpH2lgU7hN4IIvRUYDAMlZWfEAMTPWw/KhyRCMsiMumvg0HrXd0jKkdPJjdJ
tG1vqo3e4KYhKQEn+Wc1VeVkPP2D+FC2FII6uzVuQuBEXgNUKcMLCnKddwYntbGQHJUh0+4JEY4w
Z2mH6XdbH0aOWRv2XhrZqj65iMGW4MRzty4Sq0Ac9vWZVK3prW9moNXL2gRFbSxS2XDkng64aPvB
dC628r6bAS2WLdwg7wHGdMjU3AldLKXglTCbrMLyJEUPI8KIYqsxkwClpcR/IvQc6uOekkxDEDW4
CzoVpLyDjmycMbhbowvfrH10hLx3s1MrFhZPfDWQoNPG66TdSHaDeVMSxSyw3s0UgD1OfbL+EGbI
rV0zrO2KUatvjhY9gJLvEO8/Uyf0QDgbcqkDBJQDaGJym/PrAdPgMflVPkYtq5OX97AVSLI9Cc6d
Il4ZU2f6jboHL3PssX5FAwx5ni4E1hux1P3YWO0BtvayVvxqbq43oKGAOlSoD8TKjfUly322I4pB
2oWCQ0DBxwORA2hptZgNhdf6YQQk968yVZLdDKF+N774I0W1ZuLV2Fraize2gXrcrNAXVTmDlj7h
Lr/byn4HOqgaUzHX8mlX2lU6xhmlH030WxCtGe78FWJOYO3/1bE07srcb21NeVj9e6ALgnhWD7QW
g/6imDWDJh5sO8r2M9aSBHPiMbFvMnrBpkzQ2oZkK9cGMwtMflcgN3dBYSkdleM855CTINmVMh+Q
Voiem0/6hYjCBdiHIGrxaOpCUjrAwgxHPyAQgvLHMKI+vjbRdaIIE0cpecqMgXzS8dXBLqzArPrQ
i3G6R2LvHY2pbWbpA6i746sDXConIQCbZ6P1F5M4gGD2YaK9wA0zgDFLLJHhPGvJbtpXMyz8ENfm
He8FUU9V4tGk2byJWyZ4sVlWZtZaVsbPORleEtR0/0dcgfYDsP8Mi46LjB2YG1pi8m8/MvNUoWpQ
rBQFF4t9zL6wp3sqLPDEL0ZObaDAtjdd8Ub+6ekCWdF0CFVtQiWHMclVVUwH7YS+wA2idZ6aulST
HSG5vR57p/YCxPgXXOQoeFoESdhTT18crmEYSF86VLN90j+Rvu755hcdKjtwS6ps5lQ5/6RGgyRl
0/sp1qBHl/E+HLin56+iPK9E6ZSXLaZdwXNIMB4oMUIdYHIkBiTTmM07jcS8zPUvtUzhIe2apGO0
UpANJrUfdLo04ubwgWKazSBpilYpgoSIJPV7BnXbX/aqyI5Hg+aSc2YtK/5FmD2hYiFOlAZStq2O
z2gJbCOhay9bJRHr4MALPLd4kdU+RcCfTuOAwxrR/XPU+m+EoOWznQp3iE0A/pxM3P6EJkkiAJs2
frMcXxy3Swu4k4a0ocKnjR8Ahn05KUDd+Tm9NXZfuvVqVebxDsO3TuIIfpAuJC8AYG/iVySvte9G
nUo2/q/ygjV7/AZ8i4TpTLUfqlBt8FXDMQFlSoCWzedupgo+NMVmzZYCl8USqwxuXvaswbbYpUxs
/qDNxHhqo3bHFVvReKxrhBgKIpNKWH+UQ0D631rYEEwuI+yYh80OMgJk39sZq8DmNYF08LTaOkMB
k/huNFVFDTNLFbZ/kE8GqMfL6NpCq6MIGtlFc2M840NFqtsW0+n1KeQYQm6MLnGavNoM8gxUtftv
S3q74OYQCqagJvSwcq/kFOnD+4/lOU7OBrORxI0ltyQzcqgPnYmmk3lDfP8K7ejZZRh1z+uB93NA
C5iNbnfTCtmFfZ4/v4ls0qJBKqlc39T/IjKhO3P+SCSNLUkJE/7Tagk07m9H2EBJcnWBPSP1+wXt
VJ+taT46Jrrj/gq3oe2Wz+4YPTuCGflNgQ1Z04+++VqZk43AgyZkzbPvfi3N4vnx9+DtJslMthYr
E/DowlLDJPWIsWs2NOOt+KBRcv0j8iNI6NOAybhA8Ua1pO6aHuylGKCr3v3xqYENO81nIGCe1fCK
g5C1cNIcEsX1dWYPi3W2ZUcGFHrDf6r5+g/ElEG7DFyEEd6rUqMr0bjS1PMpNa5G2isStEWgaMLv
A8ZWve1+Q3FllYSsF/pd4f9/TYXJSi3FtX80ObSOn9/T53x/gu03u2RAm9nX0wX5N4O6N7xV80Zc
ZZqer3OHro6WFAV1FIGXaeRyfOdLcxkdDufctx3c9B9hZtFjPoT3sarDg3/qv/AmfzKQb5ewwu2Q
7k+BpBuVDbPlpOMT2s+W7NVbD93NIB8jlvXq4QPTr8qAqi2RGq1Z1+pO/ooox2JDJTvcPtNGv2hz
TTe0e/ait3f5v3t4a1SL/8uVVjITlx1ecyCoHx1a0c3PzEVaVQ13551XwXk09qvJRSZC3Oqpox2S
wNywErDGigYBnco0ZjRb4WcO8NgqokXskp5HkMn1cuJMWPqvxNXKBNKnk+qljfQO2br3Y2CGLmn3
53daTWYC3MZLXzi/U04P55iRl1TTwOv0hiGSA7AbTXcS5gZ8NMdtHrBOaGJMgF7BFmyNZMYRep28
5X8SBCVqH0x+d1BWZw4lxoY3xCknBsS1tbBX0MIe46eP4wYvNxm4+mwwJ0P1V5rdTwVOUJgb4U5P
61stT2RoOeZGfQLYaWk0VVy/p9RQaabeK0GbiKpYFlnKmXwAtePNraZjfUzTxvRhMVxDTNB0ERkc
w1vzGK1Qt2767BS/prZExl2QhD0o4Sz1uGMoi8bEhn2ozqx/xz6lsvTAiokSJjlKQve22CKV176b
FvmfkPEdcUEEXoLO10D4SCT7Wxx3iOHgPEf/kTT2cl0gfd7qxITAkIWaSE8CKWIX7aVVVhvATReZ
wIKUe0KinPS256oJyG6tzRvitl5mcxAs4Iw9kV0mD8J7y12da+dXhl59zzawvsvLd14VHB0V87qG
7n60T1SFSCahdq4LPSuuc2X8mDkvSWO2dBH0ndV/RsSdGFHNvnEAU9NAXWoGc2iaEIww8Q1IHID9
EAYrLhALCVB2AccoZsg0xqgn/A58ufJmek0uyAWB0dfXTU2/bcTraGKJV8ftZmjDTl61Z7kdZ1ut
O18kXr4pMR8e/HNr9Fpob21izM9DBnq4G0wXVWB2QRQ4PGdKrcp4f8GUuKX4kcz4fY4QNKLMBMYa
PwLAlH3Zvb7yI8z0FQbu2ksxE1m0JVA041b12dIf7CCQ25DMnuxjwEJgGDE+7y1RDN2/GhDTpshd
cl7waW5ryXqxFexdMc57eTgDn0QxoyVRb3LC0IffWoO0G6WX9m/zqfUy7rH4lLQiK7qFZu+/1Edp
V6eBV7PrG7/emxKNoCTlJfFhXWsl1rubo5g6/paXbExiXeYP30+SPkNhddpdcQ9jrQhi7VpEp8Ez
Og/AIIkA5t2MsbVMRqhGkp4N/g5VYJEyr1yQwGBxaTBZR4Cs4dOlrCwA0XYV7Z6Ohs/5kqg0REbr
7JKdPrjU6GlzZb6EttvnHVi7RwASZjtBocCbksy/XEY7HDiaUVh071HP8EYLUNiokHd5MxqXp6s4
c4Ts7FWvVDwtAiy6KUnKTHX/UPNcNnQV+MxYajXPBsOhaYODWmyxNATY0jcid0w2Oo1JvbgRxElD
mrzJ6E8UjRDwZlN63SoUKXlgb1wB5fMi6pPLYxdqKQmzDOOM4HMYS9WFn/bRJoOH/mVIX2zIZkaK
wKXSObWwHUe9fxVb+HFbglfff57ZQ+8U0eJY+ItjxJOUlJ9aJbuhqOs3cy4Q1KJJn0BYN/QM/v7D
BjbJZ3filkDKwZ44z11pwuVXnh5eLy7z4DKrL4RqwecFCqsAHlyrm2qxA5oIKrx0gQzm479voROx
EjsVFqLAz5o7ps8FlnyL+8ZjhTWyxMcEFxblg2WlgblRtRk1Xm/PeqotUaXgOH83cLnxBmalam8O
M0yv16FdJT97GhTNO8o72AmPfo0mGOY/K3w2s3Kt/De4tj3TrZ+V1FeZMobGS4nZANos8YigT+eJ
IPWemE+ew5nmwOTazux64Dt825oXSr8+dFLLspiuZ0hSCb0SNFgFcJqbaZiRwHluNTyz/2eduCod
3vHOeQsfCCNVk6LPbSJp9AkfCwAdOOeY9CreBmSHDyLalZWw8xEof9IH4JWnZWPYjGtHelvQiUsS
oUiQ+GwtIKmLc+yZL+KlHNUwmk0cZ3eSVL4S13LEajCjr+4bdW8SI/RtasL71jUey4noVHF9qHvv
9HxF6Id7jElb2Lta4H+qEgtAJX58mydFKLdZr/Rja5ttvqLrRE5uwGCTpOs2rZnmtmNKxRsWI+N+
gNW8NLFH6nKmC6EUwJi2VFua81moc8bvKJfBoFDqBJP2tLgjqsb8uFo1WLvWaPGoYpmRAvJhWvKs
+JUqGy6jUhIlP28pxxP38oFzYv+6lN/Hxqq7JGTDXeQnx5kfGvAF+PCayE0jHzffIz2QB2dLALZC
DfR+Pink9TVaVq1SS97vYIUa0RctRDS5UY4+VlcRFCKoMqWNS//VbeLHE1woXcsi8poj0wgrIFkg
8YfVmkndnZOrOgDZTamug30USqSJHGrdbQYjfXwKTro12xL65/QZ3fMJYWeUb+XnIAjm21ZcrTdM
hL0hNrt4j29b4SlUQ4azMdbqkgSUoJgNpqMZys14KK3fib72srm9H4n2y64x9nN4xqgqcxsaOApq
uTh7Veb6f1OMgeGARjsL9wiJw8qrdPu8WzFdlwA2YCuFn4UVxqcblAKa4sYKJZ/iHtSmcPd+ve5l
Vln6Lx7GsE/eLW8D0uebYLXiGLzarWUmzjch4mNmxxRXLhDoctHHVOjE3Gnv2XfZHHXcL5C1hx2x
5ttgojpHqTzFHEFAmvpN+o7NUP6XSuba9l3j8fj0GFhk1faqy1waZ5b6QaRJMdtVph2YywxGyrXI
5p9S5+XNI9MotZsCr8P7bLFZoPACKfgaZxwjFKWqDr6mOZUXUx3XNCOmZf47MSBZN+oxhkvl7uer
jwzAzbkpxswFL3vV0juFdB4HqLMFH0Ybk2PF+W2712FG4svDow1X+G2actsBksV2ZvbKSUFSEuJg
F89L7a75xVuKZAlb9pXroB0f64d7sfx1Jsv9vpZG58f7U3MMf5tJT2W0Iib1SjXcqvdKElNiANfY
5bqAvWEKA/p2qUOxtcQpNrWTTXOCinDx8avN8mBMAnYYhwuY5sok7TWuI8q3MBcCBIEdqXsdI1pl
SNaI5GnWfsVh+QYpfbzRDPfei0uhuxvLWLflOvR8Fq/6CcAg4lAqEtbuc/4cRpb1dhugGblPN0j6
gMKFMEQLHUkUYK5Bygepyss6TuWJ7cVaAP7YWPRvVti4Vy/6bBUVatGMWuViVwZitV/HZjA2lMqY
k03omxAxPsZGH6NnPD/HdvElr3egJr2P52dlnsPk3g/yYwMsMCgCTnFCe7LoIcWgKymx8Pcx6f+X
4XQAKdOXEsVkEGj64DiNWX2amoMs5LFggCJnzMET1gPM4qOymq7tP5Rv+Oxj1qpxjVnXlud62RKQ
XMs0tEKoKiBK/J1k4ML+m8xiWurh+0mYDKjS7yvVsT7wZevfbcLYpClZfuA+NHrj7qgK2UPon2/3
+EEDT4U3UwzXy/qFI3NWUSwMwMxLmLpn3ctKIXZeSxsL+w6+vjk9HV6zrsWKPZ0WgoDPsCakOR5U
aKa1+7oHuXyYCUQgMQK18NUSg8DjdNwpb7jphAa/VFAiozHq0wyr3M2/4UNMkchd3Chnxv9w02vH
NQ9EWArLoHNqZ1r7weToyh+TRf8MyQwIB+nx0+l2NavfN3AFfkjk04KOdMdTSzxTy8Dc+ef23mrG
o3m0G0d4Jr5bRPd4Lnb9qsbtukAm4fWYjSdh2qEzY00L66mv802PCrkmhUcNw0yrNJ996skuuZjY
B1pJtma3rJFPVL/GZjBii4sffrPaKZmCEpJq7cvyxcwgc8Wd1zUghRTJVSZIj6diNgPz+q7ER0UA
vk5Nk5ymEIL+J063QjVip9LYpKTwVqfsaGlRO/23Bbo43dlBfCHxslPDmtXhXyROnwfjXz9PudOU
qmT5UAoP62Ct5/MuOY8tH3QIDTrYRa6Wd/3zreDZaio+auVof27RMW10DD6P2bPjF5MkBMX2kI+x
P1k57Vffb08nt+T5frwv0UhM+7BcV8CS6ZN4zeAvsCfUmUGmONYyEO9nGRqH6exO/SG3hzw5pPvf
F/knKfVAeGAl8YkN2tOF5+SKdeCRYarEC+9EgpXwrSaI73t7qM91Rx8Dt47PqAjoYgaOB9PHOv9q
2xCHHS83Y6w5mt0DX2s4NL8IVUIkua/VSveJSIt4B7GH/xfPFihlOuTxeWy6P/eGHLM6Y18ExSEM
0weiXMEOp3BsgVLITxhPjEn+dRxegzhU1igiNPAyUP6b/FlCH94I89LPRg3/kQNhx07woYeMuS0F
6x2cy0T/HLo4iky4oT9rZ6CMmJO5BVZaeuJOtTB+OkJ3ZUqcxOLgKPbu9nqnuvIvAYbsCwElO7qM
VbnS5TDPT//rYKBqgj/P4dnJxdkfiJ4nDSQTsjT6C0J5UEYyfyRr2GTQM25yqnQLPvMUZV82gE0P
6WE+XL31EasipQ1Z9DCWYOTRFEHuXhk56TT2wADgk7nzq2Aoz3HE/BAnWNRm+NHBTWDN7TtbNS8C
nImKw5x9p1dcAqdazkhf9S09ZxLK+EVP10S8Rqkon6yFtKi3TwWOD4kuedz7OfDoJ1BvHCt0Tpnx
N+DezSbvJSrVRPHwaMiURj9kf67uh12fH7y1tZU+N2NN13XAQ+u7p0LfG/grqoen30Gn10bkc0I8
XRGKKzBI//nG9wBuo0g5FRwLI0PRapItxZnN9XxwiaIZoIbnFxWlPROUkL5vYkKcsLgHf7K3Z8MX
+iHPGdGLjzfL1gfPvYs75K58E0eETgKXr4iRCxSUDK6Gu10TDh8I7tuwruO7zPIVdQgCQVaLw25P
738Qr/h9p28FlM8cCz8Mu8mWddX1kobejnIzO+m47VuSMZAoKNC+wDTF325sTMvHct4nq4FSh7XI
jC3YeawzkPE/8NHSAhje78JNUeQ+lEyrZfd7zxG8kxIr7jd+oaVAJHE21RNvVne0Q/K7CKODxqxZ
M4YOvNhPxFwGPUGjlIH219Mq3ukQ8p62StdSacWPPe0xCgrNzNrdt/ZKP1LbQlgwGqcG1oAxag0H
GkObqvy8L6GM0ecCRlom+uYo9yrZtJZD7GjU02ZCvSPWVg1PD5POzByyOx/hksNJyK1MKbPr28sO
NKO+JSTRKuOWvFZbcaxv197NAP2F2hwFxTgPDolEvLOFuA/bEh3vua80g7hBYDUdJae2o1xyq+3X
WUDVvQPHL9E8I3NAdiLUGei+Z0am8C5Pjoywx5eXnAfZ767/2YMUmy3c24anU7QdueeCoqPa1a6G
37ZzmeK87mluQhHivmgcNJJxzesPjDME6jojKHTdRq7pcD0tEbBM1rfowOzyfkCxMl9z988sD8WV
JTy58fMELRQ3QS08md4mmD+vns4PV/bUWyrL5/6/e7EAPOqBskPNW3kKRq3feoO3yXWG7aA8KIRV
iQgMDjNawQA4WXV/P3vcfTZFzumutlr06Dll+1+uZTFmunHzuzQhFQcZ7SOQUD1KlZfg2g8/zQvK
0XMXoJFem+4q/uK14N5nf9oORFuzaVIN2+GcrZXGwXe/dCMsWLx2cNuIofCet42i3WLGyfo+LLYb
xthvBX9rDNkBAy4MfnUCzk4DQS0NhTjd7WsXW+Va+owseQkoNVCq+pASgYTQHGHEFCCqRsvIZVAF
x5OXF/zIVAEjkm3OG4jQ5SFlU2b7FPyg8bDRXFoHUp+znwxjYKjXA9JZTnD5TCtKQkqVyvaLl6VF
DCbO2cogSYUMvpm0aJj0D1fB1g3PAcYC8UO5+uVb5X6LD5VYdHW/r292If1BbQtVnFzJSD70OU+i
PearRol9sBsB44h855e2xD7fGL7vhjOP/sa7tVCwn8zHWo4chWma027y2pEdg/O0jyyXYdWAIVys
RYf6sX7cBZHbj8BAzTdmnAF3QBjduyQM3atvY67WDz+hycBC6jsu9qtQtnyv2g0HxlyO0X9U3THd
ZCh+03X7sLYImaNyy8DYgXyBfnRLfurc+vg9kPIvC/GUqSw2fETxKDF830/g7tK4SYbHeHnzC1Kt
UppTIiC5XB27QspviwgXX273VpWhOMc2NbcYhHXHeyQpTIiFHFk3TG031p56W4MsMBYvBCtGA/EF
WePFkEL9sEWTMPIUxKsV3l7pMrGunNOlUJmykWLjTcotvPoRI9jrswFSyVNJ+1+w4xe8h7V/qOhr
f4kbEWe0QWJCjBghH+HcQqalgmwbVbfUkwpqhzhODvFhcRGAGJOccBNwn94ltbw/Rj+sjo0G3OEl
PDe4gmRcxNpIVVJ6NfjoUfXcLpeAYS4r1qe3DpoocGs9rsBbXRjeA9o761J1Z5jU+kpK5zoqckCf
d/5VZxcIMWrXgLJ13Ew7EaUqYUdwZX7SDQsTw6NGs0Ihpv+SlFklXxra+5iThvPZjn4CCnEWoxiC
GRxi/EzsMj603fwAeMQG2aL1U4+ZCyk2qUvBEL1wOJDYF8iL69DM5PuI/Eh5Za/RGWau8kNOAn/w
9ZDy0CPmLOT7Q8pKlD5rnNmReE5kW4uHqCW4xfrSZpUMW73RfYaCx8aEvmU2UN0AT0aiv2dgkPxt
5WwNmSTpwoL9LCp+QdiKuK5Wn7iczUfBEgWiywkAYBcwjhZjCw259ej/3kv3Tm0yR/mVthuQcj/k
423Q8HgsI49Rlmpxa3sZUqOEuh88cVeFl5qiGQgyl+CgfcCd1vgaoWW+lRdsoVqvzQpBvGK4DiK8
5bx2ikz6vF/0taFaAXEANHd3udev/rNR/hmDpHxAmY15sIu2WhlYLh3e6jhXE9Xr0jmvpGswVjSh
68hl3u5VP5wGdQmFHWMWvMwbfyhxqjz7GayHhbAAij+oMzg0Jpdl62/povlhLku185p7i2LGfFE4
0jUqZLiVW60NBDQDfDerJkO9+XQGzGdr9m7bNgnJrdVuBRQzt8lMm/M8gtv/O+EUQ1jwY7JPuIBi
ZVglw85DCICxhzbR2Z7uqL3L+/yoLUJs1WZkTbyTlMZZEn76b6PugAd4v9XbcKpS0Z4CpnLyfS2E
4Ob8J9xwmCh/kj1AvhUSKc3qTUjtrEu3XVvc5gcxmjYUaN0+OUvkNDjgx7pqjvaLVIaw7zCZaOvF
OyWsa2m3zI5rXxlB41lV0chasYpyrBSjbVLEsVnQfX3y0mieG+bpcNeKO7skJCaE1p9fB8RaEUx8
GV24KHhqudg9WYWG8GahISdRhvg6mixRvW7MSkV4HizjxlnLdCMaCUten8E98CKJCKQoeno/Mzmi
IilAMkd1ZFcUcuRKHlMrLpUCszhMyt5KcNjOSYzbCW/t5f8blkKi+66aZHDXLrdPsMCCmdxnqxmR
HD764UJ4Nr0Yk9BYDF3pX8QWeoDGyqp9/0kRk4Q19hkv78525vaAwKWtLrmJl98pXh23SYXm6ooN
V6cHTuD3b4UbM7fNYJO+e7bi0wSywOYzk8WUonaoOHvIwMVX5fvHHC3+a3YRzgSWQBpF+BqaTvPL
PJVe5z/zWoxTPcAcRhvXIYQmQXegjv8C/mHFnMkR5UEH6kpkbTxk2kT8li3OGEARMe/eawBxjwyL
ej9yfsFrWoMYyOy8IIp0gXMyVTD7CLEVkfhVAPSULKsVF8auLrXvf8XL2DB1YPuKUutJtWmbgApF
579aqyt8AEYbDpo+p9l0p0cQKG+W1kvXr5u21ewq5LyGYFksu2NzuhRKmkexsJDo+MaDqRqhdd2U
7bsXKuiKLPzEZPeYaHH07y3rDzkRfHdgeKj+tY5UlGKKrAL8AK3JKpU8DsqyqMLN5ysFGrUmPCdA
NR+6l5iGZ8CmAEsEeJapoyDEMiTSnKkg7uZxQ+s1on19MHj7JIx8BQvhA/WWA8kTbkJCVK01zmL6
lK41ZiZzQjy6cpPVZzA8hurQHDZ6Od9nZE/o84bgsM7g+rV1q5GWah9x4soimjRV8ZCP6SviZw7Z
rZfo4lV+/eLPEy34KKD1vmaYgS8pqgLOl8RQGINn3xBd5vz8GfyZpXPs7uQ81jd8HkobJeBbKPBC
IgRm/mR7VH6TOTsmk/EGS8qhPaZpl008+/bUONK4CjOje4r0kVoraTzfhrKfegDco5EKI6Qzggk4
z60ypUUnjYkaG+Vhm/sRdabKZ4wtG7NaqU+C/damFHnXEc01Ocn+wObY2jQ0nNkrx4AnuXeXRxup
QS19oFfknDaI9oKUwo3EGsCkYEtQA3Zt3l8HAHLaLOqOBprtmsEC8hFVZDLTDsiymrqBoWnUzqZq
QabwjVQ7lL6r5zLckGtkAg0AGDNTn0Ffk57c14llqI6lRGzrg7VQRCeksn5S4xEzmAY8hDp36ul5
I1xgGDzhViyQSXg+dXCIlejuiFKEYSE9RjxKTc9aw9NwMK6XQ2jqdz+Ss6zWJ8+TN8MwAOlljWD8
+SlG+K1h9FDeuF2O1jkfmeVKMJ/3Yx+1Y2S4Eh1ij9VAnXgLlVQRJ5//yX3H93S3stG1ovPSv5l/
TvXuHndqqA4KmnXGtVkQWzxdD3pR0uVatjOqwq6VYXJY91npcP2plWbNagM/hXQ2xLQNO0njTiM8
m9huyhWuVnvfU0Be+XxKDkwVw35+8jSF5EpdJq6cBL8rF2QYPKc7cuyfsmXVL6M+Spcpnll7ir97
Ky+JxABruKelgn1LyBKofbEYoi1Z0LKyWmVbrANmSPTL6Wo0KsKcZbKnDHEksZlT8EvWapY6jZNs
d9vneL0cjWVDUYy5KT18JT4iPuQD1D+W+X7P6vSkxuslPGqEy73xu1+BCTZ/dMBIwYqmiWcM6Uxl
iMkqeI262b661AqXLvt1zk8yc5kQ7Zh9OD3u3Wkf4SIjyZ/AEd9cujKw6HiUWyqhswCHzXSHQ+6h
cMHn2RNKRyRpkYT1W7uwtGmSLbkCnKZwvRdsWwy4agDQu+VuFmcZ91Pp6IibUIsrD6Uxej2DutdN
8YFkbXd1s9F8SAuIRYkTMnbhKYO4U1WImh3yOfa3sU7IrbpIFHG5uz/+R6+Z71IVBvBKZu/7bJqU
jeOYnF6yB7gytgDLLhoYZxlqdhJVfaed2HEzuyPzmZmEQDwkedD4N+YCUKy+NAOKyPBSVoxRTd9+
B9+TDJ/ZG4m1T28V2Yy48gGDQlV6V5fJuvVCIQajl21A9caxBIqMmQuvDAcBcBBPQE6L9mBQ1xly
3Manit4BDKy5r0C2hUV9MPY8jJMbPsBm3r9vH2Mcy4+sJsDPxgc3IvQW5rDZ8AZCyhQnxfDK50sp
4+LESWuM60SuCTRIJNnzfjiywEKUlcBkBVpZQ29tpSYA1FZYgiavtWAlGUTH9sy2GpPKlxHRxfng
Qszz186bmeaxSJ75kak+Jz736P0UnDjJobAuF6JSvCDdID/7wDAHdVWWWL8qt2nh+71K1AHevnNV
T8rAdUp5j/SJ5HKp7zRz1WayiZMVpSFq6C4XGM7vReWEC9wlGQLL9v2XM/KslKOS0jfW69zvo6XQ
AsaDXJMMFqb+XJd4aAOs48xgnGJpZzl96wqQO8DoqT/N8dQ1QeEFL+zjgTAWB1A3+rASnS3nEnvu
IRL4T8P3JcxZfn4Zm+/imV6VmyjH/Tq4Jqg6KifO61q6v9tZNUCon+9NbedVCCAVX9j1c3aPofel
fxTp1x6E6fYtjguFnhkVaU+w5BI55rj/VtfS76lLR42bkW3oIOXdyt2tG4FUH8y2zA2WHaRtWv8X
pOvW63G+xuPkWeaJ5xLcJH3qn/SWEJiDiXLhti/DTqht60PIOrOIpPWXm3rV36qyEoh5CKl5dTH0
G0FNpXM88CeCuFD0AE3ZdWohOHK/TxsLGFFZmefEFsZxjYvzdD5xSkSphE0ZFfR9cMGg9UYe+Van
EoVxOdMQLFrtbpvx/UB1ulVKwDaItkvt8s0hsG414LenGa620E5GhQD6skLn39ZtMluX6GsG6LaM
UggkLKasGqBW+q9U+4DfrxkHLafVdG5yHcEaaf15I8IQUayEMz1nFubVG5gnIO9HMWFtb+G0aVf4
I+QDm+xZfhtHKxSwraU5fiPgSWMAgZJnOxPyaF/5AX/dIzPaZ0Zv1Z57NfDpG8rXopb1+N2VigI8
gqfNm4v3KSRKOk+PvtuVfNqz7R2L5HX6O0iUJwAlDBAODQdAnql//aTWRVa/ug0zmZcb09r7sbFe
X8fhkcGNzGbwl30u8D5Oyu6Ie/C6118Gix2ZvNJOHS3e22bDajA0L/PLTAJhk5eDbtXny0cF5/vE
WXxkvfG7Y6vZDOR5E0vmAXIAshOTMR99lcOFq314RDDP0plSzPSKuxgn6RpAV/VP5cR0RGSVB+pF
pqmChCxDwPQAaPn6Y/p6xXsQPvAe5fK1A5zxl8sIhGI87zGFZ84CMK0ZWJz9cfn6sCLF+jfnUr0F
quBuZ7xoWsKkf0+Ys/0GG17UdkcWDAmq8J+A412ptwwBozcBOWcmN0d4xax4R9ceBICAFOY5sElS
+LbwnQASs4F4LqWuQnCT4rE/ugsMDXmTA3OJLhpvCKarJj9ThCQ18MlWCCI2zeznwByusib2A9Xs
7TE2BhQ9IzDAQ/CNE2FA9BoIsTsDhWw7UHlM/sOdwLtSP+afTmP3qdnXEVClztJfr8TgH2g0SNEV
nI9kTr0MBo85+XRnazHLql4ptnlCAsPVvg2QDiPzl1ZC0Kg22W5gSeuggnlBtJShezUGLwunEqnb
jWPa6IxjXH3/EfvjIXa8dfZhTuozNxpYO55xK26SCWBC7uUIkHn1RJwKUBE770/1yz+JgoLzNEFx
ExAtMPbVcPINZBRzIfJD76mpS0BZt4P4u5glfP1wYyeI6o9r/4nI0pd0Pdeb4UcJ/Sn9gLyIoMFI
7+XVX5tTj9EabVxp02QoMZGCRQRlqyVPzp7vJY8F4OhWKCdBcSkLFoGuDhpz8JQ4R+JrJyJ7q8F5
Ix6wXHH72Ro0CUO11jCO+WY3UHmhFW48CE73epJzTdxSH2lYe1p2qGRJDghw23CpKnIMAtXg9S6Y
ZWl8F7GkNLQxybkAX3VgE4kuEIb/XUfrQpvzskr24hUy7iplKOhBBRP8jd66WXlXXGG2Pnpu1uV3
RWmE7JG+z5Yrvv9pQChxMZbRHMCchWhOQkmCbXdYM4E1VZwiLSEYCjdw7RbSsp4Ty2QFYCQl17mB
mgKZb6QUbiaqWogMMyuI7mc86wp3ej6KgfhwSrOCh5I2Lo2c0QCvkHwei11i3QEyOOgh99C+wD7b
vgycV9Ww7V5GsgqIiO4nEJsuCOEwTRcoDsnv4f/19L9rYbDN73r/7HhnTXVbYMvrzuK+FrjnURj6
aMWndTFpNkTkPr79hCYzBrxVY688yFzuHYi8oC4uVaR92iv8SiBQkeFMlAjmS/3dPhANIhm4uAW7
LjwnK1YA/OjJObg5sOIN5LG1bxFogvRjb6FGMh+OuXcgEE1Ro1pe0SWc48Z1sQ40d8ed4zVtVQTN
T8nWzqywA5M4kYVoWydkasUG0LZH5WIcXthdmLC12VLuspKAahMbfONhy2fDssXLC/HfHXYOxJ6P
QwlM+rqT1Q6cZ+mxa8633PpUc7btNnTbGIq0NUopfVTUk3QmQeC7nAeSrHUkbAGyfToyGMAXXBFe
u+1+5Nq8oDwlW2Som9dEB05d7AiwWM79PwVnkQmjC6ybWC8XYfwq9yiJlN+xGcUHd15MSqB3H6S2
On1WO4L1SpGKv3LBl9dnQydLYsd/9twh8dDLrsozwsE6uU9U9EzcLQB8mHyIVhjAWDpE9SW6jPta
zNeG4AfP8ps63QBRyomj5Dl9pCZQX4W+UCbpInepQURnkCFjEIfMG32lTKa6el/qQcnco8xT/plR
h0TOFs1I4SUyVpwqJZyz2SNZtxw8pglrQRgkVNStG+jjzAFfUg/2M61BUdTNDlNcoPfNs7eE/76x
fOhuVmsRoB1uARrG60FV7rI/aMfXeS0Cay8XepbXaS+CamiBbIpF8ZLSG430/t/mOVacWMQgeKj8
hOVc3H8qn/5n2dX9lwhy69OR/dYj1Neqjs+xtcLo4FS04OfyJd4l10UFPWRqHU5Df/oSt7jy92zX
WxWsFZx8XQMHsqtxdc2NNtXXsEfSGrQ6M/rDTIsZ77y5LhH2nLCjYz9P2TQHYIHmPKMXpEJFadUy
9ONteT4LccDYFgNB0hdjasCrnjDf2LqXrFRjSsm7N9II98f0iWDXAmZUvy9veMOU8nMZEa0/+q0t
caZSqYRwAV652Va4ET710MGbkNUsMfMSxla1fmdP7hseh5W765DqqGwlh4EV1amQHP1L2dVG+XPx
TZEuu2UZzrrfN3Rfomd8Acd+dEPQ9R9zcfrE0mPBkNz0BVNGGoSzqTN6fvimOw4jjc5ri5EChmfu
JPR5Q8DzNN4KXXl3Lr63upCBo8pdv5UoGcJhqiuQNdWL6tUKcMvXgBxDMpGNXbsiOWB0OkHfjYVJ
Wnt9REQJaKRxnXtgVfezUHVP1V+TdadSq7g0PKatVIlYJJStj2hFUmIpRELuWPFZZQD+pEeZskWu
d286qavqBEWdPT2/jNyU22fZRH5fhQHSWR7q4QrtfQA7SqIiZb/0INpQG09V1W9PlPE7o+h4Obcg
a9LaxYY/Z0sL4V7XtOUMH4cVtZ/diHLrZuLWp95lK3xnlj01+qlH33fPCmK6+OgbEVuwqvo6/sOb
wcW4McKdCpkS4Vxih8ZWjjfskkXVlDPsECDAjUHUFVMVWpvEQUOWoSxQ2/L/fuUDjgZ73lY+Aj41
BP8B3g0M8hQZ0qo+XAQMZrNqvhAhaGy10Zx4FTMotwlo7z8nwN6GnV7YRJ4ZVCwTl7UBi0ysdVbJ
7xPkslaaqcbY8WCh1pqetPE4ZqDULxzRs/usbTWcS1MTdSYSFC6W6oMaxCWuh7cEkSN0vQ5JZRWx
rvBbGhk9wlIJfSZ7bEX4KC5wMgszOQkCalB0+BCIR4cnYcmyTjRW2hGinOBuV1G9q3EALJ9kqzY/
504KPcurJOTiM5RKMU9KQtPqJ5VX9ip9UG3wN36z4WtWmb19Qk41LbhzRy3o2R0ez4CU7b2Msseb
/kbTg24dBaxk/8u3BRKonnVO9czpuzjWJnqVLIRrRtnWeSy7iGV9SMrjNxMB66emLHS61mJZy/Us
3+HTNdBu5AW1PTT/tv44rwjhFS9KlRvEXtAuWaz8N0tSWG4lkriL8YLi6F1OuDm8XBHeO9Ak8Aqd
5cB5PxHbSboNGwG/RbvomnpTmCro0lexjkPom6P5qNbhW4/iajedhSxjJ9T1MwYwG6ZW2wCo3HLX
3/K0MFguJu5MfT7qTRc2d6XRmxMmtb7/kx0Qzj3rEPu08HaDc2D8BF/mlemMRe6K+gJg+R8hSBmJ
nqXPzHLMYBX0rXshI8jU7oF/wGmhXuJhFQ0S4V5qPF6FT4mkWbmg6iKxcOSCZFzXHeH05Lyic0LI
1dWMMAiYsOjNChEcaa6Q43tKkNEiVpW8S8Ezq4X2E+lWkPcL0QieaQaDfjEY6owJs+ueO5TYXZfv
1GfaBfDern5Nk88ED9/cO26LFwepp8fLMuSpRGvJTFozJVf65LDuvv7yA5KbSaGiNmPIVpeKyeMV
FLujpbkN7YmTzliwT/kyTi+bC6awvsL+vitmH1VHEkhZNXMQK4e1QietFjIp3dCY+mCYMQGVjvKy
p0OvjF2BGP4cVlGtfeka2cIS596d1x39S+BJ2Gq2EamZzQCVOQJf36dckmhdm3wEVAeXlMlqvtfW
AQ6PZH74kw/hjx7B48y7398pCrTQmvgEanqOboP99ZjnSxpPyREFyuKBd72oglVpE3r0LqtctV8I
fc2opb6qxvgQncowy7w5IAy6Sew9ralbQYSa4NfIWgxVS18CqiFZcsX+9Ot4wOoBre9kSUOEeVdz
/Db0OUtAyu6xdq+usl5J3xx8bfTaqlBu54rv8puHZKQ1cErm7Ha7EZ0HsG7roR+wLH+BxX3X79Bk
P98EQeOS7OLpdstbr184s27WuFdGALOGWGAfeMfK0nrI1zh3fOYvf2lbgmMmCxQEugpiYkPRJjUW
pMPxwAXm+BDXRSplcVVHATxHedghDZv2xV843MRt3OY5mttqjSH9PmQ94Pes1RAJnh8e1Zgx+aA6
bTU1SsE9Y7i3v/GHEtJhPVdMcixCJwqPgSJHV5Wi3RhL0rVRlOwUUDUwsK8QIWCAtw+LmElk2der
E/J00nOdkweO5VFZs4YZtL0CvQyHUagv3RSy0XISc62sBo9s56l0zqeOEXSOe6HrN1byMe7wmrCH
+2f3UXUcCRITBZBlL6XqvjumQIg1f8Fme0KoyKerj1+HSrf9oPInI6TkdGK311ERX4SbIeH0JE4G
4LnC9jueMMKTioizb+xOrvD7o5Sks77tk5C9bbtwhcmREhxUAe0aBU9wW1P/sHM3Pq0X8sb5yoOc
T0iSFf1USyvlzqrUJzcBXFhNiy2g9PLHIb6yTX1Kh1TGkE671TH69IkRGQEBwiuYelkWFGcKZlvg
4NH8Yyos1Z11arcnhYQnyxA9DjHoNIt7jyrXapPje7Jmia5FgJKl8s0NkmLJnNA2yYKR5HnSb9Dr
p1TnTAr3oQcHoGD38DNQcWsf2NCl/mY3jR1/ZV8Q12b5k707Dxdv5EINhwqE3JLTuASJEcwWa/gf
ysvZkY6/lOM3xoYxlj1rLHLSdSpZlveXUEFxuU6iCFaFYRJ83MqUM7fJAwy5kqyUJkFQORe3Tfdk
C4MJvYUqMzUEhZgAS5BIWuziQ/qNPTEu3CNMJci1aeiiPQwd4i3n5iNPAi3mPii5B3D4PHKQSh0b
bcyWKMm3vTthkNiyigD2As4ghAVjiolcxXrjZWqU6j5wJenV3xy2Fc4FgjV7X6uV6owfVNPQc5rg
Mut3aIFVl1H9Y5KVGulV/31yamcAaY5CIGK5Pr13GrGrgTyhfJpE7Guqk2uYER7Ch8gPVxQVSQRa
OYOt+N7zlT7a0WEYvmnbk0TQ6PYa66AvXp+zKSukeHRpwy3jpKZey/R/UATXWT9/8cCmK0LyxgfD
TOAlmCJ5s2sT76JYeVhtUw6LDCd0gFlsZCDmMhBCNYl454LdWCryyLoZ7pG9wJC3yhNJAT8vTr0Y
EuxkUZlK6KH/Yyg+B9JhmaEO4/acqg5JuEgy+mU5CryQNIHuyFcGSjGv6TqXxXnzrJCNpFQvlF5A
jYLSjRL09tVOnJ3Q3nAsILq1jHBfSNi7a1B54vwdSsfcYLB7/av0EeN6ig+mibxPeT7OAa31mfj4
gflC8dUEzO4yERswqKXbd21qwoZfcKYyjI7yP4AXWjtmcwGtQs7WWS9kOOAPD4gngEfeBtin1jfq
kJr4+bj8yrF/L1nBBMUAi67H6KbNch/AdAkJK5Iaf3CLpOD8JbGCmVU3yiRT3C8z2JnZB2KAs8KY
eIPEYL+LH9qTfDc3mGwe4ld9LSP2jar0DPBL2w/YUYMxlzTJwFXNXGIXpVvyCrUvLykRnIeNdCUG
FD2uR62urKdk4fq7wM3DzRqcIfyqOLXEZtG/v/Gt3uupcWNaQoRY15DPtug77nAheixSZdr2MFn1
J+ewvWxUqE296Z/Vorn5ljv46y1JTDfOA36MvkFLCKhEPE/z+OccNoOt2hDGz3Zbv2UlFg8fQ840
Da3AsgYsnIc6LhtjmzDCKdojYnt/sb6yQtyNEZY54wK/Wha/+R3IJE1fFiCzCyx/bnAvQVTc2YI6
DzrQgi5Zr4XhVXNF8iEaR5yfKZyynrF/arxDyZ1sBs1RJS+S8cee9n65b6iPJUWuzE7/kP930pJQ
unS9W5NFrHuAKF2Uekkp2LGsaMtTtkpHoeiytn1MXHIru3/ebbpJbjaW43O3bJZ5vpnj/f5hb8ph
7fvNvFhxTrlEy9fcUVVj2aPtyOxHWtomdrjV7ipFWwo1itdonTN4/nrBD6HdE1O+Ub9theUmu1Ac
6TC+NzNUCZH1MTaoOLkMFZQgOLzz77LW6PxvhKjj9Yx8P7GEmKLcNKCogTjB8cgqFncx5TcOrKtE
XjY7MVoUw77URF3yw2JwpgJI7G8yBuApLyhrtZzmUHGiQ3ELhCY0TwWN1i3NCNzgrLNvZ1MJhOi9
DKlC7TyCXS16EF5wbwBofFEWoyyVHTfYUBfBnpmEk2URyYSnduEq4WHAwBdnSQmCHQnCxMGO7uSI
Qnc/mg0epeG5siw+MlZ3lcx/S5b8y0Y20DbNYnNwosEoSuV1jGoXCfFgIRh88qQsrYNRc/H87paR
FhOTs98CFf0g5Kw0HGyCYjYZnz79OdflD/0+HtIcUwWCmyZTd7fWcHLEwnTRTqXFjw5p3oK5yt6e
6pnNsxqZhu5hC3lvo59d9oo32BmOIOuxmSYbHvqOlrYwTuK7GC4d9Dof/C4dQaF1lgTu2oYi4iu5
ww+W6voIz3PkZqTAkUU7hSYh6z93TDq/SWPrih06bDfDF7+dXsiIkzyIvIZPLoq3OlOQr/Rp6bmC
/cpJXxBslk4oehKFM1KFeNCbMemDiAk/3ATUddRcq59E2mYBnX1Jo+2nRwgP6KbJ68fS6wAoY6/o
/jI8Os4UR6t5KX6FqC5KukbeKh77q+z9HNtDUHokevWDRuZeTMBPaXvkvI3KAmTN/3UC4JZ3Pqw9
Eqtkklv407IIq0+XloDtm6hEdV8Hygg0b8wiFL3e3wysMaof7rFglJIXKMAKBFLLzEt9JRcb1+nM
p0id+aQFzdGal7v/huc6xohXwBppMB0R5wRqM2xdgqmprPMVQWTxS7EDTNFhGEDvAZyvepAr6pIt
pAiq0Yun0rawP+NkD04oZ7MkE0cmQbCpJAbHJH4XRtfOnSVxU/aCu9tDMotHUM/vgm8qkNxydZUs
DehD4VKeu2zEpfco+R4ypL8lwNXRzrJjcjJ3IfCo1lKZxYw3BO6w6EzqEnkZnTSQkSosAnGvj7DR
mxobNZrUWbScpvAu8kY7wWfUhz7g5O4D6/p2sgFbsZ5+pGNhePcLYcZKgtfP5GncE0Xj447nK5Ab
pJGuDhmNClqVB3vEImt1f0sCWOOJbdbAWDY2Je8NYJI7sIhwhoYSRn4N9ibDZYFuzrocW2XyXBmX
APTsHeetY68NwOHgHbczeIVZSOYUp7CacKaShf0gafOXWwdrs2lKCXmSV5u2EQE4AMKqmR8M+Yis
GwYymMZFziXTBVZhkEeBf1dPwpTdRSnaBytcXg35ESjkOQt5IqZOC37eqnFuYP/op8qGk6rWVxxS
w5lS5GGQhVFRLZrnd6tisppIWY8IePr5o2kuqbnulm/5NegArhoVQycR1/F6qRYOJQt/mDgDD/i8
FLC2csLxgF/6E2lJdoR0GodHi9Wvb6WGl+zr6qp/7W7D0/iADQkaOLLNhS8xCH4GCor7RsnvphbO
nzD6P6mFpaU3wwOtu5LgK2KVDqtscXWd0nrVxaJp7qvfPzO8z2eYvhekw71M0jP7dYbEuNTe7ixY
GVf6WbVL/c39BVLBLkQ08hT5SNJjymRICua1zemPPcHifr0XA39BhGpyl4ybUe5FyubMeHCD9IEA
cUAkAFS2hjeo0mWmWKmRIk3BwOEC2/sVmI9gw06GZipINdZlUwvyqJsWbU+M5g9qskNWRAqMhoAH
RRBDlJK9QWLKaZtj9PgT7kay0c+YMhXIRwd8dxkONocbcv+1osDauWXfsDTvdeLHWMyqkTXF3xUV
fy7nY2HVj1PO68PPvBZOxfCnJcSrdkvQUDCJzIRVWGl0GMElUZ8IWCrU8XqvMyY5Tw9fi81BAe8w
547f89WVYrPVaVlX6Cu5PwZ3zTs/JnT/76T1QbnI4OiFB18Ca60p6EHw2VrdhlKrkHDi3f5uMZ4A
5PsDDEgMJ5D2sPDep+CD4rX7tAALurxrZOb9R6pZE7RJv9iJGqV+DbqJyz5srCFtJM0hMZ/27Ux6
dqpf/KpUdatlQmF7JGHF9AM8893JgAfjbC63QgukiBoJabH3emx07A9+LV+N43QjY5K4GRlPHv7C
USQPAywbfBDq8zcJeSAu+oA0YAGbTy7sL1bU3/SmyYL9pcqwdIOfsPI5Xzx2hzChJfLMWS1IZHji
MN7EGzwo2suopC7tNoLleLa4YxcfYWIZVoYCQRTgmAK5KlrX98WpKM8tdhLMdFVlPSVt9fBef1Ki
GAL6zRtusiNGsxI+UKBFKzciXSKCSMt2eoWD191ufr7fxx3t53cTUaHTi840+Lp5ugc/pcGefFcW
GKJnct4TcqdbaHJajAmPOz5sC6IT3VTK/15GRbqruS/Sk7heUuQ0cKUIA/GtasVwQ/g+uL7PZoXR
w7g13w4DPVq84Eyy010Hm4Uwe6597uShloqh/vw5VeUrEUaNKql1JItlqxE8TXBTUMAo4o5SsIAs
H5+UFU/oPDhBtsemnrvqNWL1XzDQVoZBtY6N/aBbc7OQYmvFcHpdbh7glmQrWjyu7OdOcArs78yq
tj0GKJhbAWuzAddsCqW/RcW0Ay0uf3AxPQwu+lYkcPU47sIJ4mfDDf9DJDmQVtcqCz5Pvk5RjgdB
toXoe3cFeTy/0yXOqYFjKELP4W84Q07eBw/Pe6gLBJX+FKds2kFWSPvEjcmZGuQpXdlka92vHbJv
OmyLf5Rvsi5NbBgUCMiVYiwWfYZ584CCrVtx3RSxWhko8KNOH4VXllkpOJSURrVotnM4gUuO83pq
pQ0BEFZAA5hNPVHhVSlaIPTHu8RBoCS/81SDUlTdHjWFhO130ZZnNkKIHPnwqa9ODzEMotrcauAH
dn3+GnLkRmwnrVB8xLPylSe4lVJJISVI8dbTkkJ08MiWpV4/lh5uCgl6883ln/4aAqgd887Z2vQA
xFTt3Svn/HmbOD+y3rVFa9SzzlHVbLIIikZsCOEYTkxU2zNPfvXY77NGa1FtZw4QewIb4NOtfpUA
fwvVbsx2/SV0af03pO6GMI4Xa5f6KPQuaWNziWCdozo7uccPy7JqFX2DwQLTlwKfdESCe1V6JlGD
zlGkdopFl4FS9rJ/uPty5E0MDy/3NbVc5TzdOcswjx+3eWYujNRxrny/aKLf5mrKMeYoLS/SBN1k
EQcoc8zFvgepQZeDSMr+VSfNB1rRnS4SgAlDWJpgfFWh/EVdSVyqziC1z7ot8C5tp+lA7hG/eLZ6
tS7npSiTLv363Ogm/SxWgGGa2i0EVYf0eVTmiMvCPHEjRaVUGL/4V4vlXbimKvFl3ZefFOcfOCnp
H7X/3qqt6yYdkVr8ijdQbD3+3KjT9A57XZj1kXcl2yPON3nrB/xowiY9uDWLs5Lbo2bMvIABiLzX
LA4dv7ilnQhcUXw58ZJ+5n4T3nUt8XVgZ8VCmTtnfOtfMAlNqrReHazsv/x7JkC3VY4KXXBH71zX
SltKHBmobH+nDIv+jmKTj8ldtx/lHtfMadLKR+ZBaFEhD9/Eot9I5LfektzKN9gfo1kOJqvYfIK3
+fpuQFNcowMFXqtni04/kqiqI05jj9k9G1a806gVe4Fwqm2IzQpi8XckFupTQWcEzyVUjnq4BOFy
Nzt0hhgstpSFWvTTVghDrzmbz8WOxy15GYEZTwC2kNXQjCW28ilnOTrY7ewT7+qxhKp/+/Gok9yz
K/3E0a7gX/ZYUeoEGIiBjxZ13F6UIhKQuhLiOK+BVWjFqetalVUp190sD9CdsT3xQt3eYgK2tyhf
yu5uR99IPM6HrR3Fex5IGsNPjmHjd6g5bmjBuWm6CTH0KKFnP48ZuG6t3W0F6sOyyBwGxHxt5l7n
BaSUGt7SsWwSRjDpZhwcLNAk2zpXk3WXmvDu0OrEqCRa2iLUP1en0tgQN7PAehHInKGRbOilTX6F
pBtaHK5Ba3qtzgFRItFyTkKSwgXwfH4do4pgQXE3PFtpYR/MJJwnthwVsdYT9uaJKR1y+3R8mWG7
IazPxmrO7iZslLSvzmZOwgkWkfy8iawf1n446YYsG46vIeyxWfw6IKMcCfq+y3NWJnmkVUVyXFE+
bZq2z4tQLnanPVz2xNOctYwu/+LulUbyJA1+9JMEXTSCpgJ6aYRni0NotUgutywKX+thxrljij0j
iurw4OJDVQ+Oc6AE/BSX8mgafpFlY7AsyoDsyftJ1a12t4LBBITJgpbWbcS35klTOlatV6jZmAl8
9ODBEojFQC0sd0dZd1Tk5yxjbGwNZijVseq/lmjQG1NbBXUEgWURKo/hzRqjqDVXa8qye+lpXTrc
I/mGCtS0d5gnZaQENZpN7cSdbSIf0WmLdRfUYDRD+AhZVOa5Wg7jUZSiKPTcgyxRdnujCIFQLhSw
AZq3BhZ26Bk4+2GxkbG0cs2yVpmRn+acf98sQzo+MDnobVxrwkhp4uxN/NGzktwB8+raJTEWBt+t
rIieYBR9LeH6xmqbguX82Ck1KzEiUXLRTrLBoZNwQllx6LrTbLfjbznhr71IlwIqxoLb9AElptgv
t0jm+DYxQ/QB8S9tfzwI7y6iaZmdYPalqEzBKrms3XgBG5NGAmMj6Rql4gVeA6o7Ty7wOONsvzoe
/qnLJ8zY53DZ6GAbhuNOQA+0HWWUexTn4Ho7a3roJ5Q/RErSSgxr2UNhrqsEYyfBg5eJWX8lq2ll
GqITkcXA1vlwXCEwkMMnLN77I84SYxeZ1RChZqcloviScfBwXxTEh+Rwazw0fNTWre+IxVxXv7PD
R6EpetAWrI/3rFU5+VE+hzA1Hjs76vD2zHMKkAElsoy/vJ0683b58noqirzz9K1NADkDS1AOSQa6
000oW0oYTpeqTtdhf8/iaBaqMC+id9LoFFHj7FEl/H7CmiwUnIcVeie3ccoTYF/G9TXP8p1gtfBs
LcgkxKYCCstI8vlVdnATYoC7RwoxnR7a9UT+48CnULoY0I11X0rt5gu4/bOWCHyPqLolBCVQDm07
rs1xCwluihmAw8mOAsr+D4HUgmcyOFgNQGReq+s/yigbllpoOIL6SfRXXs8SWxUS0z+/TBPM9cWt
CffJv0wJI+p0tYAHgj9tjWci0Fet1M7Fvj/ZsGVKqJdLDMnSy8SW6EJFwPuO6IiC/k2d8r+mzA/p
5KnV2qgyZW/A3QOrSLDELJ/lusJ8wKR0NBOrNlIdrseZIs+0sLVso1x8Bi9z92TlVdWsHNblekgl
wiAUZ0rs7wEw1Npnoec3JHS3QsLP0btYDj3T64UwTlbZhmSo4L5/21hH5tSaaj78y4ofYJXR/DTU
WC5m814jzUi8b5couRRWKE9Ym3QkwphlRvZxjAnundbJxEQVsB+7vOG0SQQD1eGYYD1S+/7yumnO
EYAw80cp4UDak7cnmQ8NHB50J6S8pvt/VUzBp1SR2dgzWfcizqyeSdbDD082cLFzR9OYzlSaiQso
16Hy/kx9njMrLN2Ak4Wx1kMZeC/5NjWnYRlon4ixIu69nuESJgIY4WRm0irPcmv0xItQV5Hj99+E
UlFA6UWgCnkMKw44FvoKb6MiV7DadloxaR3PMQ1A1+Gi1xqRb71TWpBIDTkhcs8avMgdvu+pj7Rf
huEM2mwsHhgBnxbvIN3XmbM2yy850D6QCVl+uXHO+eZO/fB55g1N6MqEX41DEcfoP83XfDiCAUFq
9aT9EC7t/mR5Hw7jQhU6yAxAuBxd7SwjsJ2scdFQkrDR+ivKgUJPTiQgaQn2RfxYubOFPZZKvcvN
x7KN12J6O75apaYADEMy2yqf+yNgb7IwxPm8ajIyzSh/HawNjg1fIMtAsxz27l1fgNqR0V7ww22r
RqmG332WyllxMf/W44ppfof+hYZlwPTIja3E7+2/N4zGCeOWFr5fHsha1Xpc8xMhYcC0qUeeJDV8
ZdvC/8v7hRyrwdFgznzSLI3GZbcx/IVRbtL4XZJPNvPfbfH7LSGUNKk4gZTF7TsWgJfreThEAj/m
PU0OOAIWEICceHHU/NPd4ZmJGueExwb0ftfna0iGo9HMmZ58hXAA8uCX9k0seA8a7nmGeq9tjXeq
39oMbHUoVCuGBaJ1Cif3h9twdLGfXGBlgZ9hCVXWgBgbBmRHS84F86aLTrfv8LEHO9j3J7eoqF55
dwhG+b9ZM2SRNtMMi01HXNR9XIpOa7iLemvHPmSHzmUIZBrAzRAwatfH0Cy4nfI27YHm0qBkDH3i
wOqNccznv3zA2djYxiZUph3iXO8GTr2JjSSptC82G8Hz7BLICYZMjXnh6AXaHrf8lP+GjXRUCvJk
hIhs199WDX1sJQs7c0C8GaT4eV3bpZna2da+IQ9uMsnEXztrGcyQRSr4EIiElv5zuNy34SHTRNri
6mFXgbMLY5i61kLwrbedobixuEubtf0h9an3OQmCweG0Ayw8p4W6U5OH+qaGIzTZ6Q3qDMmFm2gd
YcXkKc2uaUFuIClq9r+YMgGjIL92lJbqDU0J3x6zhB5bR1q/wPAumW77vJ9h8t9JkO0KpWg1ISnu
NOtIw5ZK4kA3Xhbw1G03gZC07IveQfZAJWypw/yeqiSdmzprmzLZaKbLypkQo7GsdOLk+7iGZ5/l
qSUB4ZqRuDW/KrHXqQ/E2H6GaSgB2lhBfeB+Z31twY+AF4AJS4gQ8ZZe3Gs6pOIoivmJPoq3pex0
1WdE1NqYe9aU7sakVSER/ceRL1SWLVh4sNAF4Jzl8zIllQBmKOr0HIGMYWYTBoVHkIvMH7aTv9ro
Q3YTAPTEUTfRm2MjkYnOiUbDu8a2zFbZygujiYRJcuqBxxNkrlUhMeVOmgQJeOIWvNAKqMDR1qXJ
Ok77c+N2BXJYi1OhZzbXNN9H3XosJBuQ3ry3dOkRnWwIChq5jwQkhAaHDUdDYWJTFfW3giAVkbfo
hG+XxH+nkP2dO3Pzf/SjcEbRt/EI7GPk1N40sfSo/ImoJBAdMVAx9zZ5P3PRuvtGXxLfA/g8uhG5
rxQF2mtcmp5r5GZTI/R4vGZ8opsfDUec3PMNc0nfbDqyCJNBfSuEooahgUeURHc5bOwzp5PfrgBN
UYchyLflxkji583VjTq/pS25uOtCA8dEaFFlIoM+qY17u4lpU8ircPYAPA3hNTcYJJRmWMroBlQA
o+ehLziz7Lx/fx9OUuqdW5klykCNnZkN3nL6NhDC+oe+1In+0ORsqmnyZ+7tFK+1iJwb3A2S0yji
TE2oaKvK0zlZINJcFkaTNQIGBav0T+C9HS/eP0rWb8wmJygHz/GRFE1Y7Ere5lbXpsIVS1rEwUz0
i+gfzL9bktq/2z92H7CmFn7SW9xsJ9cJ+qlZMSmuw+4/JDJSlySVH3dS9UL4zbdKRiw9+TKtnSEt
pZbTNLkRWgrDxCi/bDtEB4Cxd5WJpKEBlKiBu6m74waQlFUdVveLJ3/uLlH+PLI2cyyrHw9QlkQn
/ty9yB5nUQTvCX34VH4spZRxiBoPDO+WdXxn1X9/YtylheT5I9dUlLrYOEOxTrwwiqLtuXhfzUIE
SHjmS+PXYo2PLH6tAkRuH6RkYPWio9y8Zso5dfpLcDdnEoreneHnr19o2G05Lo0fp5Yrt0JnNSco
Ap7/Lh3jDIkCdeXzYyMDaa+U0UM2Ez/skZuY7w7DoftJuX4y86TBgBB1c3GKDStLoXKN++GuiE4R
JBDw7MTKZ3LQ3Pa0pVH9GZBPkKb2o5jWpdXiP0wKWrcwcNp7W5bDiHPpdBtHJYJFX37ATpMFXRwi
Y6D3a2/EMYIu19NUktc2JnTNQzYFecKGSEPkicb5rR8L6p1c82pmTBhoiej1Kr2GS2I09J23nZ/4
0GcOpbutQDfBYvm+woI3gj/0SQStxOF8aHaEwUHdtYjBf8WEjPlvu+DqAEXS1Rhm0uI/WfpB3Syx
QvWaWFUs+H4VmQuXNzwYbWopTjw5MZoGqvZQOZFZqmeR8D0P5esBJWlcCm1QRZObDybCGkSH4kHi
cq6mkZkh+76pxnTohXp79nImueUZRh8ZvmEEKTgyvADmfDbwmiN35ar1ayN2UB+0+nBH5L6X8Fzj
bgUTrnGjbTkZuU+6jYY6oWC997Oj2uWRvfAmZvWm5I0XjK+f/sQWat/lSjOjfY+XY4j1R3u6UVt0
3eYLvCY5WRVSkSqYkZmtLV0Gkme9skJJVkoCqfAFBnDfKan0qq9mh/m4QOjNmw6d1I1ZsQqNHGrD
qF/WZ06ve0MK/jDct4tSVD8fWEUhnjYIQfvGZfuDqNtPS+Q6fqbzdMZKyusBBiTNPDkXgjU9qA+G
eXp/Odc6lXVZTCoHe/txa4v/XhU4AzSHeXEMx/ghpEyzSlqlE9S6kFHyZJ8/ZNaZuk1kqmkETTo2
4aRIPaIv1TT2sDRk+NZs2T3cDENRe/UKTwBjLnfU1lNqRv8BUzPJqzGz9U0x3TOIayPkRJILKnEJ
QqIPr9J6d5okuQxpnGQwQvC9+IYAXdda8ZX2VBpEFpg3pIBoH/3MtPQKuzwJ9/9qfS8NJfmQqsAH
rCDZbgBJZzzD8Za3lrUFh8QNLNtEEaOy8reBUQ/jLQ/IOd2PXcL2y9K74W4iXJFHzyDX5w6M2/9R
OQazHcwvmnK6X+yiDkdd4SVgqev09dQNsborVCSHCaW5qbegZaxERgt/+aU8ORct+uBaWiJKYguE
PL52c3sh5vFioKo3K4m01lmLHCcTlGfjHspnHwU2pTlhNrO6MJvVi3mY2Nd4AVyrI7guVDfnmGDb
t6Yvx16KCBJ9baf+QaOvYcrzyS4+6tEZQgRe8TDrfQDcDiyJ3Qqoc9v6XxcVHGzhspCoFATKz9wN
yPkdc5Kpzr35+J8aP2PKa1WnjaJFmM2DPzUDBDYSVcHCQIzc20XcQ3vh+siYquR5M462vUpy47X2
qhdWcc/i8D0lSNB5FbVvG13k0P3ya2bZ0oRDLd1RzsSaEilW2ExW2vV83PnbpbPqHfB8AdmFZTU4
2/MD46uwjkjGrkeOb0Eal71BIPAFg+GlMnu5G9p4yWKMLPGleQQxO12/VzcNDkVnP9dPyhulgCaX
M8IP+ObMtoZh/1BD+VfX2vSLWH+27+5BTEMNNx3emG6Lafg6waagf8xmcF0lEMmr6rHj4bjOauSK
8YCANC38pxZaUIz4SGJxQlV8l4F1w9wOSqFE7KwA4UNmVowabrdCXnoPO/qSgBMqkP9/FMt/DFJT
F/216IRnLXtP//oSGChhqCsQnP4RQRrFGCQwdoIkok/+Xlpzev2jK33oYtIJejrZwzfx03l0Mdcb
Y9Y1zZUygio8ZfTwVOcxq/mgGMubzOX3NXV/7HSQHFVNaS+zqk9JC45pc597SZ1+ZOmeDh+G5GKn
rd9zIsJHrg+sQpAPbpQcZLZ9olc98QgWhr7IstO/sRoJTRF1OgBLVb9A7AjuVisyqhlufbf+V/z/
/lPq/iFqVgAuwK8SpPzsBF8Q9qudMy6CDlK4i1aotl+fD2qvM4N+/Wo6KZbmA391/Gh3GhVwdENf
RALVnUQl6JIob9EEs0IjWG5KUWvvvTu4NwHfTNcJpp8bnUgU2Liep/mCpFyZ6oPZcPTGlZcbmgKx
kBswRYFScEA4HErb6o3tn2HlloLmHkaJpYtFeyVSoIltieKYBcnZP6jvnkCbceHYEmyhQ8ObAfwC
AtoI7bR9d1FEaEBuTReQRtBTXBPCzA4fKpk5c79XsZcWE7SvbuMFjHflZsXpg+3Q5jeMa1j1vP1R
ZKfsK4d4xRzf7vJOupcCutdr0b03R05vZKnjuUgX99lQU8DqnZid6WNTpJJUrgEcb3HSfQN/5BBq
dULDG6gIkZdIu/3D4TYh9ApfcikLFJ+By7+8fwH4sqcekDwE85qyk3htqmor3BDOPpvmIPZDJfB2
ptjCXAG2i7o59M1o8DHVkGa3NFh2n3O9hNaBAcXEgG6u7bGxx3/Rnofiq87Wo0D8H0miUnRXjQW9
X6jZpOklXN5xJ1oSqk1jPwAEUpcLX8791RfQJ/bQsfW2Ydkm1v6Dqhg076Ampsm96ILQGPMwy2Lq
sOVCkh58SFNUiTrA3dPSv3A4DHlipL1zYYuX0dICkQf/tQsJ9tWUh6Ykj/zmTu+4YIkZMysyyLSE
dZWmCt6NfH+gXCcTMy8Ba5vdrE2ohAHs/S4TdSt6Gv+jZDKIgBXH9n6vyRD5BCxjbZuywI7zTzj/
JCAaCkztDDHVdQAT+V0yTzu6jUaIrn8eA5U8e7FDMcFhE8rfhP22OVZQEATMIwqXaoRJVKCGaOQK
AToFf30tRPUya00mTJRfNRsBRhvJ4Ay6+ajJ0F4Qq8mMclYrTkGdybE0GFxWDUmZsO4BtlBtmj3M
mN+6UCC9rEdPSdBWrnA/4k0FI6YqQk5LywfTSwgR5monTA//PU12rabG8PiZIsLTu1Mr3NlZlk3e
y+oxGbeJxdnruizML45toINgoiHm/jZRIHfIbHYcaABsswzOdl6r4acpyu+fvAZzCrSr4FCGclge
Z13+Rjyr7uI+n+p91WWR6hWJj1kZrNIpBLMjCmaGbMei/Y7yD9KZfEeOfwUPV6qczPkx71Mmgwsb
4uiAWHBuFxg5kbP80LQly/3mGsLlLGK2hnMNocqvpWUnYYPOfPfLdsQAMs+xT5d5xBIB6mSajDFw
uo9Tci+6ND7lU/J5vkuXLunYQ1dPHAwWPTzl/xi8bffcFWMcgbr3P8chEI5l4FJ8Pan9GDbWIoYN
jH5kkSchN1B6RRb6BBnUodEEp3ol116ik4aZFr5mz4rPBQtP2SLfICOgY6oP4A1rEHDod4c0CKS6
pz9lWBb0l4xprEZtrm5kgKtnVIxKE29qYrZ/axROw7CRMkOG4AQI3Dxb4Q9yR7Z/gxQMV3oqHeiR
rOj5QdZRkET/ISxz7TZh2IzTQG0WsRE43olKr9dCcyKrbuX3H/AqQvjM5JDiVFenEtMlcURT6K5a
3CP8jh+FFK09gcreKD45mEAO/1QeSA+O/iBPI7dIEfF58AIA2vXXisLCXjcQd3a5CM3aj62fjHTn
VLHlleuOUqe5S7j++ZCpthB8Lx2SBeIhTDzfiioUOwNz9XtKwHivIhz4ILP83Ms9OZ7KmWqXcjC6
6EBisKhY+hdyQaQEAA/cN2Fds8RB0xpjIciQdBDIf9K+p2DoK8QmZj0JW6F1dQlzCZBNcbWnzIEo
tg/9daxeLrtsp2oSzhOiTzici8vlpAGXzmjYNp7UVDHx4KtqCko9sKGEbJjlDFe9jcx9Afs7g6Hq
E7Ycx7x1DQ3t9AIAZ6xFgBEZg3hksuknftJxcRQAmAD0GKy1btJNXiNYfWh/VS9mZAEzV2S7/rqn
gdh3fHCBgREPfF3+KzJIHfpbK/348OWW5iZ+MtRnf8xMwTt1hLOaYLhQ3yr/WKmDFBwn3497/SZP
3m+R09UW5MxbOJOpDqTzLm3OqtOk5cTe3EizDFItqtVKkk20hTE+VF3/Q/HUwqFSQM7zLWm5fUr5
KV0kZPGTTJ+EJBWuxG1LQQukV4gB+GhJy4WwuCjgMNDUrRE8qUfUsaDGSzOwOt9Ry3BKZEaG94FM
2pwQ75FA0MeHCkNrvVglofrXRMNwtrzXd2049K7Kq5DOfikw1fJzuoe6bnWwRu8Ld7+eDVQm4NOU
VJO15S1cmXzmyCIP4lQLCV+SmboQfHmYg2IpUdBpZRRndPLoUo+xZiqc4zrTIB1fkE/LpMXVSvDW
f4HpsTnMRy1T+yKQVFucwpQD4e5mBh7h4CW9skwdiC2y9h9kkG2CiXoaCAH0zp8/gcpHbngLi7oA
UmWGBA5/s2/Lf4W3h+WIQnUPfzBSE1JjR4xAmLvdr0gW1wIbfs17cftM13M/JV2sNuB4yISKm6vh
oBGJPxkJCsaYxjJBrC0r0ODKZxoMDj6dGfHxLhOVcQB0g5dfEDxTzKzPNaioyC78lTAViNZUjguS
HOEsFSbYrctHjI7Z5iT/iFOEAHDk3e8cs00gezg3lDmBZx+yKLFEBefoIVEzo2e487mwX7a3BiWe
9c7LXZp9TR9IdWBA+5Tv9nmCcOvN+1WMMxcPJJy0INLgS9vTyX5aj/wdZhNnUTY7pGzG7+qucZHG
wca7xn+fyegT5v2o1dlklEUKWEsnGpU+sqUmtAVNpYJ65krQZzSVLwE/Z5R97Ll9nWOlqxB4ecor
v7VxDV8pM2H7uIvMtcZXDB437Xg8elZvjdQ98JIIJEE+2pP0SB2mdkLIJfoEx3aMtdYs1JtovKhw
ZcOKpc/qiAN0g0fvWnxHPI/SVokB0ZGqn6i8Wb1hjwK8nS96sozr44tu0uGBCaja4sslnUT9xVV6
fNnYvxuSeCDAI5EawaBRz3Pa7bzb9nCDPXjEkRK4Wdhr+bDp9wBeVEnFk9YOC4X+xSvUI8qiafUw
N4t/xxhy9wlb3V6sgZuMns2Tb8yWNZK6d7MWYXsU6cHnfAAISzZvUSYl64QdveVA+6NA/qTDWxK0
hvAvhna1zyMyc3o77CadAX/z0kA87rjXi7ZPjmsWethGWlZhw41/6FC4ElOpdvNoPqMfQqMIU/f9
h678vNR1LwUIDEmSESUIgA34+sAjqevhYXM7+h2dl3g09atySBBImSLxDffcFYHn+Dt/oc8LiZir
r0SA74EAdTWGZ4DmXi7BV5MG+yLsdms7RAeTtcdULuYTorqGfFsrQqM+BWmfayjzbY85nsaPjDKw
jkL/ljPzEtpzavkqyioHkqosvNDUEwuNZAhAm/TpdS9k8lPsCUjJX6hvIRO9QCEHFX10+eIygQaX
5T2mIhacOQ5bHtdKPrIIfApA3DcHmQdbHm5SKA9wTSmTCpI51qIKKX1DuyhMNjEfdE7SqpGU3dPf
ufdNCzOjZO2vQtLCFdrCpEzsrChDNsAARdQ8OFNAPuE1Ql0Nw9mJj6psnwmZML4PJDPdXFw66hbk
mK/bgdAUotq9zBwaKnwMKtET/QMNfJu5Yp27AFMOBPbVtjMK8G/nkHi5nzvF62DupuKeXSgdTk+K
/tHX4WlcKf8YPxRLC6iiodQ2LAX7wVeKNCfSHAYc3/ZFs6UBbc8Wa7dxBvMbn0FIEns8KB/0v+9f
HFx09jABh6qOHDE14N+BnzKTvaKYY2uvQeHDX5EzYyHDjWL3dWlGPziimwFL0xq5dn7nVAI3+oaK
1GeqFy8/vgGJ1xmitjy0FafnN5VYxZILxxUF9mSR38bOHsnCbaN1ymXj1m0c/6CxEaHvG4cW8csi
amKRURD8xG7I2AMwJ8tlENM48wUuM1xKVDqsXLjMtBj/KUFVceEO8Gp7KFcTGNLP1tIJdud3OrLe
u+rlKuC8rym3BniM0bQ9kMtGdYKfVqviHVTmBki1oBoTsJCBPHLVmpfmSQF1tQfxfNYCAze0vD49
y38vKqlz2zDA6iq7pFMbiAnNPprzWAMSbBUX+jEmbHkQeiRj0Lifg5AYphlx2wrQB9dvsEl9hMdU
c7GKJa1NtoqkadErS+1El76TZsSeWK9FTyU3OsVBTsSukElcGdK+4LI8P2+YCV5lQrrEgipZ09Wg
pB76DrIuqwGiLqR/NVocy6YKax4Mv/R7lsMAAct7bCDMhQTeScCa5Je4HvI4C7qsLZBI+0o+SwR+
zvv1DxY2kIX7xMi/lWYyvn3BegbKCHMhuYv2Z54abfImsVBm1ki6qT0IGs7DsqTZ2kXsMCitn7Yd
oguzWgvf9+8QNaua5d7nz+vWuzVRfg6PvSEa2jlrV8eCRo5gl5CtIH4QeoncJ9uMLE0lhxsqAAwP
e2orge0FhBKmrKKdPTPUQY2v21WPrtwZHvFISbBLlnLaArK//3K2OLLOkyKT1jmhmfGU0CzGporJ
BHNTIA+flhC7aSSPTJLMbx1h0IPDP5p1zoL1l45++WpI1wBkJBX/CZiT0z20UcwX74bumZoxg/Ek
zFe0oSOkdknMR9D8ICd3SPnme6BdMy0qby/77UIDE2W93svYIh1nTYMx4LQQ/+mGNcBHvaFSjsCi
Zs5tfLUqPzd7Q1po2uDc1R6odUurxmMoIg4rS2L8hWO12XRi1a//HxTiMRRoAri3BlrWDE0G11ad
qD1ioyfo0ti3EkD9PeCzIQcZ0oF6Wb9OKIejBO/eWBIy5k+yHabq6jedrPOVhIZmeZBcyhVyCoY1
s8m35v0YD3D3PV3cq9mNxaAmwdDzVBku9YE+YifgWC4FF2jzBqZt5xxybf/SqgOEPjY+CrCeobs4
m6I9hRHqOMwgURW9cI24SbF1spD2Hjq0XiIiZ9KjRLrlLhoFjtfqhLrvwj8BUIa7d2DzVB4rKNoa
N5QZeuPzYGxkTcRQxGzmhbqJgRh1an85g+xpwady4Dkh9KeqAsYzeOSvd0euKXj/AvivxXArsYXO
qaI97pg8Xge+jBUZI+gHg0MgdK8OnKDxP6viEUumY86kcn2t/U/Yxg6tRIVdPCDIOvNp72iTrML/
xKyLOwaWHbgEYiefgJUBEw9OCZq2vRXZgMFW9MEhlSa7cVhQbnbUl8IUOgw31eknl1NM2BprAtZR
RJZXzuFB2RkVMnzqi5TyjBoXkuOFT0Fq5Js02vDr1uogOTvePLXPWHXkRZUnKTk9UT2wpxS8tbG5
lqtpS+1RoJ+SInkYEvROfndiJrcC8a04cuqoHxh3EtjB2lUgvZ2TaUU+jKSYdvQmh7LRP1K59MUn
qa73znpbve1VeAf0jOugUC9GQfjG2+hAGIQKVBpoZAUl5iOpH2c2ELCpaQr6zSm6ANVdfX7goC0F
m5zbWLr7/BmlcsgdhNZoJo5XvqLcNC3pqVEQx4apUG2YwcU8SnnbR6U9MIo22czyfAV43uRTI0ME
fZ6njgSKflTz74M9odbr4RiS5o56/Cv2CM6BSMnoXOtWcKN1kWaEvF1+G5T63Y9l88b1DN/jzS95
2g6ta/j1LuYXLeZVYKXsKDNU/YTxtQ+3jxNOlJs+v2/aJxeRlGOl6ywSQtv9J0SVetrRZOgemwkr
8VxTixDwJN8E56cBa3pPTEugMj49qbJcXY9W1MfGWZZHg1xQgF8LHytYrANp3zKKxrDhp8Ppk520
63T5rZOWU8cBQcBPRODIttRLktd68cf2dEzV7h3wjwma7mYnkbWCYW8UC8qnZ+FknyD9dTAQ/u90
xzdKopf99+TRqw2ZTnvg15hLHiqiuysHbwFmhkTZrRq0WzIHUG7Ef6pL1gIQRjMtYinZx1wcmLys
4SceQsAsRYkBS9CLvx9raw9N6jNk+txQNHPwm5hUMUWyNuz8kxVnXbRbWrqNp9FsV30tif/yp0hK
GdAX8KcH1E+/ZnFlU5Hcuxfw80RoBnTZe+EhNe88GveI96tMVNkdDeFLvAbRjiXbmaYxISABK38b
31h0VRY7pxRJL1JhLXT0NcttlSO64luiQdE3N01GCIeKYKdruq1Y3mxr43kh2gLPI5rmMslBdAY8
lca6Gk2Za5IgtW7r4CWBRRSpaINUNA8BRFPuAC4QTfFEUO+b2+caA8xPOI3lU+FdOvtQ2/3wYkdI
QA5fce4El1yXUq744P57cYP6GXdWeb4hzb/ndqoYD2uHeR5CrZHl9P0BGppZEG5QI0SCAKnyaZRQ
YKQyGiT6ml/imFYMadIM8SDLl1pykZ125dx5xhtdJqhT5zDaN7nwRlpmZpTqKF3KrHzkxRqfAOhJ
sdDEHT/AQjrx+0aXL/dcfJi3Q0a5MyBhTa2UgLPjtazRgdzUSB3jV2VVas+YTIBKNp9euweVrB+7
rJcbIcKn8LgCDeVitFV00D7f4nUZcy5p3+ZhRuFIMEsxQn7CGWY0GOD0iazWWsOXq+NBEl++wHnS
pUI8xDC72ui2JVHXi/QRI3YJ1+i79BaSqkrpsNlKE9yNI5Y2i4EAZMDVDYTkV8z9LTLQTf2fator
LQDrHP9FQq+1hATlCYmFa+I6QxDGWGNaRGYWLfCCUb1rDjj4MvXCdZrGZHrJsdk68SHEfdrRH4iK
sEXW9ingPQ8j6bGwOhwXWftydHs7Zm5Wb5T0KseT4WMIWs5xV8nNtWz3aQM4Oulcc/K3J7XR7rP1
57klWvqAXvY8Fj+KcC+Z/GnlRvDUwLwYx5RdQaXaXHIUu8f7NTjaQ4De4j7fZPDzKKeHYPgBvZAV
EXRkqFd6aay1CPFIpmzLt6G2XVIw1XvHxkVTJSPFilXGpem+6j1nF/g3nqmg2JIJUqzeIZ4Z8c2A
eE9l598ZUYCCvKKIbXufmeE1HoRe2YelWQDHEhEh6T184d1mQ4w+OCBlUkOBuae1pGWE9Ye33mjr
4MM8KRnyvViNVNQ+BVw7kPVcSxLzYdWxqO/WZuJbISmacptrFQhWiBiK0BXaj7+fSeJ1c1kmuEFJ
EffDumq+CJwEihC0VhjdMSDZ0sE1RPs/+wb3JGRk3iq/fh/zkjV3c7AGLZc9EihTr9axXcp1R1Ls
/6SP0BSnT3fD/LHM4YdlMPOWa0NsSdIGqBAZDEcm6KpfjQgMCZRCV+YAvO3/8JVSpkmZA1QvpRiN
vX86sKXdXd1C/dnXRaIpqQ2RmrFkS1V4WCLafMVX9YeDmLyHEQ6QsWnPbPjZZQptZ/1ZiE07+6xD
Xk+EmwDBxvWlMpzsV4M4ebBb5NUPyfr3NpbGi0whohPT4HpWwoLiWSihGr5P/EtRodZCpW7NrJKd
VmGK3NtP1UfMnTK9mie4F4xvEjz0HG7sttuYmVn28CrIj+5UchDczCMJNC+CYIwoZnJxicHdjpHe
wM4MxT48+J/jUrtuF0uXE7HIZffKishvNznQZRBXprbrwCtxvjs972y3nR8QH7Fy7ko0b+ip324i
BjwpLkhIhl+MFfCJeV2NvpLJgPh5evpbPEx7RiLg2joiBxjPLr8nyECtY6ALhC+FYlozb/LuCcEu
OpS2STanMc+UstrbgNR3Mk3JDyUD2PmZWU2g65Cg5o8vHq3OGYuCeFG79PXC73Hkc07R4JM/h8mH
WNuNkV5BrcGEJyWfhZKDe96wiRLTG66WhRZ2YCHrvZLh0lnzXMVqhGLL6oBVGJ3HT0jYpJ8jsFq7
xOhOMtsBkgsBKXK6Efsg0E9lNdJeOb6vrqW8Vyv+0+6Tj838W4udcBnQ/yj4GtTP/6wwKu73mD3/
Co2TUmTv0sj3tVpPW6SGWvdQHIEi88Ms9Q9XdoiMymNkl/rtMUdp4qbvF/+bLpAIwpopTeMhTGMU
WRJClyTLsTu95pSsIYcFwEo5CMOaSi8qVE4xZasf/wyAqVWjg/4MDrisTjUz3OkGyHxLI2AsXNta
IotEGXs1gQYGrm99xNTviVFWyrJWphkKfryoxIstgUkFv3us1dPUbjghzZWCxG7fWJTqeosStlBa
8NAqVwlQozhDl/XzAXHfrTviQvw/+MCmDYP6jLM+9SDGnLopUOvHS0SXmHhCy9ts1hZfsVevEOEB
cgKUE+Uys9cdfSy4hqgNba6jJr8VbM6i0c5sbfgpciw3aa5bYkitJs8mNmfNk+33d0cpvwvaNxg2
opodDPzL4nvNAqfD+22A1umL8BZ58mbFsebD5lZ3IdOWHVQoMPWAPbZLhY3XgCK+oIijkUZHs2bT
NwceLVBhKDEf4ZNTCCVYoFbZq0uQ0OcePLUggxjPNo3Ep3AoSu3yR8N/t9nRTYQepz4IMn/gXUUY
8DSaR/Ba4EnemIbcPI1WxwEY4Twur7WM9j/aUxQwhm5S+xxYQfSn74LHNwivL1h+9B3kG1s3tTyo
yCn/41rO1Y/gla0VhFksNpF0S2hWtrWB8cjrFrkgSogS4hOMIs3yDPBCpoI0aV1UoNVIgSIbaad0
iBp23Dk7rhYTaJ76lNoR1dTsGKdZXWNlHX4u3DXQQbc2Jx/HuzeSjnkDXpqTjRl+TAsgDRYSEUmf
XUgdGdJKpl8inDZUkE/L0p9D+NoIdA9rca8IjFCLyPtJb3Op7jV4zLGOwcTc0dwb+smcpNUU2zIl
pL25Zf/IMMPnnaJC7C6vly3prv4Oru2atfiOMKCqC4h8eSLXSqq+vuYkgI3olcPCJUMpjlRMpeR0
+30AI1ZUVNU0GW63z1l4PAT0n+6suOqAeU/Zy7P2Bb6d6f3uumdJ8WK2+Tz3k42s/mO48syWnBVp
2p4pNKTQ6+W1L4WScNgI58hiXzSXSK/5RkwqCqMH47kT7Ln3tOLE5fuBHMAUPMJEwVLKGhuixKwG
cM1CxaaK2pLFizytupIL7x6a6lIDULTo5zfQlwFjhs6zGsp9p6gUsa3QbfGBYa0Xg80LNRPcZYF5
LKYHrYeB8AFjaU6t3Fu19nzwinSZx6Gs5ushegpkkg2x9Z1YIrlO2fVQs5NZgRwWzkhxaFx5dwLA
Z3iIeh53TVEcm/bAKnnhd+Z9YOvFSiZNGC6XUQRwzD0c0xMwpUwLwuNyVh9ZhPd20riRTwCPt68Y
0hxNPxLtYg2129U50FRLzSYObcF293Si7zg5o64YWCmvF5uOAtg6mF5lFJ1hlI7lKpmkEudQ7BKS
KVwOZ1bNcrPa9YUciqEARwfzJsBdsm1MJbPmX8VdZVBmYeO6qL3+oOcztl2pDoOa9fCjstzjPrSP
+M/kjIAch43Ag6oGtd3lfFMFeNFKw2nM0KY+99OPBGubtb0YjxrhahRJEw8C4sluDtNuHf7bK4lD
h7MX+YqcotD/uTs17T0h4GNmdiMG/9iCKYYEHt/VKOSdZfzxlX6zLTe/JZIJmShQOpzrC88owoRz
QnfnQHSBQD2J+TBmFPOMziaUcn2rwgs83msfVT0gvC+K8uysKLfAZVwP6MYN3d3WJdNV+ZqSQsaM
JCyirFb5zMML+uDaQ+3NtCndOBvdDPuw6A7eMU5n+9qcm0zxlxbhdQbZ1ZcIx//CQFEnW/aigBhJ
dxSJqt6eE+MZV8yF2H0oxEzJkm0wHvvTheWWu0NFrbixpm/RIvwIxE0ZTRDsh4IE/GW0EiCpAQAO
R+KTquolWsFv3fp96xcu45uoo5YOpHZ2yx3OBU1pmqG0ag76Fn5IIjxU31cXwh95lByhzBUETh1H
JozNJAPibb6o4uAuHZMc4N4USeBpkrzUwXGFBCR3FhUZLm7yP+fGVz4KEj6c0xvA1T0RFVfuiN9X
Wjr5sA33tCXlGnNm51F+jADqyYQkjpXLwBoOA2rGm0Ak9k22NIWFrx+Yz2QBRAxLBGxiGr6KUzaE
eIxa1Xo0AYCe5RLUPuIsfSoaok/6SrfjAa1mtbq8W6Pvzk2mtzJgyHLd66gHAes33EiN7kgmvM2Y
Ue7VdfSkzphdz6rz8K3sBHPAHLwHOo+KTbzCg0LqI92UT68SSj2KpEP+zqd0WQx9Z2Woyw4gSwT/
pGO+bsAfWJtZqiEbUdg/hRYsbUxI1vI12mMaFWyvHJZ4o9g791gcvuf01F6PtysaKfl+6h67S9nj
KkDqvM3L+0j8aFKutg7nPpcMpBWzhQYRGjnCYEHJgyoZr7U9QpXnjOWLOq6BMJ6hOJL3POsnW42J
xDrz6F9apVKKDiU+AA9ZVgj4vOXu+5B/xMQLaoyNbuwLa69M1tLXDVxI0bm4kU4vAps8IWShCMtd
D1HK6JRfRi2PfRwz/vjBk72HEQhSe8SoetnwKDu8iuxk/94VCM3utzSmoL+s+HBUzq1qcwLVRTV2
Ag2YYY+q6/eGLgsJouMgFQsN/Q/FkojkXHtEeIA44dmizQciOwD9WwvekCWC34Vdv4ZRclYELnd7
eQJsYDN6R66KP1rc5r/J5tUPvZfnDenLJJGW7U5SFA3yyIL7xdS0i5y/twmBkrzernNVQTnESIzX
OhZ0Pjor2k/PFimwjg/ImqjtkYIRAySkdqnDm2McaKSGd7Y/l6yYHli9Pu6WwqmW08IPFNbCDDfn
KpBQjbF17VrLcF6uVnA1z04gcpywaKkOqicZvQ+H9A1uIhaN5m9b6g6XjaidHotL4Ue0FuGw55Wj
LW2S7unU5SH/XMaO2Jd2+KTtlVoilb6FKljp0yiFKGDyz3F97crA0M0IGnt7gkWIxYes6bIyovDL
RXhspjB+RYmrS4BK04RtzUyCi7UNmYDULOElZZgA8GhD+BEnS4wuzmJk6HKx7R61VFOOt1ZAi8KN
I21FHUmmwodJRnoe68avnjfxNLNb2PYwhuSCS5/ZJz9qncT03jpQUmjTkMF2bVVekCAqh8joUU1q
6e77Pk3ayyrfWpDStD/Jch4WqvmKlCCDgp4UMFtDnRG1MlT5C52YJH8XBzjI/yTu1+jR9xlAfhzo
OuA6g5LpN8HXuyeC73layGzPtJK0iUxePNmDMHbc8UsZs8JA/NFyt0d2AjxgRWnZOnQ5e1S8eRss
KNsVGeTozdk988d2OxueH+6ANd+7UgiqbPU2lBqZB3qjWCP/vI/RbFD9aUwo+jfxV/xLXBQ5a/zh
uDvv3uLkATvB/Lpi8GrmyoOJxwZT38ItgbqNdoU3Mc++wjY4gFRQ6X7J9poYytnre8iPtJkUdtGl
4Ff/kAbqdb+whZL59ZLBacwh0TvRySCx7IxfrtMb8Ul6JIBwLexe7QQ4osv6eeWzpGgQzpTqPHlX
Pym7quuzK/+fHEeJ4KjQH5myV5J37D+YibU9MVwjbi/BEcEHuW2os8nxQFV7QSSfMe2wwkhPPoH1
MBFFZ2ItfTICOTJc6cjJztQas4BiEKk1zNWa+dfBu00ZAKEOvOAnq4kWMgbW/+TiMbA6yxvze4fA
KncgfF0+xi21pyMQe4wh9Wr7G1dT0pLe75rBNzUFrvAzhAGBYpgVDNuwf7gJ0pm3nTeKSr0/fYqg
6+OZnWJiOLX+iMt7rjETSzPuDPpXqMOjjL1zHNbKu1W5hPbrHXXWRRqhhTsbM1iLltK1WzRBqDpY
O3zScfXLZIl6GuGN7fEhL4SiZSw9hJotwBg4iyCbnFvEglRC6bRFx7CURmq1MkjenmxK/B5TbDbg
FTIhS8kNe3M0PR8Qggs5HLj/ng/Zbec59WCAQPjNASnOOd+SqtO56TbZNIlCTDGjHch+RSDasziK
TCaYNOt9sxzCqno//90ACo9Hgu8LirdjyF65WP7jM2zidnQ/qMJaHVfDUlOEulVmsxExRQnynB3i
4Tno2WgQj99E2fPX6CmrZPfoRkO86yAgyleveK7ywQZz6p+We6DXT+/eLePip/IgBL60Fyn08fzr
ZWM/iKHtmym2a75MVzlRUI+0w4Tx76wKw00ZtKaQ4j1v/b7hjahHxkQi5PeyzuPUtKZum6HfAXv/
42RA2wjbfJgW6ouF7BSpEaf0QQAybPO21jNx6+PWG3zgC5pEg1gGl+48rrKYugv/+KIgOLf6GtGZ
Nw+GcRnjWWYSrNfJXqkw4VibekXTfDLn2wHWXt3TDULc02VkP9z38+4IX+aJLR0bkcCxmqwXetL1
am/CndRR4Vh6bl/nCHYRryO80isg0LEBn7rxudEu4dNNkihwBRAP4BkxYFb8A+wlia0twjS8cvu3
M0AOYp/P8cSwAthIzg3qjUUis1XK5sAd02V8OoCxuWCfZm1e2uhytlYoxcm7PfRySaIJqp9NTlqH
CGLenzZxrY0Yw0aw7xs2WfhXkxW5eFkyIsBsLWKyNVT+HX/1agKcedCcOgUgMRVFSly23vbJPBaz
dUeZfZFG5gmo5LkvQdDj2+Xh18+Sk8hG/uJTrXYRIT/32+/i3SNW/jBIIg8q0arqqZzBDOF7iR3t
FND/X7gsS14QDtyYRuhfABcSV0N4A0s0H2JbACUZGfbCVSLrhywIMOPPSVOny/5F//VVy1bNldW9
+Q1+lm2NQ1FozXXLwbOQr7ZtSkgU2Mb8iZ1xh3XiZ0eaJoxUlBoU2t14/KpxiHUWfZXLqHF2ZhV5
rU6nsp93MS95FD5P1jR1SeRLVed8CIqDGDPWc2MrBg15+b3JLgzfIPZiAlurM2f1Tm2hjICElIE6
ZNDBt7ymge/9Be9fch2zkkMVA67WmmiBjzUR3J4Sxjcz6HDtb31abKjx9l6DT2LsSbx04FgPVM3L
3c6lh8HIyMS0dW9Gcbq+nbMVmI12runMABD/wF+4FX7ukJ5Jd0sLwl/3Fq+uTK7lcfrXVwBlNu38
ZYCOvlqVe/Fs6KTeoiMIRXyD5t42j4lM6jh+nqqXNMIjbdVxa9oIya5drCi3wzaXlVFerYDXjiyT
oCcHCbkXrWF0s4hdl0lmsQZ0lvYt1QsOOvaXBq6YKaO2JSTvw1hAB4JCdKnXWc73fLvL8RVS2HOu
D44oYtS78XIQxSb5YRFQyn01J+ELYnLVc1CdUgI4ykOCJE2/qBoxZ0Ydmx0oWD5YLcbIVqqCD5vV
i6JBrz5cCfExjPgBmxeGCqE11Mc13PmeQlRIQ1ty0innY5IOLbH8YWdmemDgTRE+WWrbMBNgdcKb
nQXPVubJkKT03LDQ59QkY74/pR7/DYEe9UT8t1QwHFYJdpa1d9QmVSMOsyceC2T48Yg0/qo+BKX/
CcyrUkk3KEVWuOJn5FdlgXLutoXKlE1zEoNrtAzjHy+TooNWsSsMPTeiFvlSYn6K/MwHie+pzmy+
25poEtbsuoEIKT0W9ordndwm6yXlO9/qq+hYVoskJM6dfME9zMP3wH9wCTUB/jgOpcyeh2IVzLhd
/nkqjunCaq3v8lnofGcx+wJ9H/g1Bjt7JjBqZipfZFMw2VoWb8MxiIUuIXXGZY3sDXsoSfq5Vhcc
iF9FdBx/w3mxUPAxAJ8A5qwcCyEwwSlfzfOWqB1WknLwZBbKLjMu0/Jf1D/8lqnSiMeX5Sh4zVmC
0Yr7Ukn7HulaS0Kh4MG+L5zEPIvvAZvrc0o8ooFGRHb6cD4ph0Dmf6OfBsQpy5gnp4BzJnZFaiNR
WKUQ4utpkpdGEaWY/dUyjTpR3xyVoApih9q7M2GVnhrTNnmzlu6wotbpq2k+WO6P7x52OiyCQPNX
DSxXB8s8FmxL9Vl/s6NFWponiFGNdXuOrUubNvyRLHjTF57E2ILbVAIS7oLLikS2E0iHLxzcjqkL
PUT0+s/ME/R2j8AdfL7rk2FtFK4KKsncoQ8cE7zS9llxLpWg/Kuax7vH8bhz4Z/PuFhgmuhamsIn
XwspdYvQtiRcwu8DHDZqAYkKQguutrYA5eRvJlhB80K0UWvnUfppDzKKJzFbKqXZpeuPkvAuNjqU
Nc6xR0iv4b8T0J5ewIf99QID4b/SDXlpH6YWQcIxnNuThY8Qseq0lYiGNej3a0rPHJHKB63Hessg
9zJ0djuT0imIao5Sd9pSvXiRf5H/lWjTR+MeiwNszZCpClrtVuqQszJIGfR0CUCsBd2NQzcOTgDp
AVonDKW3tduQRzZXE9UNUdKMIk98Bh6zDqeY/k43U90rXOhJgCgg3o/0vEnuaiSnn/m83U6B3Z+N
Mh6nfDbsUzdacVbB8ylfe7TPw9+2dM/bg5KJMTeYsqK/TeWoZEIJWwg9fud78Or097g5qfyd/wc2
fh69dQWmWRwamLE2+yiv7v7Z2jWsI1S7NZcaRUkYW/uFdqEWsT6AmK44jtIKlsb4+igin7VuNKVX
FYk7pi8AK5Hw2ogs7kq/CUi9Ge+mhf8eaItsRTXa0k1yr4ScdX9AHGTtVTdBADiM3ZSsQyGgiMaI
2/Mvs6fh+H1TRaIK+Xal4fw8N16t5xQ22CFY3Crfa6A2XdW7DvZeWblDsPozxYebYrya+uLvxaTW
5EypWv5I5Wa/QSfuVgYT1BXJBmEjd85D2OFR6VzPV6zz/Uh5a30g+v9TBOFF1hwN0Pcfo1qBtQkf
7Y/+7m4YvoOr5wGaO7p/NxoqJw8G+002mIcoMyY3EMMadxJeLN7JaFdn29G98QF6kl8zXD51YThf
ibr+tDPiacZJecPHiAN2Dmj1sW8LaOHg/jjvzx6nH1N4MDMjqBRKde7UEneALFlcwBfdOMq1Dc5I
GIx76ZOfalhc5EzgWrbffDev+9JA7NgWQ8nAWQmR0OOpTlymaSRIun/vTUDFEEBVJt0Z2aDAOgEu
+S2p5XfCmCBUpOYRoo5r8895mYMmN3dReUZVE/6fnx5J0fL/U5eG0Zru4L1Z3NJoLC2bzeXIBlXz
QSnhNrWC3CK7tVIdOKnWl4gprWQIq4DT0EKRJ9xqYgT5n6rJiuzUgwV8vMFVoVgyr3G8UohKf1Sf
omTUHwu16IPBoDXA2ryBZRD6/jEuoRbnZ1X2OfXCp5dfjVOznbQFYPJNDeSs4AnRzQPZXYpDYw1y
b9IuTx+HrlkyALLta0At11KzVUBeE7lTPIqP4hyJ96KOrfLXLsw6zmFylZxAbkD8+cQrqXGmfYFo
KX2hbyvTt9HdJLB4kjZnURhq/5xtCiyMEcu+WfsFCiLYZtfvFzJrbQ7hXNJj2An07TRQJGPq8ZzO
RXsf7sN2OBwVVNInXh2aHL5YT4Jl/FNOBVqF2RFmytLlYTGe1HT+pNfdhcD8pSV25YXLV1UZQzMd
S/kFE6/4UC2PKDiDdGVBgTmv9iD9UTUw0DJIKwTGO34s5nSLhHPUBc5nzRQYgSRsyyENcUgA4aEX
qb9T4L6qgFXC4jciAYrcs9zJ2EkWmug09IlwK6Q7+1GIHKuLRrqg4jEknY6WfDDbhFkBElCumkD1
Y60dFSfgDY6WbqN5ix4b/92ICdzMmZRnnki5kOz9gELPaWCpmIMu4/qOMlVj9gtrwVMEdSm3TGP0
oyrFpz9YE5oipK6S2zJkO1HFTjxe6oo02QBQVECZLyM2s7NIYbYp9+jXiMKwwl1ybTWi7KjbU/ch
1GI0t5qBsbNig4D6HhNg311CTABYJ/KKmLQwrAI8Q92Y2e0zISkkmYka3UD4aPoDwxaqhbM8kceY
nz6QJIFmovg+Jml10xQosmExFuAGCqDKwLcLWZ1UbQURHgFZhVg3vM9cEEiOPJZzk/dQM78e5aqt
hJI0HJ8FbeGj7OXwwb2G/c1pU1Q4p3U3tGvllRf68EkyWij7HH8T9o2xhsHLnXPQGlfwpL1B+/Dc
KvlDgeiyThxSDkgZbgXgDrhcO93t2mo555Qd7g7aGquJJcyQTNlUAEND4h+IanR0Xg7tXRKQ9qIz
omZblYTmSSdaACf0B3m9Wo5pK5Rv0z+U+lV0CJH/iG4ziVc+wzM8WHoBHHNylhLyii/zwBkQ982L
I79DK4uozZfi0NbMGurEUUc+rn8G1qnDrUq2wVL6308iamiUIKz9TT2WffJGW8uu/nb2muCvrfq/
zuSgGlWNGLe82vpzKDHxhTHua/NT5/tItB/6su5UfxA6muCuPtW9bV75KmeJYMQVJ02LZulxWFJ7
uJ6cFvWOGuNG1NFQSHS4pCIMaNB3EierW1xY8CY+00F8CWGq7a+FMFaZDCLPHGMiHJCsg90u+fhM
kAU+3HmUiWb8PDZUtFqR9gsTcUUGOf4dgCGRJ++90QHYKd+eIKu15zL41WAAYVCeUlTKTV/3eHGm
8xxtGP9Tj5fXXkgrs2qYyTZt3lZipYrSRm2iSnA1lYUE1q5+tj7zNyOqDXnUikdWXdi+4JdWWwsW
NniJ5RjozPncgfjCM41KmIRAr5OfKocUTJcVB6xSuRBM+OOZq7kMDACx59bJ1NsLFX12n6Ca2gt2
92fc19tn/YrmZIRCCCV8e8d3xaRwqObzDdxUCLVbvjY2a/adBnKfimxnYKENh6WAZR1aCI211J6i
Bt43JSDuLxMG3Q4ciKJA2ort2TNtEWaB1F/vLaLrGPProdKh3rFu1kLCxTG02tO9pzrBAW0pfE16
mBUMJWULh9z9LXmvjzWn/7tcnYUwLugsNqsnr9wOrZ+AkHqdBYcMtvEi3DQD7tjTbbua4Pjjsl6f
EpIV8qf6YbzSxXLpe9J+FR+I8bbkzoE2tl3wIPtSBhKAHPxgFPVy8dFtK8yCIKfofV8h9kX8UJaS
kCeCyggjgzcBPk3VnBEDbyXoWvwiG1U6GTyyHBgQYycRRo+Zx1Vb3x+2Zh5TRfn7YV37anZ37Mcn
Xg518UG+7RqB/ae4KdpxRgzJjY2aRKCDy7wl8kWuIhUQgMj4wjPt0ABeGHKBQFN8ra/mqkYNPWvX
h+av7o1AeDfzdK7GTiVSkOejLjSEM2pHncNoMJtiynqEMyeopvAPKCs+2h5Vdz6SXq6MoVrHGa7S
OUCq97Fm17X8OZij9RbwOthgzi0K19C74nETFIechJDBSVaB/0hfJ1Z51pWNzXDoClkhqWPRdEG1
anfTJ9wzSLMX4BvIrFyPmIEcNEnuJoka6O/VMWLA1txw1BvaYOGYlid+KRZKPkz9UWeEh8iTLW5T
mNB5DuScpbvRdmJ1hIbuNIwAMz1to61kCRD8WImw7SPWrT5WxWcRdv9ddKWiHYSlI2aoGjmiELI2
sWyEKk3bXw5zXTyZn6MiO6NV7NyovHgG/EpRufmAO4Ng8QewFO0FvWTpIcLJAPlX1CszwQGqF/Ni
pBWLQaQ3aQtxsXvVoP3KTBTaA1/Lh/ZKDkng4RYEKAVZyNci/EA/Mz9GuApsUGilhKs/VH/WEbZm
bNXH4r4iq71QN6P2dGOppMKhgd1Mxl2ntc1VKblrbmf4ccha4Gxe4CLXIk2llR5l5v8IiwCMdHj4
on8p1VKkdtQwnYzVuINKUV6fTHQM9QO/euAuCU7MCvZ9JYiDcqvnUT6D5ihXysZ6bBf5Zscxw8s0
LNOD6WKM15mhs41/j7vf5XfNcOqbAQIKG2H4NHSNM/8PEeBhMHO9AVvAFVUeYSKiVhxO8OFhW5Jw
/LyZ9FL/4SpVqKTkI46umW+KsA8QdSjfoWzSi1NYADjab+iCoQcNLk7ht1f9ik7n+4Eo5nFyiA63
vhN2qwKSuIyC15GSFO4e0EsRWjsMB3KDYlunbJvu8Ml09jECqLsWRMXSkllzajEAfwAROLjewUBp
iYhSt/4PoWjFT0+JMxyY7VzW/8TOH1OoXHxHaQZ8HknWJjgq3wWAicQZQqACJH3244pzfdTdokB0
Q6/ni1MA1exCbzYwkJctNMzZnV0oy1AcI9O7pPNN+vJw5ePtqgZxCsSOqoe65IA/JVNQYgCm/IU4
eDVpNXyJZv0a+nHcgZXGgTQG5PHNL1FDVPt63bVeU02CRouQYxt6ALQ0Mwo3gS7rrizwNopFVfcb
AYqBfu7f5nYmHvoJm4qOEK2ffh+RewHh43XAiitqiM5VnzaFi6YcPX0Q9Cw6e4TxnxMXxrclbmHG
+MeZdKBSq5gmOosI2wLEZ7IVfBm5KTTffnlywZN0QHdEEmf2hNdbeZFo3O2XFlqzhJGZlWIMJ578
eWcW78aOhxWD2vFaduFbTZziFVv75HcKrRTJsFGZ5sNLYgNsyj+EhyqSVVuh1pFo2PeQqGSyXHzQ
BrhyUI+be39m3Da60oxJS7+IcaULo4rybPKi/9ZWtOZToDYVXbaIeSJPDsddxw4kbIo0cvFBWRcw
69RtUd3UTYQXfhRFvSw2uHwuNWIGI0T9pDHMSiRb7LQ3PaSjaLkjIsBpWFxD5TL4woHcbK4svNox
0VAG9OGrBJRdDKiAulxJA7zNK86HmWAh+7AlSKYLK3BWdE1kthhJiLJzNZe9G3vn0wzi0/fZ8Nqp
VZspwugyTe5M64bJnci5aVjiGIvGaoEWekTw2YdAX9OX0CVlOHvKTmDAFgPRKQdstCB4AQ4sMjuN
bMgqC0EIbW7rNI1bKZ/kUSUJpH5fTZxl3NaFmQZ4kmcIdpcVxoHLYpU2XKBPJnD/CJLGkFc0OSGs
1CNxFZFJjTCzDHwDLvc9Y71w1vJaCKGrSKI7qk0U63ApOag6SNWz9XNcXXSHuadoqHYG1T9EAf9Z
1O98euTRLbngxx18XADokDh+DIE6stb7VGuSDCF60B57gR9Y3oxgvR84VpD7dDxN2s8kmNvV8zFi
Mxki7WChNEN4h1tMb07+ZSidwB58YJrGEas1S/DKINki6dMdGLhs5WKKSLe7viPo7QtKpNPq/voQ
IW7r+nhLYBt8tMbCA+kBFl31Kr3r73MTvaZ0T1TgcrHiW9shKGngSwT7JmCepbnNB4VBj0fsOuzb
haRuY7vDtNhkObWtN01ZKwO95UD3wobRkFUe1IFIXMNOpK+nCLJT+P3TbW1jw+7gJA4uZitI8aI4
TUCFrWvrDjcNHHQ9LCMlDcqrrUxi75LvU4t+xMDS/TcACzsGzgDwVk5IWQ8bUgltsavTZ5LVUJLk
MijL6ut4wjRPVpbE49eEeo5mL2rWJErvjH2c/dBq2A5anlqEcZCmrP9rFUsaTlNXC6lyzwHbHsZs
9/Vb2yFZeq3pAST3QnfjuYUOOeohXdtSjtNYgYHjy6HOosBORVzjOPM6Bomcj+K6pO/XVW/wxuSA
GsLV00Hf1VX8ulX4Ez1FC1TCwSgbVlCLgtz78VjiITOS67w8kmDykT+DVb6PznhugctvefPCxb+o
Hr7XRHVBAva3zF/fy6a01rstJvu+bs1+BCBD7jzBwtty/Zg0gSekcRR5o++gIPMnHYbYzXxbuW2J
9Jsoikvjm6oEJDSDezGGe7Q1OXTPTpvkxXVyR4JC6KeLn9dWAPLO/fymTTUvBeJkeAquChiRYRNg
BmS2Puo7hK8dbBEPfQbojaMxpz4xFC2Gy74CvLwxZVyRFEzvfRy1g0ENu9G20QCz2tPM4FJyzkd7
MWvTqZe9gV2w0Sug1MtXNFksSHV03RwfEwi1lIi3u18vGascmGxGfTee1t8ESBZVQBCKj6tGLsKJ
2J1qbDDvLk9kIww2C5YXAdFyCfg5MF9jCaxt8W+S9AGMRI2lUsbVFCxMU6d2XUfaEas9gx9oHjNG
KVUTyuupb+r+OfkCmOjdY5OYU9o1s5aJ2ug/t6+tOqOBpheTOsbZQ/nub+ZFagGKrBBLC6CauGT4
j/pEKZ3f7g0clArDXpv1V7nROwvDXZOLFRIaOntxOJMmdUJ6Hf9mFmvQ6VKeS2cZyHE9P/Y8OYGQ
Ozk/KLuqNoYff6PQv1nCyUdEGKYD08rP167cNjWmZ2WUdBoPIfUryUxbzuKBoJYCkfUU9q2VGEwp
+e1q/ENVoONWY6gptZjVUZkJRwQ/K+KNykcF0j/Dqy+A4gq9MQKZ+Xc/5TDVE8yFF/kvWMMqtwRo
Yd3GoNN0n22T2DyhmnXnIKsML2x5p8zLaVuSTifXeZMi20w+vDa0NsYMLiFJyHMLa9DSUrfC9cbe
tJLwVuRfdyhAQUxokvtEOo/Xh83YVf9KJD23DrnT9fqqkPqlq9e+RxqhBYRlnJ+ICAt5rgCXRbbQ
qz5r592ARaIN/KvIaMuIh9kSnEQg5ODBnkxA/oYf6295pXbmQy0Tkp1d3OwRq8T4Wkt8UzeS6ssw
jCmGHHJOAdu7wgbZIOOEcQzjvz8BlKu3lwMx1xEQp4uffejOQr6aRhM0DVYCoRAXc8Vd8eEZg/jt
p1I8iacpTEJ5vWeFmGUBDvXMjLHAhWb2O0Jjt1YKmwVmAYUhxckQpXJWhLWpQPadddP6IN0lsoMP
Ixpeh8Uh/KUKVUwwtoitBN0bJ5aTI9qy+NzuqpboeV4SBvyQuVHLbBjeOHwGk71pYzFSUugrlWJB
2aZn+nMXnlCi8tkJx6JTDhXV/wI+mkxcxcmQVlVdElygskHGhKllyzYTsjSPmfQUQDhSOP+F99KD
Dhl3xXP98YtPR6EMw+qFU7L49zi/kshKP03F0ziZNtFqgktqJvx1gInrP4rzQp0J6Yr3Oct5UZuv
o9R+lpF9OODUg9ogj0lNh4ZQG7MWwzkpx3AzoTJ/6HPniD32MwVpJYDXdXFYykN0f7XYfWJAhD9P
6TAZtzskQ5EEXKNAZn6tcJn+l43rQCvKTBJR2KiTnmdrb+7vEo2t9he+XYcBHctifXq8+V8koPKQ
Ifdln7I/EfgoMIRQSvJlTwwkapEQaov1w9vmjHtWkYMuOKvISe2eunbAYL+0K00wcg8XAmRKNolu
KGQqD1VYBjCjgMVAc2vV0w57EsJOidUOELwcS4vx1XUa9OG24M8FWy5mHrw0LMv9t2gxFK91f6o8
TqWdQtqo3hQ1Wrk1k+Ksa5KcIDV5zwFXHfRJ38VO2jCW006DmfrpSthvtud1OGA3ZlVK4k4gs2Rs
oHIIrujYgvDtxyt+woahQHnQo0mrg7Ho1zG1SaAeF0qkSyKTzpkzEdYY1yvD1KzShVbqsaAYrY6N
WBdc6GlIB1juwmzKF0KxXmdftBA9fYhfqVD6Eavx0UwOyYBz+f0mxOZZYYhRDT1LXtuZwtjPxJXd
nR170WfvpMr0xAZzQiQmIMc/BdlxgcumGmMadsefvIVTiQxwjLJn2cQ5AqRotIh6gAd+lvUSBdhz
FBqHXpWv/hPBSvuIQn7rBbWCUXyp5YycrKsNc8VdgWLchEv4ajF52dgR4yDuyFb2hxCX3DjZ573j
JMJpyjciwn4Fp+NxCEs5Vh0V/ez+UMz2px16n3iWyk+84cYSv11m+b72GvVagP/ZI4R7LuCg86z+
3aZ5v0x6UbxN1TjKiXYz4KWbkcNkDJ6yD2Ms5E5NsP4qfq3o2kvpSe70sy0/0WeM2jP35HKi8NDr
KeEMBtDH3hM7a/hNMnIM5PRbM5iR89UD4TKAQ9OXXJin7YPp5Gl3buR0jMd4G417IT4JpqlUNgW2
O6DprG8k2s5rp4ayQ1llHcDJCWH0YV0SzG/Tyzyg2noiHdoLmxi50XCem2+Ggqcoc0UGVqcYYCRU
O3nR600lKAMh/+PHvoW/m1bp0fw2n6emqUzd5uNOhV4eX11nyKup9VBzh6JkgGpGIW8d5zAjAE95
d3vf/ohXYTM32Hn8G0NT8bqjiJIk1LfShcnQOaxNxiKQe9DCPVaQAy0GprqCMQNInEl4K/zxmh4O
EbE7uQ5oduufPefbaQ6lM4ii4npmhGFccIzhR/tTGioQmEUA/1Mr9finDegIyM4+i8MtrFJe6QQb
kXFyAFnCChGTb8brA3OSdJpLJr3zlbkomsYCMSDXijAtPZJ1ZXzbvkba0LC9Sk9SU0V2w9QrFUcl
dMpbThCdmx7URqBfgsR+ltZe40xeSHZaJ0KdvnJFeNOAC9ulMDbtcCSJQBR3DDLKpkEetYhYIpgg
bORu2oMWqrQ4DryK46sdbeSURvxgq79CMApzegjQ6aUGTxXUyXVbWx4DH3wM1VL9VX8ro0wE5lAl
957S0F5w3Oq4TK4FrKZ6+AOwdf/AdTUKBebVk6fX2DVYpcrsOh2mtwmuZfNLEZIFYuIQxcIyV7rt
tWaCujlxraS6lBQHoXkUyL1piyaXzlczePeYn3venpzatBQ7QopokCcaNmL/srQqLr8jg6GFkX9Y
rhicj7VEhnGYoQMAPLfYue/fts4grBEMczD0Isl7/2izCBBfVhgoKsMDJzkHTngS3L7FWyna0JZu
9iRoWh2P8Zlj60nrV1ihW6Ciy51XndqGSA3uu5ku8oJNKBJjJmHa2pwDJ9UbLGRKoqK5Aomu3QVY
dVpxvmI+FIfGlJWuk0HHv/XzVHKlxhQpJvYFf6VyvE3cts56hr4woKyUbqqdM6E2uMxfePv3abS7
Tz40yK0XESuJjUIO6hdz3lU+HtUNdjbkWvEvUomxe8PQzEiNsTrGirjp9mVZIktpZh19lbgXVNrE
CsG7pqTCV/5vPm67wLIAmOR1BNJPhAhpuEtsCN8Bj0Rqq+cYq//PnxKWq/UmzjXmcdIPIl5iNE7G
QLEszwnZXEMyQzN2u0DfpFzaa41oJcFwGZyNR9cC4zNGVEOFeRkJ3JH5JBoy1AbcwgpiwY8qKK+v
b2wyERzS5NV+t6pb/an2IrUczIM8HStY1rlXI76Qn7oWznVGElKxVb0DsxhhGo9PUIR0bKiO61BP
Xcg/khS1k44PhKyOTchvnZJfo8Jt8SE9aCK+Kw5a6+G+qNHViJnDWpyH8lyShPTqcZ/zT1dEkrOQ
qI8PBuFG5fTKUYhB1xIwB+AJtynXPZbB48e1oeghX3gIL/cUfth/mf1UvL9wb8fFdqBp8MnCKUrs
iuSRd/dizZ7LAIlUkdB6RYEL+EXEUIZa+caUPzyd3KhXeI/uFlh9pwYq0JVkHDrtPfC4ZdJZq7eP
ZXcvuiaZs0uVQtFlYxan4hj51hEwJClMa+h7TiHSor3E2nYY6jRobW1zSPGh5H6Ny+99v0hexY07
NouqX3TQ6NZNda1xuU8tJgHQSPr3j5bXwtALO9hjWtLRVGBjLx5lq7uohx4vAc67E1/eNBl5+5MP
9hQKbF4HuxWk65XmIfmPNljX46LeBgSCvN+932XOdUhixGBlmXwW7Y/Z3h9i6aOgBMqaAJ0ZLxX1
JHQyHZifs8qHy6EJJUMrj/LJZ2C+lPhYL7MSLBhce8HkJBjeScqizVU5b+D7mkPNsnQkRBxsv3VU
7p7KL0qMR7w9k+My3ejKZw4gSuXyxUg2Z2aeSK35zZpoq7HUqBjodnEryY89rJkLX0E4SMVxHBn8
m4WSN3M0xJANabyxaNZZ+BGcUb38qcrAbRY1gD9s4nVNqdWvJVwPRMMuu0FEGgeJ8a1pJNN7nHFy
hqGpM0MVYC4ZMo0DGbjnnBnC0znbS4bx86GhJHQwfQyB4NSmnNxdEtK8JQmG2CJUZ5MapiRG+jsq
D4LMWrOaUxFgOPgovEOg+TvxcrIpZRB+7WWl79wRhufKkS/L2E3tAUN+ZD/pmuvitg6z35gliZYf
KjP+epCohv9AVGlJrSd+VkfEwkrL+Cs2ITLzdxKmw7Jiv+uGkZY0q1n7ESHHpAKQKSjegZs5Taey
F6gQnZtl0FDDWeeBWIpEZM+LfUBfjHPVkf4LyakHW5FjJYgMjWyg5CKWrLvbxT4JN9yhNk77RDuo
9xY6eWqqkamd1AT6CMOnBiXajCd2Ew2tUJ9RCPt5yc42DN0cA/P+IkFKGAAssvI/jM2M2nAeRhqX
18f9uKsShrTbLsQu0M1kR68eXBQHpw8Asrt5VCHuf9ZHfbn3Zz8nWpAVhKSHgouPD1TjQ8SDu6U7
XbaGBj4Lg5wZ6d1zevpOW/6mpB/8Izohu3TSOVHKXwZF5MZySudnWMPXlkVvPy4BHzmwQuD002xZ
lMzlSizYRjCCEFrjGHBHMHTdrUHjyBVUQdLq3DExkK1PhkITdS0OK3+KphLTCXnY1v65U0lAHFvZ
MST1Wdls1/s8CCiFHDGga65H1F0CGQV7XAIq+eHU5gXBUHrDECNJ7QO2E7HqWGn+Kvk1xgvK1YWu
ydfGHGt/cuI66uVWkVuFC7M0hN2DVlEV+56Vk/W9s3n1l+4QfrAuheSheTvMiErAjX5vHmh/AZCq
ltckuFep8BGzZ+LCYzhO5q5c0obpMPPR5oFZqYnXJNdXDNQ3+4B7Bo9usXy/wDFWxiuxAedjk6bg
mvM2yTfKQzKJqCRUQJAOscFNejpokX5x6yeh5snIDpeHHQoaLRf7ZUg7UnUmm9HPBxnXylrwPfpg
8DxijCZPSOYFFTeyGUrdADccH4RunmJyXs7hmdBg7FwiqZu7kKv66qpDw4P4GgSGhO0a1+CR4MGD
zkGdaGW8bCptRV+bcxVix9N3jCytMA0kQTjV9zW4uEN33CV27ziWFhm/Zfx7VvYh8A+72GZRsqf1
KWlOJmt7k+rPBTlcDwZdGTRbQNE6OrxZnnz4x2AcFnJie1CQ3To5zbBMeX6fxjQXd9irTCBDzlEt
xbkMCshJc0ccrs3nu+AXdEawtvgZTYKVRv6dEUY9xHn1Bvcjs/ZtNnIlisf1SfQB+Tc0MsgBtwFK
KvQIXiF0008J47K0YCiEfDYBTJJH7zJtyOq7yofhBBHUAQVQzPrsCMc/AYiQVC/lINWNZyy/T+ZJ
jDz1XmVbnRKULoNmseg6O73XyT8kPlQSaaRFVlvhVdpfqkGttst/LpzvEjoWnQictBL8gCq5/UWq
MJKkE1wS6TIcydw3wU+IJNaGGCs0FgkOlTKPJ+/fU1+pxf4vi3btr0hI4YrmRQ6Bg21jRgpSN4wX
gkBte28s6keq/r5lbgXqsvtV+sJASXreVjWcMeeYwSHlzy60xow2ZAp8DvNsuCPCnJwrLwS2K07E
5WcP1WWkSVG5Xx3KAlGeIkltuKtbOXkEca/FXUdlnnz/kleSu6FxuC6N4mLjlX7IIbkKqutFZxEL
KVDjL62Yj992tyVddx0kdnbBEzqxyMuxv1kCOCuR5tUesZ/q4kcUE6BqMKtvrvabIANFJRTHcmZ2
OCC7HMRuKCCGRNDQXtRaLKY7KMijoorllNe3/U3etTmjbey5qqZkAirCLFZLno+DIBNXch1iGI7M
OXGkTfQgj0AKZHLBpRvOGeWfQNiC+lAbl91D9T9yjY5ioQ7jLcygMCrMHJWNVhJx7w9jRMFqFFCT
pbnptNqDU8rgfUhA8O5aQElh54k+F5X/oMV6P9UzXGoRARVLJCtpYpZMzKAw81zyner9nXFnrw32
pGHZpryun3QVBOZBgwUXNqZn6qbjaqMZqzQCU0PTZEV9BEgAQk6a+rc9MCLiC6h/Vlha5yGaDRYM
L9nsCV2TKpfo+I6fAsItRSyRE7lRpQ/MdDVww1titIq+OPd8jfGrHZgi1SX88rgQBn64m37SlTBr
qKMxHEdzcHhjwbO+ON5Y1homRSgKnFqLh+0DKF/Ydb1sLVSH26CD7xRBCSMF21cwJiBrJOZmrpIe
wbEs85Z7lAteAsVnr6z52wz36mI0flcZWrHyRxJRI9tQIjiRGMNjG5wVf6Ib7rZopYqwqAr4Evx7
NhezFl7cmTwNk0vm7q0zBVJsdl7loVhCEMzG/yA+dqLq6mUmCUoYg1nsCqZY1ofvSxmLD9726RYU
8A38IRXsSkafScc6DD57nw+84OVzc4A2YEnqJ3tCuiNCK+F5iFdVhPFKbdnqdrVckhw+imw9TncM
L+BuPDbW7lZMf0tqfWJZcFAACeCVuZw+6KHAbP9UByCXh+0YjsbzGraArr5drLr1HzI0ZTd8pME7
L9OEc79ugqrmRBSqRpNdFVIs3rZnU8hR8ZuryscgFMtq9hUAonKHxeBiVEC2ZHyyAUVCqeOWB+p8
9qlZPIuUH6jQYxigWHjpDdOyJNA6sMfxqvuPkw5t0zVXyQ0UxZF5mUGKKeqpXExNHAcLSgLVI7PR
1cR+qBnBQJGZW+xkRW9Zk1EStvHpdtskCrnZxF0O20YhVj8JsWydrrzrvZFfTLUmyQ4ChvaTV7V5
AzUkXlvRjMkzfiKfurY/kVGssLNzvTd3YdqWFdPmdP9OQ46SX8y/GP+9UKicKZ2a5SCCm1TXRExY
9rDnlVr/Xt3wGfeULLZLaKr1nYH+GrOyzcin4wIZndcmgczrLc4adBP20AOifabsQb1qj3/aFA/D
QAdzkqg6EzP08BMb8UeETuxHygKm5UOZJGco5Uk3ibbBdksROKFMzPEQaH7tg6AiSurGAeKdHUxf
dY78U2FRUTzsXzpvo/OqHaUSN5W5YzmOncKcnWEfM9Ko+Zjw4Q80Jcgw9Xamn93XHxFL5bmZ4PBM
V6joHw0UO/cqFYz35QoiHDj3j3EtR0TbUP+jqYE7FXBqKbL4nR+iosdpS7xLNwKrDMGuMjr7l+2N
lTwgvHsxHo7IwIju9jX2W6I+SEbQeF69Etjk4y+HMENsm4IUrB7+de6ZwkXRsV/iZObvx9G4OXXw
Sio1avET+uEUWJNy/xSChLBN3T8EBcneRk+0FH1jvD3y4NgHYdGvgF9oorGMZIXUrE1Cv30N5Ok5
XiRxyp/bRpdkWyVJVuVzA7EhCd90rYhAJ2CKeSvotpXy2U+gNeq4rNqHWQZTsdm4yAM88ydO80eA
0ZqMRaUBjf3joqCy4kCEmuNxCEv7tyu/8SCCf7OT2Bgcl0mo+uB/m4nWbiC9993abFP7cDAfxZaX
JXCRuLNsX+BXnB+hU5lg8l24PUBSiyexOJBGPJI48YE92xGy4eXEmXa76JjRRlfhnhO9PhwAbWBI
WK2y1jC2VS7fzBxytMzlaoB7pcF0bBjkla9hklNMPlOQVjUhOVFE2EJWlO8hMWJ93kNA1VL3ox1T
9+FWnyiCU/n8MFC7BJtobDPa3MXXlsUQawWPmYgJ6CUKVnfMLjBxI3zPLvNqRnmEVpAJp3hiVLCc
rVAU6WExXnfvmgNJNcsnhx7XZp8y1UEQBbMbkubjKG80rPvL96bnOisOCQ3NNVzem0OGDrWpgXHj
eGLF+BsaL04/Pm/VcvMwT7eErKDgc/FbDo0kCeXGVsKJf515PVYd2MGWKnqhZClq+GreM8a1g4Bk
W2eKtkAeLJTbEUlRQo1Whdb6R9o2D4Qkx6hrQNoJwr1q9sdkgf5AuP97Vv65vQv4lzq/arhhT0xK
xdopH4rcL4ZdCQL2ksEgZCsIIvgNBc9J9zopPv45NKwfZ6M6wSa1DYfBtYgt1IS4lpvmf5Yx4CfF
ejc+puhVORFP8J0C9Xd8pPS7E2skWoRU1tp/hfjvORIe7mRdMUqdBxFaSmKvWjXpokBslAByGw3V
Vbgdnh10tYusYor7hF7aam9hocSEWy/gffBoa79NWj5sLWORKXahXV3FeSWyQLhkftK8zxtzKe0P
2nVOLXvUWsxyJ5kiKsrBvwvD8MSrCAM/V/7Xds2CYRq4GmlH/T+mnb03k1OR1AELt4sCdrdXQQvQ
+wjUYfh3+dn7uOy8uj3dG6pX0wt/cCjucN8smc46wu8RXQE3Qq0gXhXeZE4nxNaU5iEtTBox2Gi/
mwjw0FHMvEDmqMAXZhhrLutM6+z8/ifm9MrrgyMl13rfl9/8CYS8rGgrA/qxRUIjwBIrqmdbbYiZ
CBg1j0vd9DvRnEahTAWE6+SCMr1VkkpLHzIY9ZhwaV1JBvlbzBaqzDYzNNTH+VBaAI4xQqLxxgU4
60ms9T13z98Cw7mMP5tAEKq2vqRmy4In+WEGisiR3QBeWRiCMtHlormsLTWYwNdXiB0OHXN/DiwU
kK+nMejxoJVAs9zavDlm/Fr0GJP5/UVCTU84od6IeZA9FebUISgwQiAttyXbBy4vRBJFYKpXGVY+
lEaWYEYi2mSpssupkDW1NzQjDMYUvvrQYeqHLG0Kf1xhWXC9Snu3Q5VZ8XFa86LlUr1wqzAcItVJ
jGIl933UcpIXsY6xTvo5XS8VPgq6UouzDUL4CiprjLdEFIpjzhhi+lS/Vu9VaOGWXfFPQssZYEMj
2u/lzAmo5IqddNdumflF0eB/G9oMt3nYWqHUxgGOcMArZzJmE0VQbPAVwpkURrBRnK3j1i2Q8gOu
ytuGSySUblu42Ny1sJSwMV89YW1fh6xpf2BOJutM/vltKYcEiLf49fDe4+OdqqQv4ccxlGUr5YOB
IFWN9MbdLvru39oTNeBPp40aevou9SyxZ092Ln41J9JYPSg6SqXvMDWBdgkQReG62z7WtYrqk2nJ
7zU+QHgAk0Hw3opXmFYFfLclx/A2Hbhfxov3rVNf8ca4KmG+uQ5xV8mFjvpDkcyMzrLIec0SR+Zq
lJh5vjx09U/plG4nIHHJal+cXtjoAQ4VbHtly/BJ4+XhWYNSdu42HASSA5z2lagyiOts2I1E90iO
OGUKKqRZBFQvwjxekxuuC4zY72S0iajOgnGG9oDuakzRWfknD0AbNWcMpn+687LqoZIA/9J4xs7W
lZIgnbADJY33Dq6vz84vhullXFEfyQ5c0LgAb5qZfVORKTocdbnCCud8bCXlVePFTZ2dhv9csh6k
RVBlt+7Q5L0fWN1nbmAvRpoouLWGSMZmT65BCGBbDZ75Og01PR870Iy252sOuRfDsKWYl9mm1Kyj
0PulIR1yzseTvM31hZOWu91eJ06DbboM9dVlNxg9Uv7hZTwBlke050KiH8KLs//Fq+1Sdt75vU/1
0kl/yxWDCCSaQbliPDJkdRlL8toUDkGH2SGMZ2xt6zT/blwMES81xfCESomyM5dOBIWHsrvMnWfM
zR+YrBb6JsN4GpPW8+n3/h+ig0M555Jg4PMHP83GNlLbqd3MbgydphKHzmwbg8pqlY+MqkhNpR0V
7Wmv3TR1QTZaYGnZ0xVQpKY0lhSWTuD1ZSQWhCXm7UCaj6xm+QDtXhXUyJmRfu2zrtKDtm05bi7B
xXhwlPEnZq00s7tEDkJGZq8jqJRxi4e10KFNMAc/mUw+E9NYTP3TVbDZljq0T6hkSEL4ntMlyxeC
1Ib1+HeAJOYzmq4ruelajDIrN5Z7wYsYx9ToxkzZOOsYknsivT0J5NwC6i0HlP4aNx7py+1pl9eJ
gsjRo2E646odVbsR3Ix/HTZPZKQo0mUfoMl4aIR5Y2XKrjjFwN7yH8lxGeNiyF5rcUxW1ON73tmO
bcsAX8KdynUN38eyhuG0J0MSKoXD+GjQThQfcaxnF781GQJzgDvwwjN8xVQ7gNnVYH9RVBxwqFko
btTQNSvQNJmLeBy0hd1ypvFiaYDHBQtMdJ+sFHzAzgtJsOYXZXCtH4Blr3FQAGgW9QM/U5sfNkKr
yfV7eoOuRwxuSFhvwMIx36a7P/sjk/7Ob8AtYqec0wgeHtU5H0W9AsmsDbC2Olg9vG1mhCM/NDIm
oFMAbUS/hIbstwcIPMIh4+mQ2+wLmZsjFOsjKaLM7d35fAHMqy/S5dh0sc5h9zdETAGSroodbLS0
I1PWDcy4Mv3c+G/WY1KKUawK6kbqYYiKrGaU364N+xG3n/3w8GNGFGT6EZ0OuW5m8EQy/xabI8EK
wXIksUOKbRAID/ZGf0qdJyTFqkE1rCWD5O9/usDo+50lZzWP1dxleFLp/t4nU7P8fe3JQXGoHb6S
9PA3Zm0mSG9UeIaAirgDo1Ga48emSpukIGGcG6LRU1tnM/2nFasXVqXGyDn7ztqHfMbwLc8NOL0G
TSGddgM4oi7+o5GPNT4F404s90tqJ7ZbrJK+dDHxO1D/zsBUsn176/1x6hm2/k9Ymkl6Ntd6t9ZM
BXxO9vl1+DefWphJIdajBuPc8J37xNoacFduX7yUcp30eiguG8HdLJUKrWqO8aV0Dv5D+z7VCOg7
j9fY0SpkWLCm1+mrXFBieiQ+iUZmZOCSD5L/6c8Ov6BLFtkT1JBWIpXBYl9IF1JMCOT+1ll9qOG7
iO/AFxnDlUwsPbdBSBgJM4pgQbAQPnqSYwLUnLHJl72iNLv0iAAX6oWj+O+bEPgZWqEeIVsCn5+K
yLtvjIcZ7r6WJjNU8ZnKXmGZNa+ziNVdDXATMPfxtGXsB9k1d4s0GwVItdbnqF0E5D7xJNsO8T/2
15PkaNlUA6eFDiiIUrikPk+op8XR/R02ePjhHZflM+Vqv4OwsvOR9ZGKl0KuZgobusHfCtFiHwRQ
suPohs8xkfpTUR9rdieazCpBizAK2ayN71A6EF56nLVqGksodQZ0FdkibO8DDG05NRZYXHY183uA
/2AowZ4m/0Jq7IpjI4nZ1mE0O8bJhOavHq342NTdTqPg6P0mjbOZEZRD0vkAe8MViiyH+gMqTd0i
7U3ptr5ZKGOuZ4xbplSOddtmtjH5+xIw88SkDSPS3x+NH3y/xC4wFKLqQVGd1CrrmHfHsd9DTw7h
2oe1u89Zh+EUKtOofDUYDd+DqmEXxivyPw+VbS1GoJDrKZQqov3yn0CrbOEXvEtiRy6b1HQ2zr8+
sqB3D+88xMbOdrkWuNRTaGQ52FIg9CjvzrE0KZKatau0EPhSvfV1Oeejl8BbVdIi3fhQr/C45vNx
lpS5eEiMoR4xMwl74pVZ4FWSCBPJhQnavp+6IkXhRdBCVDB8zzUFL+33TfIeRCoHWh9t8gErzhQx
o+q8xlTvXmfcdIBXMmaCRV6AvSQrBBoPqVdfWDd1TLRKNrJGYooZlgIntu0yurJFeaMwV4LK5gb9
43nSZHDfw+Wp2Cb2sVfZA/QAP2QIwKMkACSgBKqfD32xGvjZmYIRtTsS3RwooISHvCeXhSYkzS30
Mm46aMWf0HJuidiLNkldvOtz39uGcIQDEdLsBa8m43M1dDZKzuw14q7o8ij+dN+AwPPAiJwP5dus
FUZmR8J6E4GiMkioE1FOKKPBYRmMNiE6Krlwac2RRpa020vIJWJOPI9QE4LZHn2JtkvjodgVK9Mk
13scenBPE/+n7WP+oUnHNZSUjy3uu+kakB0U6ZU4yHNC9abII1m/RgMjnDGiNd1MChPOm0wKAJ+d
SncgmBXBiB5AIbTfRLTsS9wK+KUpUiNNG/iG7sih2/Ulz85JBJpgYGUdr0jFxdLIhrz6vgUy6LRH
JzLVpM767bifICw6BIoa5cruH7NWi8Enj/LL16vz1dT4LYBqlXkhf8+i9xinI+Qm1nmJEv5JFsFa
Iy4Q0Furu+oDKf35peO6c7PIUuD0jGDPCIhw6AhDt220/SeV2TkdfRWLGqxRkAfjbpzW+Tg2v5ZS
8AEGzIP9kd9T1gzSLRa/NTOu83R39YfbmMrDNPaADGStvjs2VzAxFTnHTZwAjv3YLLXDcrzzbiua
xnbnKiEiE0PoXIso8xNoJEk4aNdEarLwPUo91oUXEbTSUkEi0lYwkhN8LJIqQNBBtMNmG3yY4tLv
7Y4mLoHXipI7J0NM8vi75+bED+Nqkk+A8tTMdDph845Ct0HIB6UAeUdUvpfmQFes1ixaqSU6Hcfb
t1C3RNS9JlEzSUyeOIP4+z9+zzSw2AlLLzdsRl6kbZIw+H4S9gGjM9psXzpVGbDv3Ad4JjGmW2QD
F0SRvislos+bZTJx9n+5Lwx37BSy2D5nswTFdWga7ZviFccY0bcKSsXXBM/EwKGiVKOOZ1pfkBdR
7l9jAKjY43PykVMbqOvw7vAfU2LOHXBTdQtwJ4MwxQ6e9UZgCzMqio9D+ipJLefDTTbki8h8iAeZ
KtPuefQzK4I4DnCeCk3iO7Qu6njQcCYpE+erEJ07P3r3kzMK4MB9nguF07NWHu2oGDBIl4sKYicz
cxuBiy6cqt91gLKfH7bzoniy2eRnmWOuh2Rxzsiq5xrP2cmNiJvvz8uKCzCu8ZS4Mv5YUGgeqqhg
M6ywwuOjP5tVaMKdof22xXDr+hu0Nr6/y8s2odSALJiPGJIuilXFO9lb+xkkkXQnlE3RaVMTq5NX
Sq1MuDl2DDumq6Wj/QMeVf0fqe0LR4aw0VXyvcFuueLknmmvLdMeovMuO3aBmQJXa996GionbPX+
1aYs2dYa+tXjfGGsNsR09OHTf+gsp4Dy+syLHkUKyVdqcZfi9wOKawSJCvRuihjSlVYhV2/g/GyL
oKYJ0A1clG6mZG4wOau28r1OCobir0aHlDvSyxvedYd9U3uo6veo49SqcjdCgFuRGqGiHkXaGqqX
5staKhutkWBhNnAL5HNxVC7h6rHgDenY9gYL8H9i8+JtlN9mEWzBTqrvkfVAx5yYo+9fbdk7h9PB
/b5GfFMVah+SDcIimZN/8bKMzUhA1+PH4kqL9OMU7d6ur6fmwkP5qx/R8dNJkK4gcVStufAbIteb
3W+WeN3UGItDAXwTfdF47OXrxa/1J8bC3xULkleYJD3RI7m73ejwY4AmCb6lDJwvG3Eddg6yIJSB
XNBl6CUzHzIZLmrypXv9nNadLNawVfgcx+L2N5LiglNVjyPw+Sy01d7MhAohi+Y0YvbfTyisVckc
yShoFm8xk2J/wcwDdNL2JJSbCbe5u13JBdZe4Jr6sHIXp1bOy1nZOgsVnnAn1aCF8Z9bSP4fj3Uy
SB4MMYhkU+W62zyN0oLC3MPRlttR+3jGIzrzpY8dvx9VnR5ajNBtKiZBKNA7y/IX1Sjr+tC2T7NJ
YYc2mG3EGoqhnXRTBXR3E5DNS0kitUVdzi0kE9kcv5UnSuVm3McyuuKSPxPsRJWcV5OC7ZG43eIE
rmIop74UK8pJtUEkSkn7AwGEgZZsUHgde+V+Ix7uZsdsmN4GcF3sSOuk2yPyi5IY68Ge+OUEKdyj
ThNmxiNRwOCTi/Or0BCWdPxR30unnfZBTavIvLyJkBjsWYxYpglcT0Hb6ofSo4CHtI+i7gsa27o4
5SZipAG+QvfEWSl6C6QRmXrmcA75n5t3fltCb0pkQiPpKLeVn50CiIGGNRMs1334cn+tmV1FaLdr
HEAZX/LTtwc7fUfu7rrrOWaIFuB5JnOQzp1CwglyB3DZMBMsoMlQ0R9/zmsTqDXxiaoYBlzzM0Cw
lDq3wcQ6HJ8sqW+gEM6rpcmAUHqAOY1Fw9Klynxd9qAfCkGnmx/Y5VRUFblPccnjVqU2JNOUG4he
3u9L4gl3PV/nfEaCw6MHtsZGDglhDHoSaU1W7r2C1uiMCdzz4Kdw0MS4PUjs9DaHfMLaSGaBsaRA
xIqtcTRYDJn9XmEmyyxKpsHUY5L0uA5H3iVcm9aymvJv4qMx7oKi1gzw1PnbLbY3b0yszqjsdF07
4liO2GXSVfZi0DUWC6uFmOMW/Pk4337MVUOo3TRrSULX/gK8ZRJvy9KoxBJTsuZF7e5rj3ABI4+G
ZwOmvZvNl6KprJd1J3SGgZ+WzIkHgJoLNhuUpA/4wlgYj9q0Xw1hVb4n4T6N3dQVSS/bOsUHoHUy
e+UsNIHcObEAG3BfK2VmYZN8KZhlYVBq6cSzG24asKeE9TVhNG1FyC+Mno6H8APCOO9MEaUwvu+o
JhQNGHXq+givy9ysIbXBf9NMN4MAn6LK5sdZaWQVdUbolXqYDBzbpwckSlahjgGHFY5riJBHHr/R
Tu1WCMb35PL0bnsYnwy9+Suf1P2qiRLU1xOOtxBecpCEuq7KKhtdIzDbWf/SK6MovEnkl3+q4oxr
h2cE0OqpqRHMgTwQlvdVS+ypNroiupPyUYA59Ou2K1n+IUrYEO5e89p1G8da2xo1//rhTZJsMvbQ
GAFEIyDyDWvha8JuJ2R5UhvQUu0cXiJYxk1kgpUIrKjCSdFSwmuSry6vFLv/4JhUqPUJM2NlhBdS
eXTsVQbnEcAYqVMalaELtGnA8un9c6E01OnxjHYfLWjg/aBOd0ciH1/WKxz110ZjdNVGudA/SbJB
MVoXBMLFl9aSQsmtos3rEA3LeeRcddzp5NcitP8yUnBpHE80XYBaI/zvnZXo2PeHW9pS4K1y987p
x3ViO70fJ54IkIgMHbeDIQYLfHis+wA2MXyUJ5td3K6W+TqRoMIDNq2NiXcVcwI5DWbP/so2wU5l
vbyStDa/r/38XWLmMqUAUIoucCxL96ISV2mjwhx7ZyBShpHJpXbxywDI+IHFlTwPdC3n0/FuypUH
r7R5f1h4SRlqwRNsIg2sL3WFsj/FDuILHVhfRup/eHdkiIxD/c6cUxlqtCD1/Ic6Q1dSj+G24hLC
SnecJr14gl8wS2XE3f573acKF87lc803R2W/oJUfMQdUWVfyvebtjXPp1kBNJOANq2F++a8grdmh
D99yy6Gtr5JhARZN9ENkS8dSXubu8F/xI6+MrGOUMMUbHEP5Q54DyDAkMHP+hNQIVMMJ+nmcqDkZ
yXtryFM8+Ue6FakVCXyCUgEAI8VSehRiJOC/Nn7BwqixgmtgBDc4jpIKB+RTvFpeDK7D7n8gzuvC
tPOZJrNt3PSk3LuzIPAMIkcGX8s84oLVOAg4whKLwnTXQy99815NAWLdtosnBUs4R8DlNarhOIsa
ZxxYaFrz38shJvDaaWAi+yIqC9UOWUBLF0/lQ9vLneieYoZiLAYkdAAKhuoaUkhVbJeY0KxDUzFE
taxeyBjrPaesr+fzO7Hb6a1uMbt/Gqyv/8rrYBRYnsXvg2n53yd6J7+TDlO8VtpFrI0VrmDrZh+c
eoFCDTuTu/Zd60RlSQLWWLV1Gd4IJ4QOSTSCOHgJtuvLSzvibi9+EnfXu9qauYZnF0EO6OcIoJ4j
ldi/W4SYpzRzR/oPURwl+i+iZEuSRPmWsbG8LOgSyakpUKxAaCH/SYzKsv1M9nP8hNzxASTSt2wY
iLCwxp/1axDQyCR2K5FY2nTtEQuBP9S8SbBWY4wK7SrwNReq+rHQUm2W1ktCQ+xeAcqZG+4B2xYM
1wCgLYl16WWBJEWc18AXiIa3pPet80mI/4U0oRjUF/wPMIb5gWYiOR8F+R3JL/gwKrtJj1zqEQCz
2j+2RiQ5NN9ri4SvpZpoa0SNxyUjzLHqESWLBenDSmQH8RLmHtxIvneNjPYyFtGXEYYQaoLsZ1e9
eufZraS6i7tjkp/BmIUW11byLkMWIGgLhdYZ71H2JA8htt4TasRHvykD661mAWlXBYPN364NSTgO
olAQQYaORXVz8mGL03YAKmVtrLCLus7+UhpJClOaSIU8r0mBXvjS7F2KmfTw4EvYcv4WKdUhALbJ
sE0u+6x9RuVyikiv500qX2mrJwi4UJmRVxPZFZMl8UB3/ik67wG4eOvZY0dsgbJ2LyJCmedbsfsK
dywF0ZXhl1z6cIECTX5Xp9I+gwhu8yC4/GfJkyKuU1gmwkkb4fcjl6rWBW5H47+9Wi86Gu2ikrsj
0oqG/7owIhyhP9WBx5oCKyUkkiiciVNXBTmQNs8xoSZ+Z7ijbnPTA5XfX1YB9thxHZHn3QuWlv0x
AQI0Yf3ARGAr1NOEXlrIdkJZJkMfMnB0b7qLTDJSbTBImwSk5pWQCtfigvnPcpIldZcQvdN1i1XZ
wACXQlw+IfQclZgQgIzemc44VaNv0pJfVbzpcs7Bdh0ElVEA5PHxkJ4zMMa8DlzH9+3dZMXQFk6p
Is3f5GYaIawFPFD9HfsK4kpxbMAcbyNzu+u8kckUg2Vy4eFWiOqiBE7B79MGjeEuZtaAflu3krjV
sCARSgKSVRnKN8UyKtlo61Dnhb2K8Kj1cbJ18QFwUKCNL3EsHUev0EfMMv+Rge3rcJr6gLUWcRW3
Oks7hIVzCO6gnfIwzjkr7T/8jRiwjIpgmSsshBt3v2Nebp9znbh1/7k8IJdcZNo9oGB9ETVZXTOO
DpClwnZEbzPEDhyl2qPOfZ93Ta0Q4d692POlNf7D50v2DHDkhCebm3btJ+3MwS9cP4GraJ0EZmpa
gOmSuLMcZPOPhpMFYVPGZxb95PLltZWIf6IYN5Bok/RDjfzpxHu72cxsqkq79SwrKxEhtdgE9eJi
g9MozZ2C9Jkz9IhpGvDggX1PwWJDmMfhAwEC11+8ZOFC/7H6wiOayi17GBHO5yW2Z3kiZRrZ7p/V
Ng9Dqq8e5ooAW0VTaQcmOTD2BGiocpjozbx5rP4J7g8DjckqBsSlVqz3+t3cftyOoLaH/G4LDJov
opEqhZfU/bO/SUi3X3QXmKTGuNGGz0LE9dmblGOusjK6tLK5RQ/ziVJK8qkjVNtodgo/4yeoW/ym
d5ymzlLtB/4lnetPQFy3DfTmo7oPHJopkiePTcW5R8NqQOwnFi79tNVigtpRSHpwAI7QF1SwKwpd
onV+Eh4sLA24WeWlweOK5z6d4QzlA4LCgQyGqgYsEBcPpuYFMky+Zt/sSTYYSFsYA+PNDwghYtih
jINpvSrQ0JwcawuvjWqLvrJUQjq8Gl+DjEcj+7DNwyHjPbeCEF057L0X3nnCoeYkOjs523cUtNVg
xoE3gTLQ+ilYbSJy9xWAdqgQbMD3M6Ls/A9X6+CQU6hFf3YuITwT7ZNbC3+TbTRfFrDIK5eCeNhj
96orvQD/nJaYkRG6X5crVxejIXr4qBtqfK0S/ZXBgAEctb/mrCOO3gEVIFKVS4kglgC5b6pbUi2m
nZVtPrjoPxHeU0v2GcyZ3H61U3iqqXGMOc6o/0vVVYMNqHMBtGF0feV2BNq5j0yVpmxOdNfgnyfS
n6gtx9RKr9KcnGFDL+/48vC1JQoIvBra4Br7mTuvHVEdMHYl4qWHXVnrQIWaIREp3jEFew4YCH4R
probF96LqIdtDTt2GfQaR5uBzajKfLb1+t3R28GiIQOxXSs64NhJcbrFKugg0lSyk8af/SiCvslq
T0Acs/AGK/Nj9dnNXYrLJH0MA7w+w26DxPtMs3vHtP4XSnldd6t43PzRZXzJO5lhVOq3mp1fJ0Js
CzucgotvW5+jkpnGOJjM03ms03kdlDrCMeP78GGikKMwvXd3kZ2bXK0EehfmMWKLpvmEWVwF7Jzs
cISblui0h1EpWB5iqLF2heU5QV3YzGVThO6zNGWbrUnWzW5T2Rn7arxvHEJkQxNltCjqVHBkObsi
tuc17EUzxp5RpUlCHXTP8G8HgRioj42vr2rZaHXrCtCM4p+hpdKIW15eR+MAONdXml0wanBXMgwo
sSlt+ibQfJ9RDqMVl/9r07z3kRetYnRy8Hq1VfxUtUwTsPfGNC5PTr3AHZCF7bgovwKP40IKSkwo
OL+E51onLZYByWjoPkE/lwt9g+FM6y9lQzJId56jo+/C9qJQc4VVrAQYa9aNnWi0CLpxoAIwEWTU
ByLVmODXB1In6Q0PBoM7C6F5VtxBjvC9l0njJvYHvL4FSuoot7unbGK5axtmxylPfriidw2CUUGP
Di1y/wtpdrmeLw6Bb+7QfDQ1rH6cRwv8oO9oRryKCBUseWMy8AUl9z+sPQJUMUb7zxwk6ZhhLrCz
xr2rbXfDANcXOMKaktMVZPZHwrEkVQ3aPtejc54qBkwE6cGSAdngFy9sW6zyMjW5yyuMs00VhUsx
lngkrYUNWQE9uqyX/5Q2lK/KOkgC3h/3qbJlR60RWBNNR6eQsVg9l82cMYahJzWgi7OKKQtyNIhF
Smj7LydcTwQ/lnauEZFI2sqAmj5SDb5yAP86Ocwdl1B2yrz5zagJ4GzCHofh/uC9JnzkeS5Td+iV
2zJXTDJKupQiVvhVeY7FE9Ze+wRLL4K02ZK4OUM/LEXcXUUZvVYYpDbcU5jh0hfo84R6JutuezYu
yFuwx8BKxU0/8zNu64EFKfJ8pRBB2jwZ4OuT39k4OF7jdyZg2uu222P12kz4jG2YUbBEu7ezd1UP
dm5f/0HvOxUYVMKoKzJuB+OAxYR83n7ifzF5kJdTdRwytjQ3CdOQgzUDrZqP07vLRCQjA1e82xZF
rEqkZRgCZI3Y+8zVzOf+uOyS8ungCuD6ZKolc2JUylj/W9g2xOC4xtiONXwrPZPJSaXBDewrUKW5
4YcHSic/Tb8/Wv7n/efFUaMCJ3kvfQG7h3ae2wt8wVbZ9P/fAZ94UJd3mA1eDJ7731OZIa3d/ra0
uezuDpDmfCKtkZkAx21u5Rz5ye1kUNCJxRLqkO6wr+QK2Egkeb0LFFsUk6JAbn2gmxy0pDgW/4Li
DBZaerCLfUyLWuzEzt/KAkZI5gSkLplPqRDvmTD9lkHbswWYlXMvn/4f0nn5gUUoOT5a+bmpLSl0
6KiSHt/NpY5HAh5QW5wZ7a5vDOguwi9b8rZGZRjVIOpUNH+u2ivtOerIVig7/GafaS65HylMyGzX
elC7eStPN4f8eFjZ2n7Wf9/XU01X1QRiSuVg+q76x7cRnaJYa5cdKZIue/atsraXHaHg6RDwLNyG
PJhdVuxBDmPPC8cDOqkZfKwQekZjiwTMLwwleK+maoTq6r/47biMVrPwe36HFJ8XmAq0eCnGvs+A
0MUUKO48sB1tNWG8572tW02yn7dfUgqgKvERG8B2n1B3FiR1Fw2fJAulqnLjTwX1TKmDNYrTa2YT
Wcw6eFNgrif0CSSNxfb09xd+ebuLv9o+iNe2uGU2rm7GVtgLjFPzHfxGuaPpT7aPaFahpXthX5ZH
Hn0tm/5MQNeJMX51Hq/bVBeDyMywTiZxBLu+DM8JBmClvvYaBwVIXaUoAMQN/9/rsgIx3EwPriIi
S2U5Enpqj4FdNfK50QFseV2ax4U+CtHofx8ynsRBOCDcO4pwAOMRDVLUr8AZtG66UMvcNk/oA2p1
BMT+likzvd3+KezP7rqAL6BxEdSvFbCj5TQtgnrSP+1R5bmSZhmvAadYpUdqm4BqqCZ0wCs5mVeR
g7tY0MdOkEsFWdclY4ST+o8T6Yvw84mGESrvl8C/XgkVjUh8r+jvPyUoxoLe/xEEm5zhGj8WktQd
XLcbez5f1WVqYfNQ10NSb+DTVmAFg0SqcFM2c3MLMThwbqzlSpHtAqbXCNyGPyFaJlwKu7vPUIft
QF7u9eaD2kiy6Ou51575bAJgsXmsTRz7SLNloCNFHetqvxRS/Z5uYXpmUYjIpa1Scpn6h9ihLN6d
cgSNcLMrtKoPbTDKnsL3qQbB9+epf6mi6Bel+SOP+kTs7DHpF1MR6/jq0ZDUaimc9EW37vhek4U4
pKI7hgahA0ZIR7Go+3rfuOybJX7ZcDEi9iUFLuImWsxuoc2OzNqx4XJFZSsah6ISx/mOO1o3/k31
EkCsR9RzRFA/YpJaqa2ZjhHPb/rjZ5T9jy6R0fsPfLHYVhOZnD0epXKgqu/0i4xr7bP13K5yq1A8
vQ5j4gfgqIU4OE5x5eKXe5Lk/oyK2uQ5M1uTO94LrtXeruiH25e1MfKMVtr1pLKMAVbrxpg1GKmh
4UiR+e1rO8sHBt6QfoJKuyDLjmahQSTyLB5y/vXQ9ghET5zVdrD25ppP5qCjs84H+ndGmeBgPxXl
x+EMj/6BJJzyfgC1WFq7lKpa1Be7ZVwG7vJ3A7ggnApja8cr7oWm9SNFs7fL33TW7wxhRcbZB5+E
/BpjuSSMVMyA192PqGFcvB9j5g9nBlc7OXUrJugQEL33biME7zL0G+W1WtB0rWiJK7cMzG/A8R73
slKYhLkaIbMwHwDjKF0/nUKe/CiSEwVwEYuNLgJThdLPDbWyX44qOPxRcRPM6IMmG6BJEMN+ODz+
hR1k1rpHntb7rq3abbCcjm5Jz39oLVMuu4zRa/E2XP6aFn6bSgXAeju6N4PklMTcsujSRw65CAz4
VCK1IcHp4uWZTU6Zj8BgAMzklBzoXvH5doiNRQog+yZTD06BsvPu5+v+reoTwPZRU4OKa6F9qVVb
3efoxNgfUrJxAwr2V38UTFkZYFxEttX3l6yCpi5QNhudGYpBIhWbJr9DbGuTUJnYAKi2+Ymhjjsm
31x2W1EISbvzqkKHJnz/F6kjEyFSlHruhCpPoj63758LmITKaxS1mDnX3M4N3I+8jv7UnRZquFRs
b3VzxcubiTo1DP8iIP2Hz/YotpsfuIi8DLihB17NnYA/T6TFfINWsD7RW/oKBelCIE25a6YkibTV
pX0qPBYz9ePm/+zdI2OzTRozAFFpnvSCA+IFagVMFttjrJKjjYgqXR1K6H+lMBlMgUzAXWIskWpl
7glj0eWdeT3LTj5cXF3jV/DQioa6UB+JSOK+Go6UlY1QI3u5eyJOAr2BFaRsymq7ACV7D02apOJk
Kt9eYAKOh+c6aNkfCXWbKURYdLJ/7FHih9+3R5vr1BzyL6ZDqO4Em7Wcyoxdhtk/1GrwngBqW2tw
cOt7Wnia6NgrYr3YHdEqa80iBHIxl2+6DwK+IXOvv+LeIAFjJ75wObm+xL/hOQxY3/lNDs8kFSNm
7ny/FDqhqvy3fYDWxH8sQz3DruaO8/NspfDJ0DFqAq5D7dso6Npem34KMGIB990P7Ebh7Ahe+T+E
W6JFuM9rwAlqGNyZNiqejBUjCoHFMf5yNWIMNvPqYQt6LVFJu1IJ6Aof8XVz2kMHXzSAGlxabucM
jNr31BlBd/oIzzu6BqIwhA2m4ntPUO9zrnhd3EJL5jrkLKYzUqWScF21MJI1AJWx7oBv5U/Z4rBm
tHE/EfjqFISGHJ+4DKGIFCp7vhLUZui601y0m+Fb0MPtcqW52dUGp9Mn5MdCegouuMnlIVvMVwgu
18yVZFQaibf+EwuSsquZrUdMHZpulch9eC+c22W0d6PFyxkIAF1iscLicfWUDYDE2FOWsS7jv2zL
F+5ezFKzgJ7DpMs03JPf5kIr0Fa7bmGKhc+fgnrOZvZoJFPKdzaDt7f7rD3IhuGleITXe8Wh7Scy
p8UThxl/G+TTQYA5cY6iQ9wRmpc+fmiMJi+4gQiRqfx2LJAhZMUjpsg7mKc8GTpK0aDYy3j5x11N
JAPQGE9cSGCAoV7VGHq3+findjoMEa0EmjItkhK61i6rbmK/5UuNm9N0ez2JMQ29fh9TKHmewEA/
NucZLMgDpXQJG5oX6nOtiURSlBSH/muZH1yrjdBVPxhlreVP+YYnuECY1akg6TqrjAiy/AdCPxfO
PRoCMKj1uLBW19P19rrgZNIrFAWGaQ+nLZVAg4DArft1RYet5pnhIp9Yj2MfZAVFpC8/aY7ZgbJC
tJWsT8cdqGKcFkV0Ewnork66WLnk7I8KuGVLIXbnINzfCBQpJHj+bO7+VVF5R8qee7YnvLUDjBnb
gKdK3ThQAokst/7AoNG1maXlr2FAxZz2l7a1K1pyrzq1NLVQYsTX/g2Kid8GSWNekgCMU3bPU7u5
nrHlTUgaj29ctlVr3SMOnlmlaD0MeGnKmpvr9OG3rlkz0blEXsKQFOX+hMxreKSNXUlzFoxCKxJ1
kjlo2/C0Zc1HBYIQdA/8vdgcDGvg6lAwjRQeApO5TgohgQq0MLLDyy/dLSJ0G86QrkqTNsXyzNnL
BM5HvpCaxSM/+ZbIbh/ENblf40Abr04gZ/9uRqSLrRHUAvcB8ZrlY5XNNaFCkGVQ27Rwi2wiXLuM
H4sub/BurMxGSGWnLa2AAEjn2C1FeKGdlPPNy9TL2Du50yusLRk2by59sTLi5O+hRg1rdvuO++ZO
bRlTprZK34ZTVG80R8bVDIip7WFxpRxPQyc5jEAAGvOWLxt9P/na3Atdh3PWC1E0cOklFUA1dA0L
n1AuamAA6L2UJPjkFvV5rAucCRc0XCsSQh28jvCSwiBteVhbm/cWxV0wn+oxbH/Y++iMUp4WSKHE
94SkoqgH960Nl49eEl5ymWBK1447WANmnOi5lY1Yvjftu+MrKpbRZIfLhboNOOEbJQQEO0MY7LDv
ky68kx2oTuqgSm+LnAnvWZoGBVJYaHx9uNnJ8pQgmSsrtxGDMbYagbFaooCrFmX73w+fD8gQMXZT
B3DOGL+s2v0SMeQg0zcUROn4thniyq9hbw6AkgjIF8VcFML5Yei4V+vpBHhW2gWNPbsiaRAc8PY8
6Jyux+jKXlg+OcTsCraBMqnURYQTFEQnZ/ZIz053rVsTVYmuRljWY7sE1TqBTCSwCqegOUO89oaP
NXviZ/jeY05MyoIOy/qfTX41+vvXs9t5lXTVY7RvEC9m1CgKTCrs5BbxMYQ1/3NCzt7Q9T9S0Rym
EDEfitjC4P3wpx0pYYHHFSugKY32qSNRovJ2VU5QCrqqu3OGrTtBou1sJ0UzNrUeefZ6fosIFY2O
jLvF4bc4uX90keifEKLM0dmNxKvvJODuXW/Ygr40J4KmFuGinE2RYwKaQIIJBO6zgirbxWwL4Cw3
XhDJzxlBFliqntBfuX9ehBkJJOn3Mmb4JFkTkW3I0m6+UIYKlsMOTnpg+bB2R/GfCU/+8xPd3Ts8
DHTfJMWpyaxzB43l1ZXUnOIIAf1fGaRWEFlU3aPzr079ANbySTAWVOQsmG/A9ezGXBSV5EHwMk3z
q1D+lwRus8kWB4UtY/8aC5nJ8UhPh6lF6BAo6S0YCeM1ELb1TiqJh/mF/DO9jmG9Nz3FKk+S9zdg
2258niWu1jEJGY1mW+4KCDPdILzDdp92Ye5QTLTkONtr45RkbMbOkKIyrP4BrBMS9/ZKOw4QrMnx
knXWByQ1XTm0VycrefkIRF4wJCpEV/Sbw40fKMgvyDSjBaBo0KOeYo9qZ1BCVDMyq1hcGrTKbnKC
11Vz7FNJzS5uyqNglIjQFeAdq/uFL7lo7ZmGHqzkf7t7G9MTwPv9qE0k9hF78wHAnmrzhP5b/WIS
6e+IBrvVi+FJwQC78IwA9Ixz2XXq+geQoBgJ9t1P0ow6NOQORKCEr7PLXarVknMsBpdtUQceTCLA
1SStmml1NR1BleRCmbkxAxX2tQI4ZXTB0vuhRWEl+rgldGZ4sOfpWGKmW5pnzGxtTri4vTFAXJ6x
jD6C1MmP7z2syjxhgt8u5A+Cdx66mT64FVFI5hxdOxar25STuWqI3/9HcE9PQKztpQnyrxCSUIvr
4nMDSqppejGpH6iT3aGYeQxlyNvMDAALtviin56fS4hZfGh/fx4pKcaNNZO/ThbE09sYuckM7ldO
HLCV/wYkN6GIU5AIZBRUWTzLHzqjZCN9t1/DzLKbAVj1vY92mHRx8LwNahXZGxUmkyWqATBXawPk
fQ+dvRW0d2N9ZkqBOQHP4acroM9WfRSNW3gUSVnJ/iaxIRUQupc2Ok0NZW4gdoktZfkHNbjEr+D+
wHVAVNoCkAe+NQeaO0tYtPMd9DlljqjKtmaN0AYSza/DHSnq1zyAMxYOti/Zpkf2EZJjlgow16uu
4aElQzF19OTZ9djSp6/bL6WKbOqj0mfRWNpWzJZQq0Gg+gj2k/pJS5ig3CwpOYGG6ZYUajFJ2sZQ
w4KLzwizX+262V5HjehaEO7OeftxJi92Hh0yRiht0PkaaAh3QaqX67DiDhnknuar2VKdUYzFkBgj
cqZE44e1fF67x7jkkabdbV71v4viO8AaxCLHg82FWke3b6z94bCm8AYb/mvWKCCSEaXbXJmGwg2Q
ToRJNfpulTR6dzos48LkKleeXhP2aKcgTTacyYvGVFfez2Baf40pPAUXT/wBpZGunE4J6GmDAqiI
8rwXvekPdpUQSdjuIxbWjbSfw3zBvzuxhU5NW8v1hBmamP3YMpE7qz62jj7NBn3oqIrh/mGr4nOf
mQO24ZQ5pZQF/VobORWd5GRXaQg/PMMTg0KT01Iuirsh61b0a7JNPJ/QYidC7AzEXTEC+xkdXuJQ
ry2l5tAoTUILhbfKs2ZE3CEjruO/0zbE0WwEqSHrlfMREguqNjd4YyRkpamCYAoAwrG66I4NLBH+
fgmWHmPQMZAall/fw+L3cO7fDDmqRoefxHHNMwGnDGNjlba3eIK9Y0wVvhxTLsOUob6S1/6GujcE
ZaY63eFPhUHabFPtTUNFztIbLQ0wtBhBcLyYw+tAfRL6tcXyH1AGGsX01mVhDb42pJZ1Em2yI4bk
30AoL17IWONKARZzNDpN3dBzil4YkDWt1IalreaNQwhk9kyiatnVEKnogGGNzqy87duHRDeYk0XQ
B4Qb4rjWJihOcO9Jx9xfHMRQ+J19WHabWse+m9TTFW62U7GJFkmB+UpWJR7zstbl8LAhcfYM7mXn
KtcZv+djkEHAjlahgw4i1TG5NJeqzTLqNcmpP4wOoK/jdt0IjlX1h5uUMtJtBIqebshtRT3LNXyg
F3zVBLnOaqfeA3b/nvf+1F41l15EXCkX5vC3XHuB5tiTB0SKWHZQRW4I2mSDKNMWqwE9jGNoUmFi
+F6MjnkjxL+MVsfWkJx5V2A7rCObrkJLMpm+SxdsVk/e8Bd6eNCtNPX0eTc5dWFSkeWrEul/fUdj
U+GTARiKRuwoYoSThtmRmSg6xLJ+Rs2FKi1jo1yTWSWJJ7PRUnjvPBb/2zRxKY10jj5ecOi3DlM4
Oez83p2lRrohpCLktooDETBbN9iOaf194oq8Yb7fqKglmURUCQylbejlDpl8sDdCaUv9x79CnYrX
HQJAOq1BL2/ukTFs7R0ITjBmxjNaIxUz35RcOghFISAVq470dag70MOkt5ZHx//4MP1ImLT/3MJx
7D2RdGT1cqaq5CKu0HgbIx6HUD/XIY1sqY4eR1Xbo+MnGPAaSm4dvXp+5hG8Y7G5H/Xmye22IgH3
eHvBBOjaIYyY8ZIrhGKQ5YhGsk4a9KZGJJ6KpuJjQv0CGf9Awz8G6d1TnfwTPeR77rkZ6AAufHHo
q2lRJAckzgNS4MIF+EP6ndi3BuT0lqRbFeeDnnPCVZPJZKB4M5o2ijScPXaLggZTr4x60KMTVxpS
VBs06BaX/kDHjgg7jlySXL+lce0/NHsNIg1OBnNbySPGGYVnfD2rdaKUJQ6DRVkL2l3LV79SOF03
RXhQ88hfqX0JNJMq55KGTTfzH5zsf1kJ8DCFB0bPc25kQM9vOR6WazFUIS1JStiBwEQa6Bmwf6vI
fms+1gul2Eo4EnxCKCUjPOsXgabD72yhSihiPGnCoP6yQmPXfVxvMzXJt6Snz6GVaaiaY+aak7tg
J7UJWsTBTYesJWFplajChlsLgSWNDejYLmhJa0AH5gV4Dkl7kFvZp14KtWcj2K1JRb2GBGIgUaGB
xYur8OkY7rg8ISQc6ka6msWEF/7hbce5TG+sD+7LXKpW8eRv7Ap9TuqBkH6hdZJ/jjEuwGbaRObB
5GDlEK8AECaUFTkpTlKXgC7jLp6j1KRBHRmjbxRpgAbIkwAswyZAYRajS7rCv7qmOn8sox6dp5gE
TWpmyshunhuJljfK8h02HIy9qXfGdpeOfcZPIvKoIHhyRPLHeua+jaFmrRg0Ra0irboshPRj5mh9
7lVlymGlfrY5fZoIhxz0uKZB9zKJSG9O0+580KurXN94CUErf1Qx8qlo90Whwge4Qbk9Grp6UwL7
q4OpVnlVXaT5KF/oCJTrV2A4O3uoB2YMpAAaLG60XQIJcBhJNhdsq2isyJAndJ9YrgE8v1kyQUA9
Z97d8bpF/4UXMqRhVc3wvA8IqP3XmwT+X27fUhdrFiuKYS+8ygAa5TBxBtARekkPyF/XkFKVUlbi
Awiz9jQ1gpLPkHMuJHDUQIBPNrqonM1EHH9AH4KiB/OF+U8YXgA2QU6nUyKxEh2lAKAp87DUq7l8
vlR2Qcg0U8o38H7EuPFvQF56jYC77/97+b+APNfDT6cc3kXUXeOdo7xGz9JLngLQ4lHUEZsZfj3B
sE2i4o4tIiFO/7wyfLYrl3VNp46StRuYLulIcRhhxFNH3pGD7FNDfzd3Uo46HNiRIvBY2RpwfcnW
HX4CjdzUl1ifXyZ2g/SESARYrZOJZMXtBBPFbgR9j9MbxQYthCkmoRzKwzp3wcHCtweloq39N2rP
CUiUJRgktJsZ0MPW/MzvV2p9duvNQn1CpCUA1iJQtrTvdtR3adn8fFXkV7hZUaLI/Paw4Rpx51Ss
ZMqvJM9YAz/5MjlIhclPbWcseo3zIo6x+cLzSn98tf9hKv+X3VNRe65mraFc05ysxeAkIS5nAGoi
xdQyxtpU8gwSaXkJfGRvmZ9iEXN/8Cz0hQLqvFmaSHFCAcdhSXx35CTnGNk+U3KiQdqec5JpB9x8
icFKGnCebf6Mpu0GKwDmAriEmtAygs+k87lwoAj9Q2UoJxTs5WUE1r1ic9YC2nzlznJgGNARSqWb
jbsVnnofFtuX8uY+B6U3f4uWiKqrVGrXyZkp3gI3hJQxE2dbvM9/dU+9vUFC+thXeA2vOBhNGHIR
BLqj2662lbEPDxSWvQFW9UuGj0xCSWX1az9YM4shSOWSInSqv+o19lzZXig4UX2SJYTRodzkH4NA
3BdxKaIJLhrjzpNoK6pURkZtLQhIpMm7CEspnZkCYRAxIkFruMPEjAhjFHLY99KVXb48ymSrsFcN
28EAf9aZRxF1APaS27nN2FOhn5eva9IJgfpT2b+Pt7A9qjY3cBQHW/BdaZrYMiTMwKRDWrNtrXbS
yLIIX6MoFPV0JM5tU/hqdss+28YtIO+4GnTok07w7XxRmxE1i7heyMbe96O7SHp5+2tyFpBPBf8A
ksirnTPze0EUOWcKFlrY4N4seNhdxd7iKuakSSmLtWT5zVyXAV4YqUA/6tShAidRSyOjLwRIh6XH
rG4y8p7/DYEYXJlbhuxucLtRLvjY6+snADYfyqHieNjYit5+tT+YtyyP0ByTJ9LWjXbGBHON7iBX
HW7CUUkgmyFPEVCOretQ8OuCyd1ll1UwnLjMVCXSiC21zEn0VyM93OZ2fzEdRFOLpva/Dv+daik+
TZQjaYRB/HcwUYYxCvjeoZIwpHyp8fLkAp52dBTrXszGTid0mQm3yHPB1F7n5WosUL570LZjtEOm
UIjUObZfXxqGJ0G8Ubj7W1kwH+HfSr/FI/zIMFoEoSLPaSc63k8Yg4ElB7QrOQzo0ZtP4iNFfedV
WKsfK0cizrf9ATvYG08ZJj3bi14Zo35wmOcddLKFvgLmo/89jbxq3CfiUHYZkpGmn2MjiIm+pW3K
7h+jWuhE0Mbzn65OovNp4AQwyPWe4krxDuSbVdeTs6B3KYcQN6cadt1vGXaBNqBVbxNUibq9bJjF
i2IzLgWn4zhnVd1rTx53JlhMRbIiw0AvciXfA7UrPnI5+q1Il0lvnbv7T/9V++By72xI/JCOi7b8
MwPH1V+ivy15pXxH28sDuR0sr7ot0jYkdTCdSMcSZSw3AYef//+SLDpotBzvYPO/TgNIY2+E2h09
DxY5fu+0OmORUTWUgRxKk2atKPR92j8EBQxi9lRfQXjVIJRtqCnUnkpxmck0DMStN55rJfebXONj
qtrd68UuhzXLKo9NKZuHPPfy7NV5k7xrblTidDRStRyEizl33CJXX44Ltriq2RuDl6E2CrFchoXl
vHn9lzehr65y01zTlbj2X9IKJqCoB7iF3LLpeyHiBzhOLRX4QaQ1zB8bMOz9aG8sOPsVb4fd0j9E
0X2i8Tq5MACCcxO5x8bSrOxMORtY17PnUKzECF4KQo/aG3j5gyKKfY56ZmZHzXnINVySM9VZQbsu
BtAWS+99B/S/FTFfvRJcw/xIs7gLVBKsEXv5Tmdeoy3kBZjIMNStrgW9pk9Cl3kGuF92rBdwgc7H
TzAqiGJg6yURAwV4oXHoa3hzWdJ4/kE5dFSnsG0/wCTNj+YNB3vU5MxrVB0FkkPQlG9p0CzwEKF1
sxAUI1KMswGxWmL2WfQJqsgJJex4LDEupbay6JI6QsBPOMk2DmlsO7EoUklm6lCRBhoCbFBFIcmT
VbPxwtvcWPQPOwdgfWvvR5Hsa73xjLPbK09gzdBUaaUuEnlhELnIwrsk6WCJnr7IuHSXNmtbtWxs
lJej6I85+54HQNCLqD41nHMGIKDUWafNtA9yIDmDvXsO7JwEzpEm7o0CAIEWrHVQujTMJ/YTungl
BwqWN+5eqrlIHmQK6UWCA10d0+PBc4+ZyayP1mTkQV/1tSxWZGo9WH0XJT0AW6M90ZWbG7/AiPCR
IgaMGFi+cMcwT1lfPuv9XbjpL0wnmEMuYOSXnzOQQbvXp8hQ/BgISw9Y8l+8bFrarA3I5KnS/rXE
yOMduP1gAfHGKyECNivBsKn3arT7QNti3KRVILn95RxMayXwDcYfC+voHpwZW+W0UCY4q7wFCbtM
XLUHhpB/nNhKC/txImEUUNozltsdVJRmHQSAkpGZPixT4iNdlUrhkXHuRv3gVS68zqZdgKgbUdn2
RgP61pbdxA61ynAQPIVtXoqM9JD24YgcuR04uAnUYw7KkWgoFVZrcHGyxECIJask71uxrUZ8RUND
MRdnkPOjYRfcXhCvWCC2h6rBqCyhUXu9NrqFt1pHy3sDyAYzJL5ViADVD8hB4A4ruRTg90WRPL9L
kcwn9h3DaH1EmOUQencvaq4VrcLIMqE5oW0V3OL8kzxj+EHVhrmjBQqHHP/kLKzaSLQFHMWKFQop
yUP4o3GgNE4uGaHZ+S8vNpmOGGjCr693DiH/mRIl3V5D0rYo5IBQ3qKwvL657m8wip8la9WPhDEq
65ondk4gMGPeJ62223zmVYuq402oRgSWIeS+ujlJZ5qkkldg+IM2Z/FLOBOfo/VaBSzogGpt97cH
LrUGENVNPcOS0Yj74Qbxy6M9K2Ifmjq1Nm0dTi+V8NK47jnQJ2jY6tiNMdcQcVtFbCjMV9/e8/va
kPuwJ4FiidP8fIip2QTmVKUr1V7zdl632VYIBlmhXNjMiQpqd25L39LDHMJPF/VeegQXarhpvMT0
7PoZGJ2YXDIMfIuOZTO8IG/Yh3nXMuYqXsWa275vL0E+Ylt599iMmVTV9O4emjdjfW0jvsaYRT7e
jFyUO2wqIau8KNBDCFnFUWpYQlDg5MEt6Xjej6C6HerSbU2xRWTLTcLO5pOdpKv55XBmjDEpqa7g
cEQ5Dmxs9zQ98LlgrfJr2oz/lUCh8QNl++Z56dOgoottGfwYKhsli+4hnrB76IMArZlioFiWbbZI
cg+UM9Fmm+npGn0pgSFi+hE4BeAV4EO42pn7gQEiYVXxZTQYNuEJId50cdaGen8XQG+QmtkIDnID
P4xSsnFQREfEacZkM+Ya7RE6NdQujBUEJl/LEfTAxrgI1UfYCC1UjHpkVDdrSfk6mCjuaHfe9yxP
4KDzcYhqtXJM6jcPwlg0XoNhStQEWH7mxAYMYGy28bYAteQ+sQrAX1FXoF4nneFIBdWzntihWdFH
sVXtk6ujOGMHBUPoJWk+t45np0TFzVOjHKySNLwbg4Kx6SovEy9W4DGvuXar7l+aIsHrOfmAnR4a
Bm8wELjlEYBzNKkDtOIQOvDm0+Sx2R+7LU8zC98sCHO8XW2SmOR/fict4ghB0Apiv1yI/Ec6s1Zs
8cn6gPXVZtGkk7DHGXJXAqLRdUuyuhmWZkD5BFMHZ5G15RdugTkUTu7mPOp1x6kbwlwpzfoJCH0J
zQpnVrunE7EVmk0HBlcRmdBwWxzOCCzew5uwkjbEVOrYFuLz7leFbK9GUeXLWZkYyCHAc+ARUocj
zrmKeDyp7CVgiwSfQpwAc2fN99zwo4zOXlX/hh5oHtcgkn7Oc+WQSrMbbkpOodIiBJ7Viw4K0DM2
5L6dv689ksfrSDheR/6ed0fyR/hb3yWopYL4F1tLG4DHK1P/aokbWsBhVCzZQrIKUFMExcRQAUyO
aeevD+T4NzmAosdzKLYu3XYddBtmuPQMLOB/6Rew3DgfxroLye5IWISE1YUdaQxAVcZihXMe+R14
L3eGGe9r5Rd1hiElXZ7rhFLI0UpO2XvrcCzxmZAxy0E3dOJXcpcdGje4O60uiZS46bpL4iCI1e+V
MMziVjvu6uGGS9AzG9uBlPs4ihcTG9QMjNuwg1qy3xpVxyx3hD6WW57RsHU348Hh/Obt4P5vw+/8
Ljfr7osA9FwtUhzsuISToGbdoLlc/GB8xU5IVkGHvVaOTvm1T/QJpnXLURRy8hLA1KtL1yioxaDq
lJD5k6G+MXiYO1tujJrixeyiR4YADejlnigGXkEy00iDNnEJ6DoCmhgxqfVhsGLoCFB2NbqUPf9g
+THX4jqBuXZ4XXcsMXaLD8jLAqmFyCF1unHoYdVAKpRsGpG/nLQ7H1Y+39rapSd9NNR8FCXSrfyW
7iH2CbN81vEREQ3yGqpreUbY56WCDmuOqHOJurjR9KWxMfucehLOs1tWVkU5s2HH/BFDBGZH66la
rITFEkeapJMwzzI7coQa3CxqQCw+WmgRZHzDjTWHibNKIXn2IuM/5nK2w0X7GMg5TTLrE9Aa/IdO
7pVC/qsiUXQu1Xh43XRWbSuCHdbNekh7tinwDEcsRobi64Fwvx5S0+q6+peK+Y0uFG/FFXqh4Sdi
UdYVAaAODK9yC0bwfSPbkKnXUjHgPTPq1gJWrjVunAAMHAz6+bvm6lUenoQyODPFib5+SI0VbzM6
pGwbQ3ZICbcUXGkc2I/eKIbXwnqpyDDLEO7cROiJSDc6+zf1YsfSVUj5tElQzvUHlANjhrIucUOp
FlJzRhl18jKMmQKUmg0Iv0a49XgDEaoTq/jpfcZ04K51N3W5ruls9Lrb1IzeDl/ATZHH59/xFm4H
HeRGMuVMhAAAjdlTJ9A+rp6zwKfhLMyAkK8XFC0V3uDRsry7PpqRIJsNO1n24dUcP2kN+tnkH+64
/bcI2P4W1SyAJBfw0WZPxoGUUxHnfpjn+BS6cx7AiOg1/3k4MRoGghBeQtpJQGHDxeIxewdJkDqe
trTDrbKnYX4Vdo3Vw+dLwfmqWnSrsMuISi0E4h2hYhsWQiE3dqAYFa0t/mC4WrzOyAQsBmEElPUb
lWmWRjylWIH1Gv+NisNYrSW8j2W4Eu2IhOKOmSGv28aEzrRAT+Zivm0sDYSFDYlMB/pld8xBEVxr
4av/bbmfFNh9uVADTDUOqhIgd3606lCCti3GGnYEJElyZDkxYT2yBmEVqMss8PoTxNPOBlWQ3I+y
azESv+OpI5pkxNAfub7lqmPikL9+9vhIRTRsAvR0bEpQPN+l4jxaM2b3JZsK6bv/2xcdCnV9lK+H
5JpLj09sOwrZ1U1b/ZUvK2rcNgcXMekTJtngF5rTIX5iO9Cd9n6KZms9SRQgAkfrggXxRJCjURBr
0HzkrSIsRCcy4Q/JeCwbx5fLkYAw6xrVOeNj9OnsX5eD69P2iM1WdCvQP4+8RBI2NjJ4ZGKNm9lq
D9Z6yr0JgVt06672EGraLuGyjRNQn6a11SWHNDLgZidncDoIXBk+GeyGiCkzHJPs41JQ2X9otoNL
74MEw8JvdzLu/96FqXp3fNEMpHNSJF6ony0u5oD3usITFunh6ffwit/7isVYCRuJCa7tHUzWVkGe
TRskQX+qZzAC2gduBmVoe+nQSUK9FIaZKsMP5S9t9BQMBpDIFvQn6hKHFDmCNPdsyXuY7XCXoT/q
HmwDz8Ocg044rHlSc+HRyGMXSvG+HrEDXr5yya5OfOhlTx4ieWdfW7c9v/XfpqWLgImuZAXjR0P3
L8oojk2fAUyWDwxrKgE70/mgYGUMKpFnf/Q5noh4NeXKMYZNKiE5JPOSBLkmAIcFthxxT4Hlzgs6
Ie80tJ64HOZ9GeXhxOERd4bPwxIpDjEEy76e69uJP0lliNhJtAqboyI2Af2qXjHDnyVgZBhGbhwU
HVOgAXMALnddY0jWOr+6aiWR+WkSnl7Br/TFNZariMkdTtdZ3gzBj00aO0YP7r8A3nGukX7sbwHc
oa6TsjTQo9Y6XhtYX0iA+7J4lHPT5hkSHrOQbDuB6/7Qx8rnJV0V+3ai9+R7qs3Cq1BxFPYVrtAD
P5ZC2azmLqPJ4+99gGq9Rs0H7m36quqmKQgDLNsGJezo0Veuwvxtq4EUUI9hjsaLZbw4GvAXQnDE
vLDgIrwE6pOYMxf68BPv/dGJtKd7uvnyFbd61KxKJPRza+OKbkL7wLhxCGJ2/LHi7wv4I4RghlN+
tBft/23T7ivp+e3+7CvWf0hyPcKK8suzF+bljdf759yivB5ZK5eS4aJ4PZHztu2TNuPZrR2262HT
vL4xHZ0nEtSBXY8UyKSWadDoC09j8WEpdMp1rSe2+DH2RtPGObeQ7gmWZdLIo2UqEC53Pf/3HqRL
t6ArFESbCE5lmHN1qPQ2uzLEndWxaWrs6+398brKfuponcJQ/AqcDoo7o15lj0C2vlbNuQ99s9wQ
zm1E0qYmgRjGLl+KYP0pEOkB5XYw+uJtv2xg7r/T/6cTE0MNNhUUIPkL5xBIcUZyK4cO5+8sNMR4
H3OetfuV1EwXn1M6ebaRGfP2VK0/OWYLjNSOHspiZPJJdfVxwCqoBIOz6tyS0m9URNK8zVn6bNp6
qsq1aRw2plh49GCM6zzKcQJturcnpEQ0uPYPK1nDqDfbE5eYWR7IJUo3X9JMgsi3mY1HimZFFxZS
6q8y9nfhzV6gj6kjBD9Q7KIBvAt7uvfClWqPV4e1qpQg82PG8dp3736kVqfUHOlcxeTN2mnl8V3g
lI9nkcyVauLOmP+9lAI6OzTwjpigB3sIDxhxj7OT/Uk3zlhKFGYxmp7+mh65j8DnFRXBcnOOorWN
f8dJvTU3gRWtzNLZx5FBpMh2XBVvZDxgMjNu1i/ZCxpft/v/79+JooyagNH3iUihNn4CgfssFSHu
gUrNoil+efEbGSv6j5X/Q896nOdFh/G8lTIR1JK+7WfmnZlKZfGDXCowq9xBIp81m/G8lH8xH0NA
L8kxCsnMzbJT/EM/3APlQm5OuZ8FoehnNgpfc3UfgRFQZ1YOAzPgvbs65eprsVIpyrC2W06p9vYe
C9ukyUqBfsarKLGJSWeKCU90Gn7t0xo8e3Vl8gacb2oh2Pym3oGT5VbzidxxWaJvG14IRmgnaOYn
37AQLOfPjaIC6WetzBUKr1arEDhSPnYqhDIK46nM7xZzwuI4CPYeMHJFd0HI3EU9n/SIiStUt7eI
QDv4xsarLl8Ssbz2LBcEH4GXHdBKcWlFGYJJzWfGzT2/JuT3zMYgOZp0OBU+6P2cFoc9R3ql7qGR
CoEeFY2nmjEipgP+ZMrke5qMHnq2I+t54P3aE2Y3AQY1w5+tHznQETrvF7gy4NQA7ExMtQKcgOfD
t/mnaL7vh0IrOXTQ/ErZVo21FEkO12S9Rt0FR36jIwLVjdRWWeUvE7xqkPAnbqt6SWjqhAACHZyR
5OneAxDkG9C6T7Sdj+kVEtY5LSjkoyavwdNgsLhLl9gxfIe4yt1IakplpzUewG4UvMXlMbsYMBCr
0K2qB5+NaBYxVtmBxhAzvwmmNcpqFn5FdAhKUwjKwDYcO9dqlD7XaMY7n02TyMfFW+0uZ5L7dVYu
85p2oJ6tac4/4R/uyqojzLQ+gpNE8q5rgC34qbP/Kzw6+1xspcknMIriNBtN68dU5kf1GO2G/ZIO
5ZV9KZ1tjwISY1A9kIMI87LkKNPe80cn66JX9JpEeCFyQp0P24JWN/1wnmO5agd5Dz1Q7KCGaOD2
SRi68RJWfsi3gVnfX1DGkpD6/EN6pmP29olBaw/9jZpdkmcvQGyuxXvAnNDzOp/2Ox+H/GbCOswJ
msSVVXwkmufexSF+/soT7a9VmqT/NIylfTPSYxhoPPebGqYqxM3muyt5bo5XWS73g0cLa+B/K8+l
zLqLMLetCkFIrxdwi1w5AkPemAQT5JAp2tvQq5mcrK9y0P5gGFUmPYJG291GfO59C0llV7sViDjk
ZpeKVySYlfy7Q6xEAv/GBFWubEcoZaPFiG6bWya4X/fw4aCGBM0vKOjBGlAUctOpW7/kp5oVvKAi
rmAW+qmL0mYQTlM640jNV45Db400lE+pk6JhWN+4aDEaVbx/hUIFRT+UdrPkpVzmsBv2/FR+Tykz
ebOiaSj+X3CesZvukgpgiy3byGKzSfHr+6iIpMEAUxEKeixDbMPY75ttOPVG7OOg3sV1TogyxaF5
0Nim81q2iOdNAbUttkdJUhRO1X0kojCgZNI8iGwJxvNNvO5m1Yu/qkIt0FaBvSsbtuBDs5DNspXT
m8zMCTLw9BcGOcLAFg1Z0rG6qwWfm9Ac6CgprCdgDajUXvQC/dtL6jmn5+QobkPWW7bZS9FeFOx+
vb/T+epgXgQAvvtz6lMS02FHNaMGHXoVqiXCg4KtFG1B8XIy3jVkZqWkoNbYX0uX6Mhm/R0hnUcd
8HoVxW/DO2AIdRp/D2WRiYydQxTOt5Baqhdi/IsY6eGgzBjY1myAdeZEdLePCPfI087Ev+O2iX8l
t+/buGH2vRp9iHA3r7tiCc+FgLClH7F53Tn5Gw0Yf1jzEnOtYLnGLloR3UehYU+S+hc5EL0vLWCd
wCuY5XcqhK1ZwjVifhSvsCZSrfVUIaLW9RyZ31FMk7XDgLHvPAkcpAcpaFYDipr2QDFj/cc19O/+
Xnc8ICxxoXawwguajUUO/6BtotCAXyd0InKoNvth263uHFHqcQGInz5mFfI8zClzrS538ffx8rXC
GhP7U888P4Uox4nA6T+vW5vCMhAOdV1CqHqA69KN20Tn6xL2v0Mkl/TH0EzYzeGPcrovuhEbnbA7
hsJ+4UqzmkcklnWWsUcniItngnPLLFWNHMXxGubvJmwsk4Gr/1SpjTGcPxytPXdjcEJCEyaSVUuA
4s4UlOP/qc+bRtgn4m7QUdNr9pPwrKqZ6UBVUNl5Ty201eVmFNqP5CJWb6/4YXiDTJ6Vnlftc121
bGICrWOzhUmjvg/NvHFxDDnt3EFlACiTntpt1eZFwuzH4EoCahBPyMyB1h7j3p7Y2gbvL5zAvDLO
lv7jyAntGoecc4EvwflI40yzi0gPlg4yd9Tq3yNaApWB6BKeMNJQQ2tetXvy5fOYqzVpZThSDFHs
iDGkH8GtY3ZfQoaZ9CdTSGiizw4OBTItFLmxsNFjeTQJztb9pViViDwAcfsdNh1qDloidsvWplGE
1za5ii9TLpGAADtYfticnoT+uOJCzJmuW/0jmQoVLl7zoJbcQsL/z2JLqwEHVvi8MRX2iQjp3eQ7
vv8KRJB2+X4YLVwiTwknzR3GJQwcP+6VbMudhi/sfdevV8/GaFTNtdB7x3NbgYgx7HuDcIOfs3cl
lptJlfJKKV1Xb0Z+Q+NROm8jbzyaCg4zBlZ31WuIQzAEkdUk44V4UcP6NaukhW3TjZ7BIsCHF39i
IDpuBjDOm4gdrUuNy29Is6qFyY0LlvFZtBNUPrjs75EkWNC+fOLEL4omXGO/XjjThMQwwcnI2QY8
DHGD927YuTb4z9tTy3N0bS0vrR5N7MiD5bSSf6gPcHboJ8lBs9kKPNPWiaQzM8z1h4GVbaxEWmEU
x947PBiDk+Rnvz2ti9tO1ZTXobIOxglAamxxl4DHtnOc0vAZ3sKySiIuhtAkfm9xYfdejZKQmSTj
pizEI07lel/lI7zrgxS5oKe8rU2MQsKy9sdVZsI9NoMr8PAbuNnhpAAeQ5yagsAiV9nrHMgrpV6G
hav2WSgPGiXcgjaob6Uxm4vxKQteUyLoLbVaLF6nE6XQoyh01a2TurjQZNde6A8fymL/iJlq4X67
KXqR6/ayWjQFrGlxwl4TPF6Y9iVMLbLzupUtf6O6SWbUy25H2TisIp4Hx2aYu49A8L8NKECmTmZA
u/aKqC/bYSRwzPAprG1hhA41VadMJZJn9sBh2QowipcDInVb2xsab6nOKi4QHMHV358uIFC8HZJb
X2W7JV2kQEAxhb4druiGiSlCkEnL+4Towvgs16EJDeEFgZFja3hpYOSPc7XzZ2SyoO621y65OOGx
byb1wA1CVOEz0MGq5Zh8K+FEw53ycP+KX5+v7p019wN9qXBN+B1mbThHiHc1GNHz2hZsFK+68Ccx
5A418emkCsfOOAsU0+sauCYikeRoiQ/zC2M1sq4YK5nS6pXZckZv4YYgEJNiLHhCLWvOfIclTg+6
KV3R8hk5drn1rSExHSXu1TBKOygjYjeKJh0q1iHfVCEmmFF3o93EPzzSQ8ucVJ7SmeI0yu+VQhst
d0KF2TqdQSUmAgzH+qffvNY7jKHcu4scE6TsdrNeyu67VXe+Y0BbgyCfkmKpm8AOqHW8hjdLCwmz
CfjJsWLMY2sqXi9cvx+ojs6IP2ATx9BmmRDE817sXYfjBexkV1L6t+UiJ+JTWLI8r30IOuqvWFEq
DeJ6NX/m2QKjPxIFmnQOxRTmY/29TUyH/qB+37TxAdTMrqmFD5UKodqUBMU+FUYLkdSHcPMvixOk
GH1IuhWN5KxlqDGXPw4VsL+fFTCWJP+YyHZaZbO7HlI3KHIf9cLegQcUOo44TG0uy0p86nil6ILk
20jQnCKBK1ouHbBrHh9LylqFWMvmu5VeUmZqecxLiTM7FahWjm3OPHQ7ypn78VSPV9tllpPiYzMX
loZXdHgKnEsRbUowy7xlbbxjDYG571p9nX6Dc1YpAWBUaTSFR4ttivzfoZGmvBd5ZEA6PYCB7K2R
N7maNe7oskXpqc5TICrDlOblkZ8ajLkdyz3mBvkStRvHl51N/22Ib79FXZGSrfW9cHhR6XNQx4ir
QXA8iLipQYsDJyNCxBg06Sq1MKvqmugyNkfuudss9eQweCf7vBG4hmj/MhIUWV5E90NBu8cnkNrS
nGkdspwgaXP1k3leJb3ybJcZUUiKFUk86Hv0QRO01ZBiI66AJkcseSDV7BvQUEjrYDTsiDPsedvm
lMPMA+6d/RTYleAsP5RRmNm3Rc9LDHf+kib519yG1yRU33RJVovxuu9rOfeskWJ6Xj6uJvU1R79/
512yUjbQKAmlub6a7I4l6NbFJYAS5tgxSb7JdJ6lsAsvG2NOKGXvQWSbHpN+YgHrCsRoP+jZdWTi
mxXThRMHDrsC94zTmH1OspMz84ffisk8RO2X10pKZjkr8nsetyRrzZmeHFst75hbyAJqT2aD69v5
zTTmwbeGM+lPB293fyodFm7zT5VAdYfB9SD4w+dWNoOX/B2OwCq67xzMfayuivavZbhDDySDWcM0
pIxOd/j+ZnTq0rC4nuuSkq8AlqDdt7i25Yas2XdUMTDzldEWqc8dpIkkcxBTqcyaQwYtrlhJVFXt
5xCrbFI2rXyk05e94GpgKGa9ws0O++MLU46LOly8jBujQBU3G30ES6hofA3PwvjTlpaAmDA+QMjm
CM1PdMlMS+rPL+0BG7D5sIgoiy92ocBydTBjCj3+QK3WNPfqoGKPZDCbsJU2DR6TJFX0Naxwg/d+
qzSYT/+n79aKTm5Iz3Bqgc9sWHznmxbKREwyKD+TNlDy6WU839LKNpiXn7yuhKYbY/yNkIBFvqPo
JD9cJkf/qt63Ijp0RYgwimwWK8qCIygV4mZ/plzRM2fVAnYfetpI3x04TFx/EwTpLCd6tZD3xaEN
QmD15TznPN3j6KnIfTIFk4REqHFZ0wulecFS5a11fgkGm/x6B1DK9wctCIQs+h3lxqTcQHJYRVBD
54lrBjgbArzihCt9HWxa3IHu7lStOabGsEB1vAXM+RjhPnRHmUbuwt3rskeVdPbzxFqurSXnS1QX
TT69Noa8TWwBez9rxtF7zqS/xK9vL3HnloZMZeyu96rGZDMJ+xd1BMxqw4VuEdLkNtegzJQFgWC7
klb3R1WcYGT3AgH0TIG1mGXbCxrNiZNSgWPM5j4L2qKeknHr781MPfJknBMcn8CcuvfMeF51b5k1
ktXbCZdD8VEwE/DkMN7fm0EWjz70jS1e2kMJJuwSDnASq4rPgChaRs9TRJizNY2ohmoREmkJtOsK
LmTcQxDOZdPMaVWFpDNBa6m+qY6ZxUWD2XXOslqQ/BPmPq1Qx4CTaLIM6vdQuatEDP/fI8wRIGft
/rZdR4uETJdmPgUqwPGbuS5aL45d+1j1fR1ADPPFMl2YPfOE6/BlBb/vGtcq8XSHLriWhy0xA1iV
Z41J/EK6BCr5k2rMvG47aj4C9fKyKrtzxDNQyZSU7FsgF9L0HkoVd01ti5QFppP9MLOHL9bdpt8A
0ycJ5xRIBUJkXTMKTeMzwFWGGNIbeLl57l5esEbvoRovz0ZdEXFXk3RwmwlQeJvxcaLfCwVVJMz/
KIfo87Yz5MucBWwFLI3AbIg5nTTyR1xOfAYE21AMIFEF5peSOyQddROUynzag3xyvsKwatEtNfw/
LXE0nPMkiXbgt5N+lAuEkpjoPFXhW2OYa7hGFoIbo+i/1cKZh+Smb8rLQk35VJw+xHt1mGEtKMQE
XKmYoQ/VreOPA8O1w8KppgMNPSUL5AxSoYa+ZH0jLlApdNbgwKADrcK2FjKJ6LFbSMmoYNorE1wl
kgUIG9cCZ5bhW0l0Yx30QcVmQI4Tj2/zJK7Pf8a+xu7Ruau52M5y24iwYxhV1hs8ewozBje62Vjs
WOmg3JmLiQzTlBWWnqabZld6tWEc7a+oiD88a1QDoUbXhzyv45oWmJy96Sh2CthiSPI+Uy6uADGe
1B9qZ/tNZjMNdZPdfeHo+uxHM53BAd4mU1gV2hBTjVvogxT5QSAaYVTgH/0jC23a/iXOc/i05PxU
XkLdGTNYPpWH2NLVOiSa2+QxCrtI67I1cMPzbEXQHOsLwJnX0sfH0QjKvTXYjJPcfCD/8mNahZxQ
QkyJGq6gdPeTjk4HGokG84msmufe4lD08VAooR7HrdXXqkiY6WBgfRWWyFqJaLfX7714//4/+9Ah
u0S75eik7vgbESWgF7hXTdDQnmy1Ne3d/w0QCEbfr1RRu+aiGRNxR0b0MWtgdHAMYw7edrxMTxeM
crqVnQt0xWwcZ3uzTIbKlx6RjBmE7JdCbeidX83kQ/q9OBYBeqbNFnMwNbrFcizb7WIs8jXzwg4j
kSXeGvVAJoDPyibHO2Th5Y3tdQKmj8B7Nma1HSCZb0ZRVo7h2OFQpGV9b9Hw+AnOmxOZvfp/9QvZ
nObYiEZ1szkyGsBliawvYgZrMmf21w134Egq/5wIM7OfTILuVCekaME0Aw5QVs7vf9AIlG+bBRF1
59igMbBPdNom12NCOkHhggh1PEVvxu1ZYkU7cL4A+P6OxLNhB4TwfThA5TeloHnPXiFM6L2AEJDR
ZtNr3k+i69U9Th323Q0ORbi8fbn+wZoM/9RlYqVRG61gXypB4UTu+ikzaQZPrrN9JDdFcRlvFppW
m6UFE8R0Ie/cPFsNhKv+K7P5uv4di0BgwilE0ZHWPS/35hT7SCUsnUIM+l6UoGbdgEZljKvu9S6A
H5wVOYEf7PomvOEUMUihI9YwzniGNzGSh5cUAIFXKaHkXmcA71zM36zi4Yg788ObxHAstTPo7Ws9
awB5WRDNH24vIXxdaq18Dv8ul9LZU+/OrHz+njRSAufWbUBtm/94waRMw07Wt3q+F8n1UXYNKfTE
mr3aPj7Pf/cGF4FMfQsHT0Iy3WgvLh8neqDPnlCefNab6+uDM1y4qmMHrkut2CKkpxs34WoLfyv4
KbH/BucV6WSlqiMBCSSbJB2znSgC//A6wDOUWFD+oo/IJ27L5Qu+LlJ0MRcRjx8/Ql599ZigVY4v
EjUq339OWaleFXcpeRFwVyC5YErPzkalSqRTQCMlOdMIY6tIgEA1jtdrFvoiMaboJAHjuSZrFqxf
J5Nb5YcbRiV7Qu42eCetab+pclicBjgDnQ6htgclI7XLuf1lKr/UuqIbwhcOl/5mfVibKYPUIhiq
d3doH7FWdIimI68vUQmTlkqfDVqKJcU2hczkKKe+jwBjifgGiOoOOpfi20uVk6KXMIei4A5SDCnG
Ip9V0tfCxMBx+KcBCZghhjHPG27rhXxnmsqfi0dzEGDqPtEcrauvWPTNnti5AMs8fh4EcUK0HMhE
hOQQvhY8q8Dafm6rKjYKRkaI63MwfhK+Re2I9vEqre+kGXWj/2ikfwBskgtIKSyp3xCn3zQFj4br
fi8Arr83ZkIcaYW8ZbFpeg8pePm4elynfsaY0PgEdTDO30hr0+ubPTDP2fPmWTPgGFKdd6QywoMZ
yjD610Gts85sL0hIZAHLL6T9qd/PGcH7Fdpsk+62N6SYdhP8USWMHPgROTHbEdNCBfgyOUQ9QOI8
NPKoeMH0Aav/vWUGYps5pdDjDOHn/Zs5YuwgczX98iU1SjvVj02EubuQxCgI0Z1sebIjpng60CG9
20Lg0AxJz3xmwtzmtNs1PchaaIhVukhSea1UN3IH+cmEPkp/cSgMpVBiqeL8BvZGgvbcXH3gt+hC
PnXSAjB2odYFFdWyEUBqWT6UJFdqpUIp6dXRR+TGPjaI6oeJ88u5SeApldBXStzty5mT8jsFF3vv
9uzCI0Sfl6qN1Yih2GpnFWfoNyQdu/2KpIQaYh7/2HwT1FMvKrMgqeEczS+I6UgsLEcAUs/qPSkj
h7a1CEPSSxQAbMTqqtHJp7Xm1oP1r1+EyWhX+VdlcvXsEVQyLSajN2cxcxpjgPpEHiTvWm39udr+
WBW2lAFdmmus45jehkd+SNB5IXQFcn+SccBNmNeHF0fgCj+u8v/KxGXQGQnidr64m0H7KbPeYDEo
JT07/uduvp8iBUTsHiE913Ih5qs7rZIoQC//cd71FipCoe7++3w455HOUKZK6Wog3v+NJk5eXOAn
wGgVd6Guc2teKz/F2Mk18K2K/1zCHv8sCipErxutRGIytYAgkgH8iKkIDgVCa9T76II+NuzWcesL
VtB9b/HgOF2bH/bN5MBQZ8377eKpEanxC127B+99QMTVAPeSZKZxjGrh2/dHnM+cvj9cVrhzTYcj
v/9h1RCmGw9bxCs3RbY5fnAA7vBRFNJfE9H1DEBjt/eTOb4nGG93aM1IC8PcPwBRDsrAUgexBYqj
WUTlznU180mvvlR1Rz7VzEYY52u/jXRVcQtuNJSZka+V6tNjCEZbODzY2Ns7x04vfsyfe5j6HOJp
+HdBcYf9eWrAD4MKZoWzuRXrGwmGBDay/lW88NWkQrYcxo0rVraxeuc4jk0IT2GyIh//j3UMnchK
C9PUK/jPNuC5A/CyYq+zMd3/TIoIBv7lqJa0BxvqSJPJrCzojafXKym3B9aLyntxyWPYyHESgZRB
WCYKk/BAIj4MssXsHInzI3e9NErUI2TjVgKRhMnQU1GtPQbqt4hkbgEFYPJSCsYn6tPjEinVR/gm
udZkgsb0Z2bmrVOHHnTDIGpOjA9e/PdD/jEIgIttRKyT7Q5g4vic3yvYt/NcTCxC+rrkPdyEXA13
0L2WmVCQhRIUr6YBQtv8XmwDqAQrSZ+1HtnujM2kNqDbZZ5HJo21hKMG5WYqXFD1IEtoLMCl4rfU
hCwslppZRSGb4tWUwMcgwknR+T9FX63wH4W9+ZqEroZnxxuZvf7fjTnSYfzh5HBhWUgp5fUejUNJ
MgU4jZJwqLEcTUUlZtygA6MnZdkgyGb+nEFcGedpSwL8CpI3Tg9LqFOk/y/5IiMZirpOOcT2Hxg/
77OlnCHntwElH9O6J/KalN2uG4StsbAcymGFopKyZiZ/Pefz0jUmVBgqTZpFA0NXU4tqoVXfzw3M
5X7CxiVoMK+tT7KFNrI+O5fRSeFGN6bfkvcImrCaseCsH5THYUXYiT3MPvqT9RVCNkpqywN7n8xu
g6/vD04rpKYE13uXPzYYht9SjFVWlCKkluiv1VLj6+k2YXiP24EUEmL8xMv/9B0NrpJ7yL8JdT7u
C2Jvg5dBuQPr1iFZtcyEymRlCaBmblJahgG9jRK0KFMarBs+F6hXkG2GBfPIYVRoMKQ4RZ517mfh
fmr8brFF5XdkpeQf8MSAsIaRHwpQs2Z+3kk4UV+VDLu9068ehBVX9ra6/sdDpO2Ifqhfu9VSth30
r1pU5KXBXCUsJulWFkuPQf5UB8HIl63AYalI6kkwT7n0zsK+E1f43/HeIjDe+EFq6tmgIh8SnYaV
G66Utad1igzJy3h6+Wok5GGUf+jMDACKfrsoOJJ+Ckgimgi2DoxIVahaUbO+KBZ0fIIjMDRgCOUA
BsDsMKJewtG47cYem/Oy0dDxoYCsi+9vekhkF7qjrsoWZAdcY5vknkR7jG/z0LwPcaCopuU/LEmA
h3RTwB1zf3gkxZbJfHD3vbcX6h0V27Qv6OzCO6DNAaZCASI1KYSc2QPkdWUdglTuD9tIU3lR9yBf
giPeLPIIsZUBP3fYK2kM8xAsCEvZwaJceesl0Rl1wZ1KcG+f5l7SFu0n1dKtmI9iCevv+57dHFU/
1sB8MTDc/2eaazlnHB4QEUAC3NovvGQJdfhxDCak107i2vFB0/e4CmRJMDW1U2HVWQp3p6/GSL+o
cs/peK7nHuqm6ZkGqBp9+zHZHzu6kqaM/FqmkX5o+YeKvj2ynmHcnWhUc2QoznPkReTaaaU9DIvY
V+wUOOtijBmEpe7sc56tS36heoEBOVCXoJ6IEoy7bW+n55JuABRSLmt7YJ79u+8a8y1yoj/rOih2
BC5Zw31sJCQ6H2LWpT3sdyPaaFHqLLFC7I5g9W8cxhg/CdpN/EK9n+LAvxDcoC4TPGLypjOKxNw+
uujqNfgWx9NJe/ZKujg2wBHeph3p5SUtkPKyAzj2ObWKgnqJoOkUeyf1LVtMEji0iybnUN1hT44R
0xLQr85VB0hRzPgCQjo0jPxHRzNVcT4a592fFez8sBhM9/5JmYRy3fuCnDPT8zvLL7xu9ACRHZGT
yFK64Y7rsTLwWkP07wMmBeuJNJh9jjNV2i/wgsft3m/NJmUHqZk48Y/1KnatAgjZYxs0kB1kr5b+
12rhppAtbwX+8pjQ++JcHjh/IEidXZZNeiO89DqtRVsEElYpqX5dqYr+NJyExLkAThvZ9ZphsmVf
dtDCglOsPOPRqqxqbdQBGKlCL8zZOVRlWk8aCiMCk1SiwBb9kOJDmOuLu63U2TWw7dSaEWuqY0zA
Sfq0gNV6lbUzLxyA4aUu6yOi0Vk2IzYaiE/Z1fiYLGsS202m6NMvGjC5Xz3Ocp96UW+FHHqKNIww
4SsewZ4D0b9I40lYIj5V0x0Ih2w/zTR9Qg9gCRVyvYpcq5KqTnM8bdgte4jXRj3ScBW4/Zhkji9R
ohuSFuxJvWnDdZ6pC2gUjw3H2TOS3wS9wemsUdxPZBEuGAH/Um283DarOlXLwIrwWYBXVLiB5JY8
bjIzKVcmqnDfX3CCsuIh8dJzP2Y5JBK8WhzXCZS0Dk7vJm9I8XeTxtGFuSsJvAo01wkGfrb6iSod
OAOIvF0pRiMfXffmBkpzuDx0jaMFXOXfSJDh7CxZ+sl98xBBJ+4mz65KwAuMx9jy/NmHi8y0ircU
EdaBIlhVOv9Mg8GrhxWHbGphRlT18wCqBoCsVuRfzmOSHgbCbY9ufqLjTJJQ9fathEhq2WfNgG/b
Gi/me4DKtITQjCcRqoVLB8ZeL2oQ723G4+tJy507Y+G+tHBKJ+YQFD33jWw75q0KOQ5OOmgafv6B
mkIFTvQFavxiVc8quBY5kZFNJ7H8pxzn+Bv9gz2gZIWzPzHcB5NiABgo1+QozCy61y+lBqTRyToS
7GGOrrHL6XogXT6C7UnbTyZd+2JoQD+BLldo6eziJhpe7AByfGyRz4Hxta57ko0mFR5OHUayolwY
qa9V2bY0VwiPsxHkN9/qUq4YGEy9HYe12cbXItW8sFqTuQaaOwagBFCLDvfFxsGX4kkEjzdxUQCb
hD+gXsXddKqPWs6kcqY+DRfcpY91FK4rqnjeFAso+WH7oADuYodvRO3HALXITfFe+pMaJL/s6If9
kNL+oC5lKopoIBFYHxHDDa01W7KBTj7Ju1wo1PkBeMPQNIGmt0C+SmQ2Jwnv0bmDHIL/WJSqS+Ei
2eWBtODaBvETos/+8xu31rC6M7PzQlsbK0UgpXCqRGpp5QfK1Rx2vQc97RWUnPE4fq4LPwvayYs4
yVtZSRhmAdrgBJ9Hjji8qlVuOFNRNk9glVqYLpJJkvF6RZ7iMYnnDUpyKRhQZ7AsZid0jEEtGcEV
iDWTi2w03n7v3xlR/FH1TgAFkn6MF964nxE0bF0qF6PiLMXing3SQHZzPnRpajAKiyD6zMdV2FbJ
zdXv4I8eOp9A7UXdfqxI5vJ1+WZNdUStSg8FzQ5jw8w3NNXNWvL5ahOxhtWg49MhvRGOfG+SWD7m
awU07JAr9CbvZ/7jSM81xQXI4PQWGKU2qlJUvVQWKnjlq1BdFPCEyl86c4njFosMSxJB1o/oVzBL
L6V4MMH1RgESWS+rCt/gSgzKLTvzneoHlw6BexZ6aZ/lql9HalLACJdDaYyj0FTktXC4uvssoE5G
mi8o8ZimXghog3WyL1N7bQUEvypILMzgWXPB+0tLq0lPhAUIXxGbUTFTsPOxM8NC5evEdwM2cf+O
m71QijBhqnWbzbbrBcDqeEmNPDqIEC7z1Wt13Rb7dNUrQMq22k2voAoqQcA/ysLgyHe5CEwLwzXy
6hHfVIMPyiZYejUPK3geZQpmnDxgM9zpsrNhw78LV8lxNV/2kvmIaZVxogQvVw9pcbqQlJi4cdXt
+LZgfrRSLfoxCPy6iZAv7AV8zmfU35Whcv9OKPjb2cBRAWBrTMZta/vHxpCnlg+5KfxW2J5n67jk
88q3u2WvXLs+FmVChamaW0JRZVL4BuCCptpBp6i1hGM45PNfOTSRwnbFxKa0jlflnAFnwYvCtZnX
X+GnSVz5AVCSk4tB6a0semriemjsGD46HVP2FagTECemGfZS97WERmK8PhBBQpCnC7EBgkCGaMhg
chrCIegwuM97Ns5bcQR+M9XlkD8fkdAEqyK6XEFTiUmD8cXBrab0zrhvUw1XK9D974jZmoxvx3xv
DxOVEq2T3eBUJViF6qyvdC9bMX+k8/sEnD+AdcGx3wz7uAaefnUAjn8mF3S4TIhWbTXU4tUlaeZ6
QWmA6xKm36gkIOPPZTT1AUyefauw8g+NTPy9pcIR7vydOTj19B/es4OhhC7jZVynUYHMyJWwWIJj
zECMYokx/7RsDVuP03oHCCSEV55SZa/ApHNC8xL8Spt0/gTfUXC7F40sGVVI2qSTG8mSytWNbD5c
I+WdlsXT+2Vosdeq/G6xXdZVgUaUkF6/COeZ9Mntkyt1/bgI8X/GGEcC9mLlFDf3LIJA4Ge2h3GF
dRcqKAayk+1V47NvDGBa+3XGr3QxXCsBneLSsXf77NixbxevhUTDK/em+jnq1oQKU4YnOWAv0yMU
hISl0S7xq8//uaYuIZ6VGKhwv9D+2S7EDV+RmZD9d5lRpbwCukh8U2NyWfBWBRZlxIEtXRw3ZYky
tcbKSfLnJfgzY8XanJ7pAizFt/bLap7Gn3TGswot2kmU3+WxyUeCVQSMM2xfFQTTDDUFodrkK+UG
ozDGjdo733QW+0oc8TS6in6alLU48nMxfR4TzaC39+6J7NzSNZ2r3cU2bjOqTxILyEPmAbrBd3hX
LXxslkALnxt+RplPFmFIIbLVFrqpBTOMUoSxQva3e3/GFY7exrp+AhZQdSaS5bo8JJjIb7LEGh0Z
laTVD/jnXXNsC7VM57T4L52fkNhiIttOBSOFmQ7yc9IkasJjoT4y28MtALlthU2cPXnBv/ta1U4R
Dlc8bBHD6VUj0GQBh1EhbFDfcu5LwI7HW6I4mKYml3n14yY9YDmWjJZ7yDKR7QomFzOoux1hxG7Q
udJPrll9VDZidADN5ilsWW3AdLYirMj6l50whHdaC/tFVKeuwhd1XjIs7ToC784E/fMgurPxdQKn
LmQfplWAkmCm5qi6KWG5EKPjT9p2JNhCsPTV5bsqZoeGiQ5eHuUeGDsClhZUWBERtLfOgjVG24t7
Lnk2+BsHi5MHb9lOxxp+n1AdSE3MjokKt3aJMk+o+GDjXaGtFfD8D+ioSZ4TPAb3R5h/x7BUOlet
9jKhYzwnI1/mbW+Js4B7SlbFSMl4PzPF7FxvfRrWB4edXApibMU9881mdR9SxteOWjsF59KXeU45
KXLmTCicO6qCppdQpM0ZEMqA/a0Q1F3CpjYmCf7Ceix+KsN7HFJah3x/2n9Yaz17lZsqarqAx2Sc
jp62uDSVR0jBFumXrunHj858hzZYKN+MKXKmbgrfmmOw27tUBEL+5PvtO95Y0ilWPr2Ih7FmfTWQ
ucH5UwZMUZ1nnb1exMoTyfNf4wlHidjSXKqiGoq+ty5NgYYpxao/5tylCm19vy9j/k5YPq7xSPfI
ixjzI53BtPttuncT5Wbqfnbvr2hTBWW7RFxR3EoMh4iVKXU7NEuE/lG8Lx4ljTkPK34cweAf7UcI
g4otfBiuGKgm2MZY5AhdGi1nAAg73U5Eg7yxz4hRkq/MWNLN5BP2K+5ZEb0hRVTbrtnlBBYhxQdQ
QCYW7ezKJcgd0BFu9A6jsF+eN+1nnAmeGiwAYn02joBRvgET6B4v3kBHo3Sw+IHdiX9KsXFUgOO4
W03mjplCA9J9u2+Wap3ULpjNqdXnzUMEdV3XQHOhm6t53T57mnFAR23/K2NDqedc9OMLMLqA01CM
/tIbrKAOMavYdtSLtx+sZf++PmN5J/jbiOJHRrpmWZinG3EZ51dJonHJmihODMUp1VdrCH1RrhfJ
BEOGTBQL227dHI2rgg870sZTxeu3M8TrUwmbmChDwJ+tamiZJDDe9ZAwkB52oynof6cEofSB1jP1
XVjlS94oVeui0g119LTz1p1vyHEsW6mPr+641YcI2QuGLFvWZA7R/uilIQggvlxfeJBjOGbPCqf+
C92MxXW/hRjD3Rfk+AlMDu5xn+kZfSWyHobp7lXYaYaM+Sne+Gi/adVYbCLwSIwVylYfir0Z1ytN
ixUqYgujLxK2CwSQqEKWIuxGrhmnLHPIRkNi+mJE2VoPuH2TuYYYQZ4MX5bez8ZAern67oFJpuw5
F3qjgsMWMtZEPUQjMoTgo0cZUfNhyLliTbI1/ie/T5hbhuLC4fb4upknbwrWSv3BkJCDDCr3DnX8
cz1C3/t3t4kQmamiKw3VHSDRuIQlSpBHxi7nvoaOL9smpVqrVlR8sjhkpQt4pK0SiU1tw4+3yqQK
t/26xS/1jKmpDL7R/0a+tytfw22cldxGOW6j4sohh86R/vXEwQh9ugP8hkScOdMGrDOd02nZAtyC
76kPfqyl8dUm6rcO0jkN3n/urX4MMDEMAEnREeRAjE/5xrkDG8VvL0FvZG+pxxbv3LgaPy2kRuBQ
u2SduwjzXZxSbFINxa8mKW3ONiNUZW5xuwjO1ZJBs3KajlrAWmxTIeNbg/5V0ffciwtX+t6weF+6
STpO/Sz2spHO+5sRAmKJ7TceczzE3ylHxnbX9WIb1IZWcg2r9Ye1XBxoOXzZonABJyU3Qyv2Xxo2
fPfPC4btJK6mNORuxtQQXshvflGu7IQXrna5JSCyubY+rvTcSDE6iPRflSUygaYr0oqW+OXC7K3x
eiX+e122ZgJIS30uzSv5Y956G7iiFKikDz7gHta/4tiqVVLbuyvwefz65A4G7JjKzyirRjakqudi
Lz41fiil9vKQJ+Ffp4AEOMhUxvq5EkQykojyBjm7R8smWZ4nqwvpqMb7bxlrLUZmhoR66Y9gZAFC
FkDgV5witNv4Ajjz6Bh/VM/YrQS90i/24LIuMh6oolc/oO8cBOVxB540u7sioWEovPKvNlrvMbZt
kkws3eQrwGgPxPHW5fYaMfauEs7sJ3YXnLo3R1kd4j85QxVH/g1DnMSQw4507nZuEVaL/uDKquAW
yAQfHD4lIy5Dm+Oy5BPoFYYxovzfBjZFFbK3THYWGprSNWw/nOo2ildhfH4lLgi8xnc+JzLCvlbp
snQS26fjpINIlA693mVER1DRg4bwRYRTbYH1PQWQnEQ76VTku4jkxmHSQDuNEcB81kCGI+lo+DCa
1yaY9e019oAtovce8zntokZN0nw4e0R0al47tw/FOJpr4CSXVvJznEbiBnREA3XNHPi55Mf4zdqx
u/kQbawTiMH75beognnAaRFA7Jqln/axy0PDUjtLoUa7xHttPS2tmnQ5uzWwmtKH77gSc0CtmzU9
hvHYM/6VSL/kXmN4paEhkJrPXgc7ho7uGqxQCWcSW0Gb4H4sbXpcrRZOSszUZVHLb5lAovOajWoB
Zu/KuCTpQIARON3+aM7UIGGPMUBF7pcGwqJPy+JJGLZZ5rrsVnrwyj3aOHk7hqvii3y/QaVNLtD3
xJJoxk2CasJffFc3oA2mme6nqZZzetKfGXKIrbJuE1K0lNSf8gzHP6VNi2W1nH3nE1Wqjmj8pQuy
p9va0v1efg4Q9tjARwO6S0RbxqBWdgUa7JpopPArfLBojYfEF8PRsuaKw0P9EWqMKCZaxYBXXCWp
rtva3ZshIGGDAWSX8h+fG6R8WmJ1okmJVAtJO3Y2p278v/QiqnDhd6u0K3VRVDvtJ6JgcACEnvEl
5Ad3iB0ZyhRp+SSGIlWze0bqvDIJ7IM4k/FP0njPBbg+GmwKEIpT0C5wqtvHZ353CYyFitjZfH+S
3tPrVpwZVgeH8wa8MSeCUAEjE/0+m/P0b6PPGUHJCULI7R3bRupQ2rCARhlm6QbQT79QgKdrcKIq
OclwdmglYi+wdDgBpC/furvLpym69qrdSUjfWjZDWvBV+FnrGemSgCg36UNVcUftPmEGBmCHRNiC
gkyA8GSTq0qx39Gy7oOi9MXLnXn8ZlqzafPmgAIP4v0uUJrYBx/aTFJlZz1L5BKjkeuTP8UqQHri
WUynS1XtUmjHdk4USJrfygQVVYcthRAdHnf5NjOP7dt4HcsORnCMT+85Y3kELUqeC68JubNnedA+
x7Ve/NPF17+6MKg+hyxh6Mdr6hZyt0mK2e8lp8+tp3q1sJyPJIDdKAODSXN2wIgkQmAAKIeINtjU
AnQKqwD9L/N9nQaBiBa9uTwjEjZwe9XtKzNh7B5Plb+ODDLWulvUy4OAEWA8r9jIT8QkWwi673Fb
djThzRSV3SVdARbTor6Qn6c7kLT+DVa0t6I9Jl3sh7gu4PbpAHfcv2JiTcrETt1a1N85GPT89f6h
6BoNfVwDeUCMrCDGHLz50s5z1FgeBWP/crhSO+nQKv0ePNVFIfpbArTSiaAipRPHzzwGbH2eNSRR
BsTMgM9lsrZIPlpw/tOfMqTPfFql1biqMfFPKqrNghQO68saup7b6INnlOTOEJWjMAyAp+YjqsJ0
pCVF8yQKSgMfr28pCtY3mrOg7NDC0CULlfMHiiPRK3uzflyggCq5FdLWj1NhmX4bxoIpmpZT0+hq
PMW2xcuCBXeYkiwvpg4F5+t1rSzml4Vx/uRyDKNNDUKfzxbCURe+3L6fUS8e39NqisEn5eSRaRHN
i40z6hXpUlLdAaw1X4rXrJmCyglW772fPjQMTArszoPrxRioIIEAp+X9jM4edrGPpEFebHkUaIpC
SLE/xxG+1Y/YCndm1D5Gt0GnoaLxKJ0fdBipwZUsg9hiV11oT1wwbbDhYTLD4ewTahMfVwkR9+ii
7R8kQc0RKgUxplw2a18IkWZIj+VB5MunpnN1PIICFRdYLEhOTOUoVSa9TsUa5qPT7DLIlhZxe7N5
Nr96M+3z6Klvw4YI4pIk/OpwAsXKLhoU5jOFJdaYmlzCQZVRLJFht1ARMedsxHdDwXgVJwSmJt08
6nBizjyEuaReQuJlArk9HJbgsbacQCnvAU5TmdmFCvkLVTUJ0vOmTuu+7lU5oK/Ho5mBHrpPsm1I
rhy+9ufvKVuPGxUHlMQKo/XZKXul/aF0KpDPgSKaB2HGKfJqwzW3GsTMDlIsWAofZ56638xBwLRR
ZEg+eU/lTp7u/K+jRESG0ozm4Gpn5h6DoHy5E4I/iTvFDyzBOXtYPR8dVtOoaB9eQNcJGiALzOIY
6LEV7g3AZpIxpr3I0fuxjwlTmfK5/IIhNj0uIrfQdiegK7yPi8ItnU0GZPlfL5Cr5kxpBcbsBgeo
4rRzC9EUKl6qTygXVqV0C7ODiu/ytEjGMOMuA/3GwOJQwolzMB+znYIjIr4W8AZ9z03jwa42hJEL
ZhQq1n1KZ5bhl+4z5tMsI2uAxlMU1jSAbGbpYnTSP8I9zdjP/l1HQuL2SX7fUTXVB9AsaWhzjyCA
aXeDiUgen1GFEZ2Y0qnEKB5Q9v62795YOYDfiq7r8KrNiaAeiLrjxbvuF4y9CGAvnpklX3U6xRy6
wKk4AzHxHr7z8/y34KuJI3rhNVYaQx5kDHV4iXoSDTk25PCMqiiHU7P6AKITmmTcApnzI6VevMaG
ljTMiA7Iqp7u4zosklgXXc8XIcwYCnfw98IPu1eTOelcPWgyr838z6SSEESYzBwYvBcUTSpGwUxP
MPfkt0Id1o9VQ0GQnqg1PPmlWjcFpgUoG0/5/NMW1i9kOTopSUnVuTyzT67PLevDi3XF2XVRxGpL
/a7Y4TQId5rS7fH7wYMvrprTl+YL89xkKG1oW6cq/BZ6yPe/ncgthKExox3j2f6vEs+AKPzBho+r
HQqB4dYFBSitFsQaWhC9M0c+ouJ8PBgWuMJ4lCGEayLVxvk5SqrckjDLzdCohD8p9qpLrwVUhuSx
qmutnbm+W5OdL4sCHNjyUwQU/yMpUuoqmEY46OEOQO7WHh15Wd09pLnZvdbn86334AsaOY+PQRZJ
v9R+/i9WaAh3O5JGQGJuMZ0d+qRACf374BOzzIoICLr0aP218WdJCxFEqLrg6nIn0c1e5cXVqFSn
liHP5NalMTyL4Zk7qmRV57ggJEJLrn+Ioun6r5xFN73/rcbHaiuBnIrkM6LaI5MRpjgdaNTs3TGE
bWmtESCh8LWw2m2AVHg93aJVxlFHaafGxKm7usCql+LT25ULK3dENYfPYb8Fge3w84KHjW2140iL
MO9nwr5ako7BltuO5abAnVm42hApiq9xkIe83vUpJbtaKtMflqqsLk3L10zYLkwCS3CjbyGrm1W1
N19bXd4t4NlgTksWTSiJqmZoDfms4DsoP1AwoCpVI+gQf1VWTVNlmU4dEyFtFiA0CrpjrKcwnBGC
WBHsT0lYo8VGO2rAq+ehU9Ef5WSVJRVVQ/SCdVikcKcv7Q8lHG847ERRDBq0JNYWMdej56apFe/9
LoEmQSFCoucNcdKlGnXV2q21aQ45rfho1sf1o1WCcWp0kDfYh5lNTNkwGv/lnn2ekzl8vOKIgQJ5
PppFVsg5g9hOBlhS5xicb7R0hJf8KI5AHitnKUK4pLyKUqExl6JEQzRqYK4eP3UDmJvavLjSKj1/
lSY+zOzMGeiIlDhyv/gj/ppL6xZ6+ymEtrjOOKAUFA6xDw6dAV2GXrkjQgXy7p+LhlHL9RqCGm/G
pEGsudNlD+74x3P+ERKwAr46tbUrkU2nIc9mHNCRRmpXmbQ4lS+1ZM3jam1dqRw3fvummoTFn1dF
V3+3FV00KKQrUmACBCw6cVfSu8ZS3ovACwMWFAkQmiMJJQnQel6173EGz69bKGQpEMNg1wuB2GoX
7E+GUbCKapBKkY41njVjJpozGMMvhO0/tE31alRsvCuZIMsipTjpSgl8Qq3nwwfSJ4PukNgjlx/S
rtQ7Ov3TKWwClUtFr8fd8gzh/NTfqp4h5U8AAxZA6Dewi3Tzk6zbQLWhHEPhbkYITW9cyM2ZETM2
NTLr11I8EZU9VSPSwgF7PoKAmOeyVPpol69QhO0ue7mbES0nlS1XYLcJM6/M9asva1qYqLgjYQHV
HVtBNTUYmVLj7tAZ05DnsFlaJWJYfNUFHrIWS/l2UyeK+IVn1TGMji8w4pkW394eUMVHe1v/9Wy4
jdF8vmpRic8h4RFoK/xTN/dekNzR5EdlyRufIie1ZOxyiWZRqiKw0KP3ayzFncWSY5alm7F3HL3K
zl7NTMFWwmSJV9nhEqNE7HwCn/sLaMGPSwJkHNRAjcIMNGr++fUYtkekSm/uiOUlM6R5B6rVnEit
i/Js49tQJYpsyImP2mRAJrWlpWsv0lbzIZ5BtOSl7pzof6g5D1+9Dnwv3mWSQOh397ZaCCq6TcB6
NWuDWlAq18ol6CN+Db2I7ibSoTntlTCOhJqH4/BiFoBa2p9moHTTHaSn9NHSeDMPOQ4dz3ijltxn
rL14jQiRKBoV8T7yvLnMGhZp4d+9wQCVXQ8qqQZCF98liUCsPOZm6LDDGloiW5KwR3lW71J5aP+2
rkS/nYVTCmllPZk1+kR5DJDvssd2olCszr1D67HQ1CUSIwQAsbyu43ffY22HVQZk4Btu6Qe/4aBo
Z+RSWxdqmJTabVG1Jczul2BQG8mI5yswYjnS+iu4oFo5Foz5fxrErT7uzzYkjbgFnU0BOIopHNWj
hs1DAt1lr4st+xG2NhRXaowDprNpm09sOEZ8cKA/OTYpC9DWd7wnHicciubgQSioKv6Xen0VtSzd
hJ+4ywhMHZxqw81WK2H55fJvzg6dZ9wuu0tuEzKKUU9zYKp2sYh8xyJ5aIFRo/+vSfo6ft2td40O
aHZ6RNO9Uq3CWYH/naBI5dKHem90DTs+Qad40qN/Mt9OrEKrvOV9nxrbmRqCNjvaHvu/xnZkGnus
ThRsEnlz/inNxaCNc0JBxI6o1pVt8HulaM1ir4AxEkmPaVBIGPWFhM2eKl99BnR0Lys2jVBXiHFg
W91k7B0bpq489CP+QL9lRwGl8NKTczLBd6MX8gz2WMHO27FxiuCYY/6S9ZMN7tiap45blPYVQBz8
9pGL2l8Ghx2wMHcTIXe3lUKKtIh286lCxfSoi1GhMXnOYrchAfO7yDsTHxJTxGDTXdnkMaETCB2o
dPMjPH64ZSeyv26SkA5OpWP1A+0icUeTcHb7+wBmmOhGXqv2m42fHkEo6XO1sF4JzhGREZL+EDP6
+DjOcBrMDcJ8NzrHbZlkDfrRXKZ9NiafPqcJr3aULuUHHVXeB3PhWMY7wtpCvG16K1Q+1bYQ3SrE
ocs+gfuh+b6vJnQVDvDVc+PwyV08reELbJc4PUPrFg+4ye6skbFpQ5E+vTxmYnpHfqBmTT5MPM+d
LGq7ugirlgeV9ays+pBsleQz7Uu4j0CGx1fBi/UB/04BPc32LFuDt1q7eMe5g1x7JS3s0DZe9kaB
1oHC2/ZJW1/nCFrMhXegwSZab/8xn9l0K3M9CaYdXQtVwHcac2OYpOr9wY27Bqp7GEROhriVNRmd
VNNPvI12Ke7Q94XpGX7kdFtvJpiKI4MwhSHTEQOX2ECHK2BZNsckI9KSeCjCRk6l//Ia7Opc6fHX
TfxxrM1VD58nzM7C+j2WewGFYHICz5Qwm3YW4GVakT5rQbNLpe9s6RZkEsFCDyksYAhp+FGZMRlb
fEtsWixXFQG6meFHQGPZKKVxFGq2/8c8Rw8zozK15dqsAymEuc6iiQ2WzGdSuyU+87GFvnS67Zir
taT/TdrOjsuADXMSfgjnrcQiaSpc0MUtF57mzjDBOQ5jpowouErFF9C4SD1d+BCKGfZwQ5TR9kJr
Wer8g+EvnFbfMrbclSt//HQfeuQ9Cypd5AT0O32oivLYym1cBg7dDsQ5jgTJbpC+XZf5K9vl6ck8
TFzei6/eAj73koQQ9I4oFrv0lDkAauxIfctZ/58T2Kp2daXDVi7PQQj5SDE1XZYB3+cZi21f8Oq3
kwnbFtmCsNsa3f9+VnSLGXlLtQkyI7yAyLfwxRa7x3Dy8Oey+rSzbfufEU5T4O0i5F+nDXZZL/aU
VtKQxj46XXNLOY4H39rYVoYZa6P+04RMuHYw9BFLin9oYqT9P2cyVDSLZMYY4SJ6yFn9e69X3El+
m2JKYlP2VgIIJZc+nCcO855PAOCIZnr7/mVACu09mddjm9MU/qzb9MpGJ5dciNi96kWwPygUbb8S
7BLpsyt3uPlyEo/+buPUUY0U0fRk+5TnOHAn7CzEwdvVCK77GrbyEd3V077T+JokK3dN46LshZ1t
BydZLMrR5e9Oi/yni1cFqRPhR1QxDV1/HrUrDHyfcQf+sHKemNM4kW2UQEAWOypVcJS8+WJN091p
bDYNGzvE/MB+092FQCJbYoeEdFOXUv79r3zYU3YTFS/b9KKwNVwmmF31cxwFpXbeSt8rKP8S5cG2
/fQ+ETN2I4yvxKfMQhAxd8zUs+OSVUcjwb0lFs9iUhCknUWCljcd/JPkPRN1BwfoXnRB526cYLsM
U3UoWnjAlzet7Ope7WtDYpgs7vxePRqiEkByqPCpHrxg9hNOPDo/7vnjttl7w1ABvb1Rv6QtOtzX
D19hGXdaps53BNRL7iAHkj3F06ST/xmAjA+i3agP1WLPFS6iNUDv+uRqdetC6yUJ+U70nAcYmuwS
joDMMiIGLmAO1jDOv/CieAHl8iNs2DrlTg2oab9F8dbHu1qNTzvv81fyKeh3TEk/LvzOkXjyZlo5
A56OQTu3tZA1984C65Le4MP/xIn7ChBHzYXTsQqV55A6arCQgadd5RMWJGqCnaPQu82cOAu25tIp
obQp1SfISxC5kKCdCZRakICDgEEv7ZJiyfnNrFe6/ZgSUC4SWK3RCtKNbbQGAB4znzBGY6iSH381
hMpRj4IzMHy5BYCkM6pgf1jpXsQzPNR38EUU+9LQ/0BRkq7mUR1ynQtdez75N+JQlE/ij1o96f0l
XumBMPgzDnK/LFgpcUdtV1ikHpomykdoF0wl7vaZeNe7aDR9MxOl7fdAKlb4OrvX1XUqAqvnjElU
IsevcDfDdjoUet3MsdAsVPkb95WyTahmz04925wi+t76OKo+W2KPqIBzsJqmRo04KcUF8JqXGlEZ
NHyNunWUF9BxZuM/r3uxkx/3GW8TBuWJFGV0i/+j47xKkAhdmDbRCesKUSJsDzfMWKsUNY2pQiD/
gF3EyZ3qwfvOxQdOC8yOMvc9WxAI+Vu0LJml+nvdDyY/Iz8TKQB9iCG7Vr8+aoZAsIYPJRx4TmOA
8mzhp7P/9Segll9nJqyLBNyfmsaeAniaFeePQfj0+QLTXgB94j6sWGEOcrb61RVcQOWhsuFrzlLD
k/WGgyh4rLqJUeLM3418zWmJKarhiiaRyPz10jIGPq/zmjsc4AYja+MKcEvVxvOiGyCBMJ+5A6Zb
fKlyLAGwPDnTbZ66DERP9SBlYoPNqH+hQwiJ0mCYYCaLs4mtSH/3WafH58TatG3KW2iW4pkRE9PT
oPH3wQ0LMGCnovOemC7H+mgaE9CifUKpV9OkhpX+eqZ4oDgD/tEzFIfgwkpQ70DoOANTwdpUkJN0
vfosNUlaNxM2MJlvDUSzewFv8wItGOu1zJwvJ6o+Qt3OkU0SMXG5Yls/cHteLuFXOX5keDwJlq2m
4Ht9DFr69LxBjJGKygiEO5fdn1in6RPnOBijlxcbS2bA4K3O5bXjGGbPnLAIqNA4BZC5AuK0W07Q
3LBU68zpYzC1a8DRczGMIIciE07QIKAd7fR1bqyQQPdDk58BpL4fuNHR+vGssoZ0DxaUS34EjvGb
KzLmQFF23+LN9pLpRRp/RGbZ3nR+q+rtpbYRgwh7JsiCFalfYWYYgBeXLY3XmLeo23LngGjJzd44
z8TR+XeP6sb0+ECWWwX67nZXJg/Y16TQuhv2bqp3kG7yg6yIUoBMSomayzSHyykJF9WsdO8LUfGc
rUEvcZEQgvhSOtCc/d5iq2rOA2YeewAjha8wTSPjlXpTufZq8crV0+MGozNSdse3e33JEZJrdIvc
cpHiMNWZEq48Ap8HHn4JtLllRQJhZLhnZolGauseH8pGB5Ug8k/zZJ3ztJhMUgc+vxpU0qxsTjSh
CfMu2r3a5Tm4qNDpxOysxO50OQ5VVrLgcWlr+REQHwA0ELx1oCFG9i8qSgsk85Dl02U51tyKiVO5
M1ec1OUs5XUunRWs0UEg6fsfNrboZcllKAD535eWDv1LpuYqjbZjZMuElGVW/iesqy//wJbC1Ut+
RvMmpvhAAn9HThlgseH1PtKlU/ZaQdJcH+UsDF+E2dPFOkzSQ6Hn6nBBbY/s7J/rvtx/2S3BApwe
/CPpIWyLMuWxdaeLbxLA71JzviAo1vOHz0jZnTqn7MkFcIUe43GFZzLocG2DNyJCwWv+caAd4yAi
0rRJtq+sP9W/x4lJF2pMKAufyxxFzm45s8FaztVi8p6uyP8GxtCzk9WQ6eI9FFlHLk1hP7dhq4bP
IgYYILdEWGTe3RFtqXqHDFVBfehl0TXYXog33K/wnW4qd2f9Z7fQWl6RP31mKaGS/KWWSs6gZRFb
Ts1fO4WwRKPv7rCUcLi1op9FvAUEuv/JrWW9G+wzXWBgWoOSpPEfvrn8eBIrVYojhf+Cy43FipnG
UQd2cgswR8gHLDyqdSomd4+VZ/D5D8la8iy3Hclwxmc0Q1vK0CY2weieHxcXwOBllIYuUIqmJ9cS
EOFx1Jp4lyTVRie4FafkyWnu/NUHfXgIkv/Zv5jvG8EG/WgIvi8Qv+R/QB0dMoboQz445OHw3bHK
4XTEe37pD7DRIFOS4UBM9T9iUYgZ99+57Oc+NnXtnTyK5KMGQcjzGwh2scyXniuDUTeTgebjkbkV
kSuY+xBLHTG8fAXo+/vbkbL4sGJBdzDRaJMhyGgVCaB6bomIDCpY7VciIOyKjgeKd4bR3heRnFhR
6pp1mHjYq+BPmoZvJXZLC15SrN/xDuLXZYw0sm69lIiqmxOjrccwSplwu0aXSFW8/MWKG7W3tqtf
c7cEWuAcpfcEUWTF7bBxqr5yKQhYenKisTNsCZdi4/Xu8h4QbAYvM2gkISjfRExZyw1BuOGQZIP0
/bq1yvjwWpAwP8WrOkdFOkBonsISl+w9/AVT91JIaLarYq7AriS9aiw5eUHZpNf6pELTG8ui8dCF
1cWqX7O6gi4Bukf3jaoSQf5GAkRhB0RpeShm7cVMbZxNeXQFB7BMK+0Gly9JTj7VLh/lZagpfa+8
m1H8y/eJJwX/acnDwdWNKtvEP/e2pteu/ZreiuEOupYYSoF5CNEr8GC8ySOytxAsVwiQbl2H/Kfu
RMBhLC/MW2Q3CwEJ0610fu0V1akxshrVCSlJ9PxyPFQddx/qyDyLxx2kReBg058OXdwNS+uxuum0
NlgOZaWmYs33ai5cNOlufhdIr5SCYAwDDRoXd3l26riY6/6X8sBEXxNJO6zXbzAx47BWLASdXmSH
dWjSKHXQPsF6oxWK2G8a71AGAgwRzTE0Hi5rGP8RgU3QkXPfPlsah9vuJj+lVJQ5pdIXA4T0Z/pf
X0Ez4yKHtH2jIUsWXFJCdC8QLbd7jNcP54Q0pO8jYhrS3y+dU9bh0NVhXq1LNnCBmO980r38lVoB
/odLQitqUVHsJSfYaMpjdTcSaoHoQkWuRayDKVrUekcMmQTz+rZnNJexGStIc9Ou1aRYgkQrSZgq
ujcsF7JuUZ+AhhBgzIO2s8uiXDMLOGCercjK606c72D6ihUuIEHtDJQbDiBkQ2y0oumXdihgrSvh
fMO55D0Az6rk/E99rrBzx2/ZBwwosFtqj22NjNSOUbne/O+dgyr9IbBjLTawOLhse8hiMuOl0pnC
fvSlxJzx89H1oFdif+edHp6GL1tdr3CQLup2+uq9+Cv7AdxahREsaeyTaLG1h7V88Daunm6IcRbx
VQ773CVnxW0JD6GzRip6p2ZYsVEqPnN9/cNFIJgP2GCzKdXq5pIake5rkYAbVcECJ9CAn2VRpriV
Mbxgb1n0mPPVwfeD1bmJXEir4QHAfAiNaeDiMO0z36E9cMWqAw3xrVYkL7/qYZsxZHk5C1a2mU+X
Z8vQE9EhBop6bNtsSAfYaKru+C9i2re05BsA5HY5ejSO7zSwkiSUGXWGNMeHpB1fS5GLu7BiMF/5
NLemfEq9WTc3/+sHWVmREE+kg5TJc5EoYk1i9hy916BO4H/LeCKGPotnBe0kryv6I05UBZM67oku
T76FN4h/iBqK5PfUs3dl8xtdcIBjCKDrnOcPlgbNbgNx/Bv16EjRBwZqWbEncHmenF9pgrj4oXA0
2+bQUdOlJ28g4nMx09y/hYoUMytRNqmEkOiYMPdPlYeqz9n8TQd9i2eIeow1h6DgEaxQCiBgkBzX
xzOxHHpOefahb6p/no4DVvl6qiJaADSeRqwtclXuGd8vF08eNlcmjEMjN5evYz6NngjmmxHXMM8Z
W21KkRVWuc9FmaCVc71yZWzLK1ncqKdstTWvAHmLmOgDVIPpyqHYMEzAF2wBg0ZdNauvo6u4o6ln
icoWbKo2EXbZl8ialDN/5Ta9bxULpt/R5VuH6q7DvlkUcRKJu/9C1RY4ByjHZLzgL7e1G90xRiHw
8YVJGSYGvMyrhkk6BxOYdnlEJBGwI3exIxcTn9WJ7gx7Z97V5dc57oVK1Z9/17BYDcgbL6WvV3vD
ESp0e2CcNRhOd7gFyqGHqy5LKuNo0zrekEfx0s26VO8MfHJAxkfkYieRtIUdzv7Yju6JuW0Ozgru
0X4fIbYhpFKQ3TFnoobmWT76gMqMnHwSGsXSqzZobCFRn0hzx14uVssWe94o/Sx0+rMEACLvmm1f
zDRQrYhOg4sEM9slbAtOXIahZP9Ao3WeKaWeK8ohOlcxy2UBm3E6TrxhuaBnzS6PS3cIFy12ngoo
nvv1WqhPj/qgRJoUtrBTZ9mVF8JWHDHVoN3JYceQV/7TpEN4Mn0EO4ZA7rfr5r3Hn/fl0VgiDZpI
qeqJo8TntMA2FuCRAGgYLBhGB5WYrx+IX7Qr38yUsJe8mQG3t5mvdynTEMAM6oi+lMIV7dRVKf/f
asZcqGFFN758wjx3RMCn3g/HqIBKq8Du52xUY1kBcUD9XGBnTk1c6e51J/OHXFNYgDzFXliBbFIV
wuUaNUcPG9H3YbddQckW1gargh0cCITU6Zf2qnDeutYraTAZNAMOjzP8OYxnjf/hroSsQk+wLugA
HLfCkXYMTOsIOLdpvWEnR018JXLtqJXkPZRXNYut/p0a9o4Z52LKGujw1XOiVxI1dBLv+xczMaKx
XhZO5hqw5nrYJQ7bYTViftL6BlDQsHV/KyTKnFcAi5zTgV0v3udVrtwOmfWjuYQHDYX/UZEksTM6
6Le5Al3hVM0Kifnl9JukV/g66CNLD475Beutqi0w+RBBcyh/kN5W3mBk135TYBKUsBkJUS5Fgjs2
zHXByo4EJbQT1vfVX2ttiHpfbGyZRgmdu5n1gS3qKwqDHMrYS+Lk8HaqtNXtTGg2abiMSMH74rQN
a7Y7nN2feupTRF8WMwsftpcaNnwNt95Og422EamI7kt/a3ENukmmANnvjSoN1vac0Em+PMrgUwJx
DG+rcQ/oEyU/KagTF8Iu84z+8B+awEGlWXp7qw6iB1626i3cUeU2+17pg8XvfCKa4TmK881nlDCW
7gJOdKcUzG4d4L3AloPu4xaIFHtgGaHbqFfINVHkAPn+fz4QIfsbddWTxZRP6WS5zYu2kI3TASXY
t0JX3xerVgzQHEszKc9w+lxmmM3UNKoSkMUsS8riIB61E2AtAim6P1GbjPvd7GKiLLecD897xlVP
pL5/7PiKQ28Mgca85CRcKbQJnllNCs3gYHG+BC80GsnfKlN+llGTfNxQZE2grAKJ9CNJ7HdVZtEn
B2mtUYBsvR1DBMjlzsX6VTqvnYHB3jcDL6AZYb5h4p97gO5fquCZlMJQRbgGC4VdyvftQKlYj+CR
T0Jgv5+Ha+A8YeQcNPQqoFVs85zcWpfHw5oJKLb3IZpJBdq5uogXdG2v4ob1htqGadwYoG1eRFf9
n26BwoB7vKHYnkgdO0ntX07h3Fpn66xJdpat8zNPbRTH7qStfGg4RRZyIOhRVA5Z/84U6GwqU9qL
4/zkGxq0b/UZyX4S6sAreladtaTBBW2VQNR30zgHkE+hTz0yJrZC8cwWbTixrzejC8V2pB2xn5gQ
QJuLlAgJJBk/qLempI2iRdnDFJVB+nqKkn2fbemmILGeBw+c+82r/qmg3R0EvfPzGohp7a5UrjBs
Vc2CkTWVHJw5FHTB273ilDxipnjGIgff3p8NbM1ciWqkYjnbqfBzPPZuf+VWXTKzc9wwA33sF15n
wGD0KAKb9A4XVJdY6FX/Rdydl+qBjelOcjaG5rQ1Ja0e68CKSz9TQEC147G9RDcpc8T3unldwF0b
0f1rqs0Z3ghJkn9cHUnJOeoQs+6JDLmaxedBpFMkwUkWf7d4XjL+EsN6j2AY/pj+Jaf1I+nuMTb8
crKhZbVS96xVwfOtGhvsk4YYaQHkTAXjEXpesbul4T3DV+VrzdMvf8mWnpqZia5sbIYwguU75xt2
6biaHTSTiJfAB48lV93iVDwDm4fCwyPWE3YVmffRS63KOEtTVdAZLS6IlBN8gB6o0Y1WvQbxk701
IDjsyayBXyEERtqcFKpsYwoexlLLjfmqiByWiSY9uMyoU4j1GXJ/sG1FLjetloJfOeRvmtGB1+2q
TIV2Mn0iciF4ssa4m3N0bhNFfPFXv7HA6JkEPmiA797rfLYfVFEvwDDqo93C9BzGyMdnYgHym31Q
CaVd5qg3rJ4RKKG4TfCfR0yDct2Wg4TxeoA7p+vdPcu/jGlwwVYnAEXnI+nmUjoUZG9wkdzxvsC7
oqlaGNwH52FIf3Y9IEeWiMOTB8VXN100l2+kQqkRzH73zusjKXKWBdjmB1p05sFYjogjiz8FvGeB
PmxoPTdiKPBWCOx9SfAUAJYiYYoVFHMq8WytzqvInNAdV48hD4iMtfiNTpA29R9XO3TfHizbLiJQ
/v+IDJXROSn5y0D4ZjMRz1gaWefMp9WerObSo+QpBKginZy7CVQs0gY5cXMtDNepA6oTKNBOWqBI
AkIMCmdAodjhJz50GMNyKaXEtjb3uIZcCTE43KzIMJ0gB2gR7DJb4u0Aq/tJokmbamKtkT1ok5TQ
sClpoDwmTjd9RxsJLS7RP5WcHg0cSqIBdCs8wUy7ORTAnZmpvpcFX9GRJyOfsDsvjtzLu5q+RsUJ
NDrvGnZW6z1394OhlGb0y2JP+lG8i9fry3XQXwy+z8s28tlqIdmxZa9W8OoMhI/qpTlD9EX8aebG
76TD21F9Z/wxtuE+wh7BAgL6FOvAA/jnLlrFgnN6rqDKd6sMxGz35FbReTVdO+CE+/3XCwIl2MwU
v1HZxSDOoimBq+dR3I13drN9nxd/Kc0ersSl/VwlAqUsJGBTrlqtFUJFS3YbI+YOQzuAAyJL1Rn6
J2/Pcphb49nODXxWSWATexIqEq5VKuRAR2g5WF8DheHyn35VxPrG0WDVagTim9fsByQV15M+U1pS
Bf5IC/3u2i8UtVjC0g8LSzsnUs8tU708Xn+QoKqYjcLvIi9fMsgV0DRND58c8N9BCKGAbrjL5/1j
L4ofNo5jf1mhT25iMTZy1fyIEvgSsgYXqJ49CZSJCQiZxi0javL5wpDkG2GqYuqTHDkl8xbx8/dQ
hMBa1OcK/X4Czi5VNhQxFxzDGkxxuT36OMMXZiG5xpgB/U+lSPEMmzkrXE/WHuSesMlS8x/VG9pd
wxcW0eFWQTeA+YQ//Cv9ffFU19KJyOrLxBYT5iDmYfsujzHIqkcFjqyKmsn/xS6jnWqGxaHxBlw1
NlRt1Q5QT1Ibv2QHjD3OmyVn1pRkrEJW7y7O+0jjlhysnFR4PtskVH5wAhwZiMiy6FPsx8nrAj36
rAphMYmp7fFcbg3GJCfv9kwtV7kRDplBwZqR8naneTBOhlH6MCb08qzzsuczowPIuY3kFhfiB0lN
MBNPUH04icnFX88+i2ihTtQX9DrsoE1kVE+WjF6/ITIN2hf2jDFn8c1VvQreOvm6dxgIVl/dRdtV
YolpqUr5aybXONQrTm+sdan0KbParlQPeTHb3VMzJGpxxiL50M5BuTqFCMSkz17Jo7zSfBI87wn1
K8E3U478b+ASQbplPPPn8oyeOIXyiPVCbGG05dxEMtOInuYBAR9DkHYHWVUw6dL9HIPiXsoAm9pL
OunDf90wx+Mq2uVManM8egsbhEbz2cLFNdePC2WaI0sQmQLuJvDT2GQc5cYTomImphHR4afrjqh7
Ez5BEF/eU/Lh8ymIieK/DbpaWgbEBTLhNyIZencm1gzTcxqrUUOqVFAeL1V3nn0Zbm08Ogc95J0a
nmTa8qK/cZ/8Y8hkcTmnoAAwxCFbeeEB1skRljXguKb7RFRk/CPv+DIiVsfEn7fEHxeOhZ25MHec
eh88g9KXSIpcpgktuSiC7IXbirpySTYtRnVgiZZPndqKvuAadBTMCkQKqI7G8xBcNdAbhvf0gnNp
nuT29UXR5PgHhFFFLvo25Ww2ltUsr6p/8SqS3Tc3gvq/zaic26h3IAFheGpzrIp/TSubxc+mPD5D
fIWQdL6SlxrofTQIgSzFUBIvILL2ZshoBXTtQBHg4JCSPoV78zx/Qqr1qYGBEbe2DrgEHgpnGWCc
Q6qv8ugM1KqKE1FPfwExUAGZwJKySiszf9zQYW2mVPZBro6EqA5/LXb8a6O6A13PzBqQBF1z4x6x
2KsA7du7HEJLNvC09k1XpZDdlAGgULQZIPlB0NrVEyuUE8nrXtnqdjAZni3gD1rIKnuXUZQsHlly
zRVTDQDk6ulVNO8fvRes09NSUwMS87mGMA0XeKs1dc8DugrIw3IXCA5i8cNB8tMCn4TQkMKRLEfU
6hstvgn5ce/jps/9T1SnuS1w0SrXDvr73pbxUzq+4+4kqZ+oFX1FWuzIHxbFQc69r9JL3MvKlo1i
Vtyt7XNfZgpGsnWdSuCocDL8GxfKkHeu0uUJxcnu+lhbgs8c3rmFlRiyCqSjqCMvqfaeuiFzfLkR
ouU/kPCBkNTJQHLqOLt49FLHHMv/Quzw3J++EFcL3JHL0vjAHxfXtQKUhWWnaYu2mB6C7uIb/iF2
VEpP1OMqmfClMzIi+OYI/t/YaE7+3wrjR8LKz6xKnQSTm/RYaFDY7d3N6t4wHu42Wd4Ars7pjLar
JK5DeT+ygYm19PzUZqNcwIsvsxWYjmv1LOb1/wvAfWJBhswQ2kirZHSDAQPa66SrOrUjgVuYIlEP
/BJ/OwBxIo86Rf/LKeYhv133dPEuKcjuxCEN5my3DA81Ws6y96ymRnpAhX3c9sqdCQxYn0rAoesQ
mrkelxw/bEg4tkPVSxpiw/yt2rHaakMCTepGLy9G1z6c+ywzqpldg4wWnSe5CLzpJOm/oaFBsMNN
StHZclLmnCxtBFqwK/EL4kOTCfS2DlS1b4UueXV+kULTERBBXEHAVd0OXQQjZZKGi3UmXBbPVdMv
Sr8dMyauoUv9A25juUKAH/6HtGN5p1TP0jBMyUXIlI7vzbny3XDgocXDCr0G1EYczwF1TpXj4JRg
mJd7PuHLDw2+NkbeNV/Ubju7GBgQfn/fbditkIWElrouEh7fSldJ+Wgw6oAbzHPThEQpVUsMAMvY
A4wvvN6faWyEycffR61DzPG/R2G68Isk+lFXAc49n0LKQ0sVCkbpiggCHs7lWp5FvNHcmznpclgU
/9Ihm+zUepx9ApR88QV9WY9jpU4GEuCKoD+RdvnRkLtlI0E4ARTDxkozX4O0m2MFUimK9sl1Y9//
IluUBLZ62STI1MfUh8OgvVCChFQgjzYAb2V9iUVKPAeV9pAQ9yvLe6BiESB5SEBBMU4A+kdQ7V4H
tkRTENf3WcXv5m6pe0PfkVCBoO9hsg5Qoww08hgIqF7wY688KvGmfB0FKq6Q1uhIRc4Cw5vHGhgO
/QA7gs8UaNb+ogVNz+nxzkq4wyJhd5c/a5oNh5VXN/GSsVoeHQV/Wia/OpZoraLgKe3mU2QyDqtQ
63wHE+QfbblLF2hw/JAcqRubhiitltMEQl7OkadX5CanpVSEF6XASW51UV8ioKJBTkB8mX7NWkxc
cT8ywL06hVzHNX+r6y5/af+himeeFgqj+cqm74Gm4uOUr/B7va9XBQaM45xE0Xs++yVcnpUI0WnK
jiiD7pex+zztB2VYc3Cmlv08OWn/snErsFL7Gz28tUPGhx81lundfmG9vfJCQQOu8UKdoJexPIbt
x7HRqm4yD2JvxK7k5ujf7gavnnFOwCzqydIGfId5ZA7eBO4ZxHGLlhs8U57AWIrbHiCwWP/tl1RC
GhIBjOzzjp8O3h9mX8FN/Rvs9z777QVHH6mxqi4pU2nX8UUAaGG4sJdZQnnl2KodiIoL2bmXz3rb
u0nztKTk2SnlRUiC7PI0Ej5i8O1WuX5w7uDi+33rxudZnMeYhEwbtlfqv8fVVhiNASw3A1yRwBMr
5wvWklgOxNZn+ZSDOzWE4owNQ0ImOiFPgRcJ/vb+NLI1ZjvWPVZQB//njB+XPcrxWnTFAZRhB/3Z
IudIG9jK78add2CtJQe4iUv8l5wFjzNS4g71Z+nsZgiH9FoNP89oTOuD69dNwLhzJDfDH03R9D//
/ZPqSGtNgn3rdUlfPFbYLYtdgVMB1yYAp5e+t5LoW0sjSCzdsp54KETb930Jnw+iUnNfpGIhxur0
fqm/tz2u50ayMwdSplmlxVhM+I1Z7nadZCbmuAmy7mUiD8B85IhB9Jb+5V17Yh6XWN8sMdXf3GTr
QrHkCVrCylXXWTWJbAttdXk4wkkmMyMvnZjscovdPjRIRmCrxBtm75/Pvd90FwhLGphdqubiVxCT
DXDAaMATrRaPfcx7LhvSk5StGnsPKbUKzPx7WX7tVcIYENyvyqxAeUYBUuF6M+q2/KiTlfwdWziI
P65xFcW4Afm07JWJ2BSbjwNrSgRn6nEgnocZf+i8m5+QE9T1lVtOKdB9M81zHDhk+iFEhjaQqfs6
uVEEpWC8lBH5hul6wWdcPXZHOj7epxCK5WVYjWXCMPSW4w0uOU8pK3YkSMk4k8vzZSMF70eC/Str
ydv6QeqA5H3mTPt5r7/DRbHU0WO7P089pAm5lVMNGT+CKBLJpBHeTQPnS+aGZSpXQkNXwo9w31Ps
Z4euSK6Mf0Amdf1o9wL0EL4+D569RZdsbCVMmDuNgbrYeg6iwGKXeugLrL6sIfRJuQtxQ8xcPb6w
/kawjdbWu2lVtG8Pug7iTETvuFsIO2y6heeHAJ+iI+TECk1WeeCRokD656WyHUSgKHUVJgKMZdum
rQX4OvbKPUfUF2lQrUv5gF2HJR9t1lRcj0fa55P4xkBXFx1RQf0Vb8agbRssI5MHPwTWRRtgfJr2
5cuT80NA2mRQU4X/Auv2uM2Nc0l57mQqdpa4pHWfS7CVWHDDq4erwkPSIG5CozBY/AA3pHqrwJp/
+BsPMIAYDpAJf0kxvMawZ3XhLTHu03mGxTHko6YomZ0kThLlE6t/z2jLL5/aaM83tZ9kL7V7cDBL
HqYlmWr1zRxLcuWbkTvyOv2VCFJ71HndrlNuE6LuUbqJNX81ZEgU6I844oyuoe6ac0bTf+0FVjs6
rsrV66kQHKHMqss5KSvo6I87Lzo6IswuVyZIbGc8aZu0O5wwK2Ylwy+r6XZF3S0ITmDx6PPpsgwa
yl2i5pkdAOfK9AE0qV3IutpEdcbohTsd38VCOwYDhhvopuPqQ1vJd287vJLZuOnR2zI5ip776X50
P5ZJLAlHZh5FS+421u//Q9ciLzZj3LQIQeKRYyjfe+22JzBmY6ZbaQWodS/8L2qJ1mhPQZh4Q+ge
ePmmSIzB7yLj/aqbqlSf80nvrbPkQ6sqg2Ej+UoEG5QpnGO6flIrP96cilrq+sYkgjS4T/v5DltX
wmt3KS6PiEyIZbNOGyfKdEd39BYCa1DLBfOjWZS0o+jqyfmRqCHlqjvylQ2+xsS8UBx33D2MeUky
SbF0CgmlyEYH3CrGX2ADs/kZL9U7l/RuXwS3IaJpUjkXiAx2i264R2t3W/zpSPDgLkxW9r1ZcMpM
kRFwdQFAq+pu4K2rJWgKbLpUCjkudwR84c4fHgp08vyQlwYFR/a8W/lOhT28mmkXK0R5U8eqKcga
UU2GdlNvfS7lvfIOb7VjJWLlv196ou7q7maC+xQlka7/YQqAsyfFLaj68leKpjffjrMjRZhWqJVZ
7JKOb916NB3dHSlTR9J8ZILNf2OK6zd0PYiftQENUnfjpWErWuiZW9iclWBZLA+B5nnW+qybvkVO
ZSmT9Sau/9qojwtvUC8HnIQ9OqyXlfx8rSP2QmTAXPJKo1EQjHTGVuTVkRgLwcp1snFTFNCtPUzp
DJb+lMo3TlIpG8xDRiL8Ml2trxFc/fUeY+qCFd+2CL+HQ0kOIr8NP6ortx7vgW+8x61qbf9l3u7i
RoK6ilxVZPqszMehaPlQRs6MTLutsoW167zld+0mfQIpWqUOx0I4XvYPjiZHTGpS52dFNuheuZui
cXFf+a5zI+iHz818L90ZhaAmAE26ohQdKHTAxiD61S7eIf5SdwOPKxArp+eyebSNN+gtJxukex/F
OSN0OFMUxf0YfbO/bFTYTHyg0lwnShq13IADB2Q+mSF+kXpVTw8nLYUr1NtYwQ84Aa3fykXETOSU
lCVDUWVozH1Ix0riAaByiHVQ/KSoUCCvPP/1iFdA5rdaYpW5phykmuOYVemELj62Wk1QtojFHZqB
mR7NF6Ulx1NteR4TsIdHxMFZPKjpTi5UIzP9V8S7k8bN3/VqA9h+oa8d39mvK41eHrmphinPmAJQ
HqDO4olNC/sTUc0TGrfLLAUDHNC3YdCWyb5rbNcKZieTdPttW3SXwC3qFU/4xeiNYmZxYXsKX2Dj
3Oirj4tNxLmXlYPGnB9SCOB31XngXyrJRuMXxx+3DpzkOKfQBJEcQ0WMEUekhR1lgf11TmtI/V3F
rIPqWe7CzBj97rFsfFGO++JA6vjI4Rt4CEIprGTVQkF0xfjDGJtNtvj7+eYRM6TW7recvAqAzMPw
aN9GuM8cawONyQwbgIvdU60pfzPXJagEU/XUyhbP3bd+6+bDiBvlRp71sllZT2CjebRyF4sCI2MM
e1uKZQrODvA13nO9d+KvppoWu14RN03EsR/fmxgxtir4gSMUi7JWSpDX1c0zcMiqyMtwXBycTP8Z
zSevViV7WdoMrHiD8S7y4g1G5IHU10HjFOjzVrOWQrIUEE3iFIDO7ZCst3xROfaPbolR0U8Chjnd
MrYrrCJsWNVDCTprppjRDHpng/Bpi9pnI8J13VzUAq+rZ47o2mgSTPsJm0qo6NqO0oAbZQIShG3l
SLE26xiJK7oITkjsASllkTiEHMZeR2ajcomoWjSUCok5aOZ6Pyhk2+hdudV+x3wIa/hk6WWG0oez
w33M+U9+lqCovqs0oqsi1w0Z5c/0Jw7l+s8F3qjwtK/COQbhKiBo7uuE+BZKeCpTKPoSh56eViJE
6qW3uNNDkvDk1uRf46xinwz7YAGrcm+nXuA6EQ+r/VCmhDvEg5JUWHQVnhwjeA/2JlvnuWIOECBj
SWJfTg0D/IAoIUwZG/6yo1xjGUAIEmenyz9lROfTSa8kpDFRyQM9eNZWI02Mynf0rSwHoppEiuSF
QTbIeXNntYYhdUy8HrklzZeqx6Od999W5A5xcg1wMj2p3ZUwx7vnBAQAhcougUXRoMsXVkbUgTUj
M7Uh1vN8xHcpJ8KnrwicwL2L980D+wx2M1EKQu7EqIkZPqU7VVLajhAUIfDxCJQToGmT+kucv6XH
04diD6JvIWxWiDBr39Kspu17s3I+IeyaAb09k8mRkk6kvBCl7VcSt9mRA+d5gl5sO+qxsMgeGMY6
1ovYrtm32S7W96dBvHWEb/KH96veZA50Esx1QXcHW4JQ2Yupt6rl6HlXIuQS0wjEVu/Vm7jsHqHM
/+d+wXuTqCjR8B87tlggeh9U82ous/DHvXvy+nxcx62xgcUumHFF/YMbSO5J5rafide3a/J+UCbI
HAqqtHWaNIPJl05xh53LR92jmEUmUxL9OjMjtgYagOPeFfZXTb69zSVs9/Zejj1TwTU/7uI0OBdA
aZAEAObefVJBDhxd9rsqNjoyCRcNDevqj87kmixBH/pVgx/jT8IyGiPee3n/G0P9n/xEKtWYSHqW
ZB6mv78hoJ5lYH4wsHZ332QgWMVLcAOwQNJMveGrp278L2VUG/yMiOg+4KvnI6E5gwhKO+RNdf5e
6kmdbGdjWJqZD/iYx602Pl/N0JJE5El2u7YlNfnDDqcCotywCrUzdkjoH/Z3eHsV0pnVmrvve1vP
Y+dSeS5qOXMJ6Zq3YG1pcnZPRSqGoaD7/EiFv+165uyJsza2nSfcAEeoHHF7V9axcIdR1xY4ZvMw
rZKcuTUa5uwsHYPHAth8arA23ToeRIq6kqXW0u0Bakx7FhhzdHX7mnPxioXrTRv7xy99bu6xIWfc
vjN7ORbk/mzn4nsiSX0w6f5YqlP9SkR2yXebQ9SFs1+WYLKSFCgb7MtrHs4x5uvK5AO2nmo2Calb
2eHC4OTQiukynsV0lDKJKcjOM+QfzzPjENygl9+W/qTvd7NfZ7b00OxCb1pBMLcfJwRtsdHXfL8I
JQt97KULQ1Ug9lBAjn/8/WLglhTMXpEKXJjBBAbm6nRInCKEuHYJSdTwapJHUJnojYetCrjizov1
b8M/MAWqtRPG9SuQZn9OZumMHFoE9B/JLf0kpOk+8EoMBemVOxO1zpxydPKBhRFspAw93UjFPv4Y
twOfZ2/i58TMQvqlteNLv2DvHz6+Yn4LUbtpW2roBWXDdOTSfK9F9bARWN3N2U3GBS4TUgW0EMyF
xpjv/VOTsQyG2Dfgqen4VZ4g4pg6YvHXzZGEE2B8HSCGOHpTi5x8CItGxKwH33B3J+muhlABvteN
8y2r8XqiStCJeVf0gBHlb/0p8wJksxr/bbU1Zl4xkiBszd3BLBg78blUqzgrI7ZUvi/v15Jl3hNP
wbz5J8btv+0ja9XrtcJChUE65pJ48xUwVzYkx19FC1jk4EXuPiEvCsp2QsLEA5SR4ke3ABUhrcs8
4vr0mhvScrCzxqSFCTvkGMFnE52vV8HiRXt/gBkI8YUu2NEpHRjUE9QILk50h55fwU1RxwpCRnH+
1IOZwGe0p+yrtRrVwaISjMln9SKyZiFChiy5pyMc96/gZyI4eZFnp3LKlMOOaTPaZCWqdCptDesJ
7Yf4dFhneNJillRWzpDvfNcihqCF3kgAOTjfHwOtnTh64aQiSYSL3DHJT8OkAoJFZokqgIog+D7T
hyTnbng0CVjeXvDMLRnGkKpYJdLpNQidrkQFL+jyKtb8AyGgh7i73p6BY5/G5+jQVlUYfwSJcIC8
rxug1T7ugyrBUN0B5i2Qi/cmoIFdQ2UA6pjwLglLR+c/sf3eVXWTphFEn3gGsIpJ+8oIQwRZElpq
RJEstwjxPrPCASVjsJsZyEpK3wQJt8RFz2eRIMqmmSTOVd8cjILoQR/9PwfigRotkp9OhaNaTSwP
sxx4NGbGgtb3vqZkO3E3ufDSMC+MUL73R1ZtMwS0FBvmKqmvQb/OiSNjgPjZknrJQB3WJGW36Wr9
px+FS6cdiryzzTNckmcE/o4tBSGSDDpSNNbr7fnRJrtUQ8ScHeoq+L/+Tc8ywgNkU3f4QGgw3OpF
mq4zlZYiTkTVETxbLBOUhmof4QjpgG6KnCh8JN0VhW/gjOlaH4VGF5mPEJZ+M+5FB7hVGK00FRPo
3CKR//g8Kha365Zw71bnbryip93dvIEpw8e/qbU8seDcoc7DS0e2StAk8j3GKflOd8cNuTsGxjbG
MQlqkygm8YIuTvGwBqxX0peE2oKCJwYJa5gCjI2FjnJCVUF1VSY+TytW8sWFaRPPXyOUXSmuV8Tk
kr8TenB0DWNp29SeKt3nGmMCPLrhOuqh++bPRPfmOrnm8q0guDcVjAPFS6JslXEUOfVwBENj7i7D
s0Smr5z2YIrDtkSbGuzS4toV85PhpLctYmvJJwNS8qKUrIS6pNe3EMp5N3YLO9CK9IW9KyikVFIi
QG8z8ktIgC1HQsq51p8sgCFwIXQ/0JjZyz+blwOk4z7rDCMZPjOFqh5EBBniim0S5iIIajC480Vg
Au5R7UQxFKxkRZ7wra7tYkmqZTtDK255T+bmuN7gr2M/UsswFqEDEwQTjHSBZlh+JQZOwBkcTBWp
zRIYTAIkb95EWhGZ3ZcDecJBtmuUQuFhoTcGTDQCabc01exmFDxa7yhcGItTal8CUxnaYB12hsfC
cAzlrRzys5GbL1JIDSEU7TLCa/agpg1t2GlDGqk0JrFOMZWvUonypxsPfJdws2+PJPO9sjEbew4F
4t101agQGTbY6EkgPIrd5mloTQL4+APDEXGYQg/iYYDdUgjEvlXqkhC9nGhor31t/XGbY6vxsICJ
4aV6CUVvEMlOcRkp+WCy3IeVvWY5wiVTMGQ8pArJN1cDHVLiaPfZzlV2b7HVcSUMBHxIzxewqoHY
ui9xbGkSg1Y8q4sApDBxdyXiUYbJZ72jYOUOosdW9mkznJQ5ENcT8KSbb9kNdVxETXjjDJ3L+P0i
62/9+Opdjhd3syb5Tl5jTeauixN8qkBHSqYV+l/ypJe1ByM5/iwUpPWwq5KHyRUsu3U7wbUghH70
ytu7izpY5Nj2Jid9ybNa8HK3GqL4hzrZvbiAAyIpBp8SFU3CRwqUzqtkNgG/5TG1RSR+4lAHBQe8
rvBvU2ASv8YlCJQb/kHZuwhrYxiZoakS6PsnT3WlFAATOy6SxSQrNjyKqHxRf25jTgboavh1zLUx
NAGmJqFuY08NiwPe/BDFI7Z6ZPjvpaD2Kz7G0lqGvGT/DOWGawJL+FCY/6I6+LqaH+q/KM4wzMcn
aTi7RnddUWwqIiCSs4g0zIHEyHTHj3cTJ7RwLGKoMGS1YIC922jAg2SYS0IyD6zI79B6MDWdTxxy
Ts14zALhGQbXOclbrhCNLH5cTVSdDWpw80KRC5Rxnxlcf0h6vjb28QbnCEPGMEj7E3ITz9Dkodpe
mo36c6HBqpkQyECTs0PUM3nGU5wS7kWmokCO34WlecwNEKGP1Cj0tar+rvW5XxmywdUVwi2X38WM
cFe7JgVFaOmLw+SxY2O2EynMpC2NOKQTloeO8sQURMGvu4Xbm05rtc4/5Wqi42HtwSH9z5Y77yjW
BB4scduFZIUZfq+LVEy0WpoyHqkGEvKzUNC0bwxKD1OGmrdx3zeuxgUyblesgrORsq0VPAZaDu+T
aHpIHvkJ9cMxS8CGB3vroW30cKs9YlPmE5SiT8XBezLzZHFyqYghCw1hljvG6kTupAiNdNL4Lqjq
QO9C4pqTh1k5afkKIPy4DCdSVy7OMFRWX8a3glzcO30/bcnGsQDzMpu5dqOrmcmL6w3Z0XRBzlUi
EsLmNn9h6V8nwRwf4rRuZK9DPXfihJrpy/XYfTisAAxQLgl2Jz2S7+MCW5uUQ6F7WlFdN+1x5KsA
pyl6saMyGSB+oUp9uG++g5+H53RHZIH7YqNxDlZ00e2TVxGc6KTqqrDW42OknznBUmQBVj44vmxT
CRDoY0tI81KRlxCwfDuBxBszSZMKuQcP93f8bYk0NQF2gldxSgcxn3rmJKRm+/PbkxvBcGIwMeH6
4azgkWeBxV6ygEBpeEtM2TxBCiSnOOHqLj1mPDDpsfWN61GWKBs0eNDixlbGt2F4OS9bpKBt98fw
CDvXF2yDnOTRN2EYOsB2oj/CbC1Y7Pf7FgQ+s13V2RGeZFCBu9TOzgAcRiTROtzmQ89IcSZ62EGK
LnWev7eJCLaQcbyu/tJCTCC/J/rN3Fh9M5vYhLtZLxr8A09LTmbonOhUvXhiy6DLK0wYnqhlAGkf
+tO+KU1+AGbm1/pYD22KZdOi97z5VO8adJjCffstfYEWeoYgde8pr/5H5MFhd+J0r0y94wsOwewe
AX9wiCKsOG2MofYVYBtEEzseuFgK+FhcejEam2bWdVRX23NSrHxL6o3MoaWzSmUICmRtoKZ2Hxdq
G8CB0QM4H5J3s52JxohzFAA4wNmRRzFNwC7hTUk4cKJRF4TO8g6atvPFv3mkCw1AsXD7g65r53vL
s10NgsmS/3AM0d9LAxed1fT/9d7eisAlfWa2lczj4rGHbJgCEP5AbceyNmqXAKgEwS5Gq8yto9qt
ywD8zc+Fqwns0GW7SCBavRIhGjS4dg6h2G45hfS/31k7BqBqy8p/VwacI87/yn8HldOUIKgubl1X
XqxaYXVqccJH51dWPiOVBA4q5LtwOfbv3rYaInkQMlxWFJihePGNr6lCxjnm12HW9sgLziaiDIEH
eeOQQPva8fj+dtLvyl7vaEa2O2iLsK4fIvOyjmld7/X37eWW6j7zQ7DQ8cOnE6yra7WOAvSe88Qr
vbVE9faWwW92p4decTadgqT17xxwOuQATtT0gwRMZNksOgdmNVsVACpR1xYEEZO7kEZH8ijME2x5
ESIZvBONomzbBBQ36+CjNh8CssXc0zvOeJcjlNaq1Y+btvRUuchRp0v5lQMB7KsIIS2PvYBNpFqM
MRewuDNyQZ3HtkejWR70kBrM/0q+XPHidPDD9EYe+nlouuLst4nGArbkdv/gWWjbVBiJX7rvEj21
Y5OHFT7FhksT2TNgZaJkSESu3K8d0GOvLZjnkLGwTjittcGOcxoeQaDx9+zoK5mZ3IjCkBPAWb60
PuKowPJXURtTX+F0TtGdy56Hfzxko1Xuo3Jmc3uIbmWdEme96kIjNGc0Vy6Vni2w8SKmKl+/grpD
rf7yqT5TiKn0fy9Z8iEBTtzfoTWR2M2clUi8vYVLhmkDORRgHExZHyYBsr0NxIut7garhtmTes9C
/PNGSLsgMbBEHSeFn40h9QJSToAYk8zF4gob4N18NXV7A/6fnwlOEb3+VmbrGAjb9Lay4pFuIbd3
ueYJ6w90gL8mo7K9gZ5Lf4di3NpJEPBuxb9TUyuvHfkC4ewNdZYLbg7jJYxVRp73llQW3dFEKt/I
P/R/2qT05xFU9WrMm3vF2UXGwAawJDkQ/0VsYwIkL+YK6+kS+D1idntAW/UoXQnFSvZCUYAJC2Qz
Wg/f8UwsXm2HTl56W56GCIiLtLBYqngTeYvHERjkvBpq4VTSyBHHUuJtIhpWuOTNHqrDorOn2lpO
NRRYOi/IEM3YVD9ym/B44WjJmc1lAMLVWvvOZwnAnaxHtkK00eg8VhaQsrlPjBkczUYi6Uo+Q3MT
yF8jjhx/QBJ9uzE14EdmKsEDFkoa8h/ZzuYC0AWDSQh1qWD7kHtrqdPsuOqBSqr1tF6yhKu1gX4J
MPmLNNKN4s9datA1Ga6StYJ3DRAz4Qm0IDeE5+M0PcYzmr0Cx+XQyw/6FUk4IzCsYUIx5eX3K0n9
teq76sFjpx35LWV1jVgAKuOFRqpwL694zf916ZBJMOGlOs2q29fg1ETIcuAJDeRYhedTNA7mgJzw
5Q9arX7iM1pOT2rQVLt9kqzlcODyiW/WpGpCPx51+Y6VWdxfwrJlJlZLishfAS0diilgxjrSr5fG
NUCJg51hpuDgGvtgmoHh+kniPGEohmeu/fKADwVmK32maAKZIZPqwtV/yP5F78Oz0FY+jcYCfNqt
1AQD/JaBywzloY616B/eMmjm11NVM9ukI/QdwP2Spf/55sdt3rxhJNoUVG7g/QdYxER1H8DhKDCy
hJ6x2cPl9Q9S1cjzz61+peeVpFyrWSit/RkLxjfADI8ZInHVMZFThteOHs6hDzNPF6PNg/1MUTYc
+UQn0Z8mR6Db46+PzThv6oVfFE+9WZDk8+TYAkkufJNqWQ9whOmxrd7QG+yNAT0n4jHKfYEUqRi4
yV48gBO9zA1G/TgSXy0yfp742Jv4nIj5ityd3v9CLxeyc5XF48EGkoOyAS1vk88VXi3WDMSOGtd8
2NQbMA+oQbQNczl2f+IW8ivuiYJnkj2d1o5ghvs8bs+mYPoQqktK7IBnABy0bdrZ1FVUGcdarX3A
Wx5KHUye1raot3JAgSXLAiE6y7lYKVgh0bJi08iaCtKI/VCaGrVKjoV1uGaZYKBbLIH+IcT4PUII
XU/kspLvESZyxI8uHfpi/J8O70RRmXjItZp/yA3yCqdRHrURZqzzoGcFYdH2M741JiARJLsrCywY
AdFlLcYFgftxVD5Yp45d9XgS79lV/qhKmCyTctvgZbJ1CNO90lSkmy/QxQIPwWXFuT2wsNOzcFCC
JNl5tq6AbshKlxQtjwNOuLaSBWl43o61gj4XJ2iWKJKOjm9h4jINFcjkUSoLqv0HoTu4Seam6mLL
KohlgHF/+oUhDg7jj8M+x6/HTQly00amLcx7czspW5pR2IBnEDc5co59S6lXkGiXM3OigPUfe7Z1
GAJOYBp+eEnnmJfCFeAWcXylgyobp/gJfASnNtJyhCeg+DQDGpR9DxR6vr0aeibV+5FNFx2NCTxl
ynZsQ1Ll3RWIXTUIwLQPAO6vXWMAvKiUp9GxYXR+20GT4hqBKWY/G0JUHdHl+q++UWjOr3h5Vo3o
qy/LgkwHQU2NO4hFhtB2tV+C4llGCd0+IfoJ+yqD0PbZmcx7Jrmu8A0sQeDb1HEdRA0FvrLscr0z
Clso4br6dU3u0GihvdqDmaSx0mkyKTjG3hrfsu6F3HGDpevYC2WF2OUimetGaZXgHZXxkKdm8jJm
2aKyvit0R5eigKK6MgA8Xz4eNlZwHO1MnqeMf8dgWhIwuzFYCphElr0LE4OUObF14jl7MsaIdMzN
3CitghHNfTqstRRJ3PQrqajqkcSjBq/R+MGzlEBNokr1CUDjQeCIk0cxFw9XeBT7I+JT/tLZ1xeF
Rvrg7D033/guN8M0pU8W/WYD6w6Sq7X+b7N9GtyWbgz7bCPEY19Jdk7aHDyH7ipFX1bQc5N2q6c8
p0GUDzr8FGa7s825nnjHk2ynMYPlf2+S/R/Bp38Hye0Yqlq0Tw/eWDAyVvDEf2v73x9o48J31kO7
vqnrnn9inz9urm1cFaP+T9/FGrRSnVeGCDPu+/hhl+khpVxnljbkB3UmwStVOlDeL29E482DGqkE
nY1eqVHzBtkDaDX90M7YGwEbj0X6Hr6PRDO/f3+3uAtcWH210DfgPhmyFNkwbhErwMqAmTpcSacG
UDqVZkc6gBl8TYfv1WyCk5Bcm87oy8rTAgqVjsnwXLCxA2xZJPdW7oUd5aipRba0qRX3q/TK+lAQ
QHDSt53VtRo1tBn2J1tCGHUKKKRFOiuWs94FP6ND7NnlmJB0cRs32VhGD84HyMWW8zxe38hzBdRg
EBxtefF8RbmqIz+7682GBhQCqrE7EyIm8JPvwPa7DCoxXgYyWX+Wc5qnKBFBqeZuTPHD8wEvstye
hjZZaKNxRdE56wSY6OV9QZ1CgXdCQQbd0C+PzpuaWCtb9AjypsLqUsGfWqWzlXJ2/TpsAPxurkQW
mFqRI9+HN1whsK/YTsfqgAHxo+CT2l2wnqjVCXFx3xjRiuhb6PoDaPbgIzm0XGfy0cnrARPY4gPW
7wiN1IVec3VAh/5OWe2evgvjLp1cS+X2JwKJgmFtKjN/xvxSZ/fEWScja7ndtPtbUXk2aEb1Qna4
vPkg2xkjd/CI9iqayZGqjVH+bavU4jcqXlYCEUWJ3zWTOLqn65YUaTaNxOsr1vpVvio3U5Z4zMCk
l6YOX4MCtjhPFn/oEx/RKJXkFhalrJOcpe5qeb53B5++0HsXgPotzdzF+5uceoPXce0vqSTDPTW3
vAAFzKC4EftoiWzE0aVk4zbZ2OyxRHedEGnV8+iT0X8HDeuCdo3S/3Vg7pnOoWE1dPBCQbnvTAmd
C8048t+JN9leXdL8oYqZP6hsd1GPYJbiqbq8u5ZdZxiuf49OF/bUQ/UjxTWKYbnIcRMI1hta3/MA
bC/yPt9RaXgdG4C5v9Y7Omc/2tn+4FpHk2hevAgcfsXkp4zKawOL1rJxv90k2lRbTkIMEzW+za+b
gQ+JDwHgWjrGUB5zejq4cX5McxE52741oZ8GoPlOH30zrS/thA3SIVVBGcNIAqHl951n03rm5eLU
0fqwC2WBhqGjxlatnJztyOOzO6UvDUVlrWEXBkGx8FrQ5b3mRzWjwieH42yHnIL+qT4MJqso9DUA
zvTJjHuXTD/LKS4NQD5NXkGQQHKiUFFBg3Qn9H5jpKmKV1hav7lO0BYENYdScteu3tZPpN56E17u
yKuUP+wLTKmU/A2K9B0A+BCZPtuIq67T3gjAGHSm4k2pLMnkDytQG5i/meNLODO7KRQRy5sKDL49
Xg+EyzcmwKuI3vyoL9WVywR/XdUFyg7oZB2dW96sb94kj80cbCXam0Z3clG76vHyGd6MBZQACcYx
R3TETVgeSt0vZNQ1+XZRiSf2dcl7pPTaU4R0SZdFGYZQdPOofmueE4SXoJnh8vRN3+5G4E2HLWs/
1jAxQzj++RJvgC3vhCGkVWiiB5MVk746S7wMTMWLgc5UeTX15zN3r5zx75wxnseLcW2iaewm490/
Q7DXnAeTt1Btksm10E8hamGkCuwYPzERQCXNJyaee+eqNaTNyxX3uuvSTjdjyyCGfi5pLujbodVH
S72KGBpCyHZO+BdaCYbQ2lQ/wmx/v54Z/39hA+x4wZkEPz8Z9Z00KZh5w2ZamOewtfWpH6ZxSRPp
9tJHAk4F9w90pP0EOHzGe0n7zWiTQJr2pLnJb2FRqXIoTFcfuBrzixNA3UuvzLRLZZgiaj0Vs9kk
uMpyf25OBKVplkLQLLpbY94cSs1C89AMdeaQ5sGwf3uzENF8Xks1EWj6SyfDjAkWaKFhNjMO1sgS
kd+cfDkskCaq9v5pM7rge4vJc7ZaC9EKqwGUmvL09+ZRe5MZ/U0d3aG3vaIZWtG6E9DAZfn+BHwo
xHwzPag06pHPSlxyXQCISY63shBB7c2waqn8+hWjLRQppTZ79elYLY//9yNYwr11EZMoXRSWkcr7
6hUoutNYI4IBoNdiOUrV1yoDCvEx+j8r64lNokydzPJ9aP6kaZ+dzUjdTnTfGJ3yTKMSI+92SV49
KtELbOHh3NatswMKKv+h5BukS55IIwEnHmUWfxTYwVxoBa27VpkbaD6mO4h3UnYs1xaFiOkZbj/1
Do+Kln5EwIuhxF78ieCa5J4RDacRpdGG6Nn0yyQmldG50NBWPf3ZtjJyMsUqrE21pwUdJ62LpiIw
3E7qrXsAR1JJ4iXAzUrrIUC5diUYdntZtWWa6zmmTgJw0tTFZigpjTSBte5hi3jaxzr3sNgTBKnU
udp0iMCT6m07pdvRkrxnLeUyxVD7Psj461zdIFkWcmDr9ZMDhJC88pzaCAwbcNzEbVyCFvcpyR7h
XVzsoIF+wsMXBicJ7lhdjGirS3nskSja589VxEgUxlQNddFOcLMrkTR5a2zhOLC9KlMszw1beCAW
I2xaW7nPh0pUno+FJNu8yjkmFZnHSlFf1MA5TWnPyR6P6EdcAnWDE/u2HdG6jM5JSOM93TITsP6h
hXHpm2aYOgw6eohWecfu+etPFy/rI6TF5O/KsIyQ/qqqWLC6JATwPmZ6vo7SsRpoKPm/Xa/+2ADA
vYsU7VN4/CtspR2TgZ8NNV6KyK2c6lPMcBCbpn9WQquejpfEsgfSXVSmMaaHanEjVWiLFlZhCFfL
aDRyb+dJGUMKgBZRUTqJOniA3mLWI+S4vn+Ah33dyXVpk6klNdqqbXodAFfIgRwWRJt7A+Rf0c7y
Nt4gDnUpF8H48b5mhEkkN2RoQziGWVouZnfrbadUR/yEpvhvL+4mtAEfDLud+rIKtyNUv3cTFQHZ
P2vbYK9FxWYuHxyfIqv+NlP/NZ16UtfSFXmqGiL/BhG2ewxRmfNJU2HWssiD9pS6QTV3k6GdoP22
kOavOvEx2wKUL0K2+OrSd37j6p9ObJGhn3XL6DKXlO9NYqt4u2uiZzGFyK5EvnCNlidv0XahZaxj
MobwYLOwl6b9q9PtdH/vub6I67NxJOLjy/Tdn3UHlH3D7uWPgRoI2tMTttdbA8WYzuTZ3NvFVOOs
FmwI34ewSGK1EMXi7+Mf116fF4Vb1ZRN4kqcbxT6X2gv2tBw0/wsNsXtuSdvc3SOF0xTqAAuDiFh
pucEpPAdZoI7KrifYyMCIkniLioy4yiCO8a1+dvLS65XJyVcD8u2r2leHC1aMS2JAjFgIoRAMInU
Xye8yCa7eO+HDV+6hOixfFkRXpklAbGDcINntjVJc5fomTSy3904jFz9M8L5Bs5gLxWxlXcgO2Su
tFpuJ+afSaqrWBXHyTTPDsqedzqP7zqP0dtiPBnTVSozURdmksvRVUxbxLgT004aQEBhqm/p/z4/
vapNnNv69iRq23+x9JQFHhq62BIwmfi2uztdjbO8ptE13p58VZsEnjHZNatmEYWrZgZU5V6MhWXP
4S+upZbvdCffMJSEI1W4ozlc9PzyUdqjsOWQCRd2neHd8bASEW8ep1v8hUCw/GgroVRmBL2iRCxe
ei9Z14fzUGevtTzPlbAqRJsoNER+iwF3KAItlkNz9JIWn2fk9Ts19Vu/TmxnAClLLHauZxcrjir6
avEEBSTMvsMgZlFdvnvDhI9xNQcpoHZst4exFPXc20lXL2t4b6UxM1C5+JRL8t+jOVOpzWEivLWf
W9yhuYbI1Sw8G5xrMddM5mwGuFl5QwezT7D8FFqSmgc9dW2OHUZfSH2+Gs8U0DENj7cjYHo1YVMp
2MAVpWWKgraeBW6ZY1l3lpwyY/HALMHT37kzOqU+qLku/+pI/LHXMbFkmFfl4yyIktnGsdZb7qSH
DzwipZ2bipA/glYnky+7/ntwoABgVWnHeRg1zsIcnWkEPluagaV+aZzCh5+JxtPBVNfB630vaC4w
ll9s1KvrGoltsyy5mwUq0CAv/GcIs1g3MjfHhFZgvTQAzOyZoQlJn50NIiPwEL1wlBR8pw2Pm9qn
704kuq5KyWiZ0bAqjdyWycL8fu4KHxEFn7K1NsQFcCQ6dF2s3eoM7Xr4LOChuStn70GKaDRDWFBy
RPAmrcl6bIowCKviUxbPlIK1szaVbZ1HfplkIvZRFXs0TVYBzBQXom1bs4tw7JHh+X+YroYZADFm
tQL4w4nKXs1W1zY3PmrI2nKwalzd+usfLHiDFLaxWrFsaddqhkUQuCJaadxTYubSfSMeDiMPXbyq
2xw9a7ophyg4jpWh9L8C2abs7DoTJ1yDbY2Gg9Asgtwi5jPPVsGUpfymCoHcy3y/nEW/cxrfiR6N
N5xLRKa9hBmGxTO0NHa15C0qzEOQOoDQZodpOlrR7lTb9G9kiFuSJ6VJjNRW59rZFLrTwQh1Cwk0
KytZsK2eqnXa91oqqWs9v0ATgxvvA4oIU9DFXqAQ/FMI1eAKIvQ9YtfvKc39Bnv5Ed3CxiKjj8pf
2/q3rtQxIRz3XLXgihyRkhIUHs5nz+gmuajc2Gm1Nt/FbdKwt+4FJEAN+3TFvoVF1n/pnW4/2Y1k
wQYePE4aR/psX4tI/xZ9Whpgo4thRKe9GAp2g0aPMRuoav82piRc5Rg840XruL/Eib2zfhxrmyBi
babKrf2gLt4to1n9OagKBkF03byu2OC2cn8yobC6b9JNhHaHrk79rpjjCh4Og/THhiP7RrSGDzDD
xr/jbCPrmhNDP6j0/M50FJkyYANHX3yo04DJ8elz834EB5pt9kfbO4gSis2jmb0H3bia4No9+kD7
PKr52UGrKaAErs8nwtPgjpat0T0yQiGcRsG7/yNhJzKAu+ipY5kOuXLn7Gqeh+jWSxqlQ0s5oBRg
6QjUSzAQmdkvJw+gJJXSG68Fr9fcFL+hrD+bA+9Zmd6h7FIHvOI7tEIoz+Z35rbWOFJW3Clldyom
UDzTQo5xxX3PcoYAWv1Ma7YPXVDV7rnyGRVtm26C4TOZHkqe2WSeAHiQ3rO2QlAc1lEnHdwuM4MO
Fc6yJtQAAwZ/Oh/IfXrjjFQ8KReUHfQ7GU6sBjfsY1e84y6QmUAw9o6os6qg7zdx2T+6U4Lw1uws
q8rsa+9JdFnSJDbOh9Vm/oVokimKkKe75Oodd9KGX8Olyb52VPm+5u57rnfNWQ09qt8uUA8ykJoL
4Kmc0zeQWuvEIfAvIXkb9EFnCCbMYMkq1Dmz4RHNlVGThbsdmdN4O/4GMrPOtAqc2Ww8bPNxaB2v
vQ07wjb+JxcenQ/N4ETLYWVHKdWXtS3AJhr3Qfy96itW/p/vYpesZo1DU2KZ5RXQbMynSSiNq3P2
NyQEZpwWm085oIWYxsZDLYRucgeFZS7+qSVa7whrW8WWQKZHM/rzStqoZCzS1i3fh3Z+XRPKihVR
cxXhjJqlx8UtemoD0cbyloXw0VPhHyDd204OaunAM9Tv4ZiGyBwhHVsOWQSTHif4IOeOgrEfzi9M
/YHTCChnIbOevRy7mnVmd4lOmBGOVtijpis96oIHdlaNB7oznQFDk7SxifmXgO5VBsEmmgnZX8GH
Ti1rfZu0xXGVVqOcpRFV9l4/+Q5VQZEbgJM208AcSKhGs9bfneePTJ06t6g2mnrM/Pefc/R/YPOJ
ditdRh8ydAyFei4n8AZOEkn6hXj7F80DKFHVLmbMWtKwBOzs6Z+sZFJDveo0Mga1mtk+SzRQmsey
IsDyhfXawRP4zJTYhGaOCxbs94QMx2LuoWMJIDaYx6xEdf34XHvkp3joXVqYOnU+FOEd6eXYx2qU
eXUS51fOh3YrEdJbwfsrNxj/K0VgocGlGbUvG9LN4nCAekqHNa+WnsfTGJlMVDKb56xnwhmKpXw1
NCDOuK70mo//BrwqMieT0WBVkLH9GZfXkpo/eWCvWTKwc2uv37Ok0w0I65tY+deMrArqToUynJgD
ywDatQJFkhB7Uw5tGenhoaNdE6mqHOX70jYz3vfE/oDFxybz3nG+tuzaGDidFIN0tkzdlc7Hh14F
2crusKTt3TybkkAfag8dA9uCSxTm50rrj3LKR8tzcXEkyR4Wvob4fU03AmsEwSN8E6F+qT/tJjPT
tiq+U46KMigkxvOTRKmnO+3V44aHs4rk6H+5uH/jSnmu+yoVPNy0kLknLKpUchY1K87uENHggcny
Xf4uvSz9GD8vfPMKOracOeTUzdTsIFYOtmWUS62tJSVYbWuoxOb/BsuptJu+TtG1Ff62WNxQdrAh
oN/bPEHxN8uf2hNBdQiMoMdK/8rvrp7t7xhAiyKrehAob5YOv0IoVMkmnAH5MJyO9E7OvgPh5l5B
RjUhwafduVKJjShn9f1nXpQ7hgfvhaGlTr3WmZW8TfsJfcAqotDN8WvEOagJJe3ZuVvJvndf968Q
vxEQ1x2c9Jb2qHtm7CRSSKhAqInoH7pOmFvqlDhwWJ0zRqYFUtQ/a22EYZUqUHSUvIjD925y3ogu
QnvMTcFI6VCRlYebPa/DgUXXJfu8uW5tknqwkVKK4UILKfsRK7hFCCKsk6sXmoulU4cKKxFDueOF
jDjN0Ktz1xml2Lx4D3QkUThiywafJLnPHrNiDnKSAM4MOdS/bDumQEHbScMpvXvvTqEUmSXy40bd
kfeUUdRJPz9d0ngMWE7P+JPCkj7I6Eu8QSIfpY0WdHLCmA1EljihCYzfGryhl9rGjI2bK63pu4Gy
r1a2Wo8fKOU8JB7HFamHcCcLMFTnBoNS/eFclcTlghaG3aQcvJiftMH3yc08rebApigzKsmWtk3V
evkYnb/asn2NfD6d/Saa5FY57pFRFv1R5Rwyujh5jRwiSA4xlInWmKRZQnjLR/NbEqv0bA5Cx8O0
8/WKoUR3tuvdVtLGopaptOWN5xjR9/Vgyx2FB665dQXm5mC0y1UAnTTiQGCk3j9EvaRfZ8mkrcEE
IlHZuavKROWDk/M+goyfAuDIgI1VSvEosdybjn2DKxLm9FSXoxCLm6FgrnSLW6/bjVOAIh6/tGEX
gkkdftWLBr0y8xa8urbYk5qWzBbG+G1xjoI4KMsxtHN8jZZL8+7WFkgT6PDRngQ6GRnVke3p1B18
k/71jScShuOCJl6yiJs5Y8dXI/FF7nMSR8m741faV9t7CoBGuwihuqNRdYhl4quy/5WzGcLDJlqD
nqVc2jsBarE0FWKBMRXDv5Z4yfnqrk7Tc05NDSZPs82d3sEcKWK39fPiZ/zKbb0StbzaC3vzdq6p
Pl6YontBv2DShdI7S6Ty44q8vrfJuLB+s5cbI3xfOR42Mqm9e4K9JOd9VTmiDjiXXgQ26qS/XchN
RjHqQRR4KB4MUbz1GyzwjDCWKMYcEiJbPkHn7ZTWIn7I6n4lPafduhB9caC5fGMFxR3uceJBetTL
5si6e422yLXe+3Aobfm6EQ6YOZzuGYfm4q+HKoNdqNtsZWou0athm+FmRXIYTLZcY38dbrOOsyBh
8zo8Hb6GvNFQpLspFBfHN7K/jJ1OqewnjSCnCnjRsNJZzIla7OMzC+eNU0TkW1xGPNzmB/Ypyk5J
F3l0g+ZyxiXrrcssis6HBxW6Qn/AP8VAa6R5OCkJbTRrqNGi5VsR/dQrSJZKcE2V/uNJVEib6MXN
fkzGW78ZiDILOxHangGFC+Bn3OatSOr8b9Y0texfOdJ5cxNXb1XXKx0Ya8Vd8DSPn1HeEez+NJfc
iOHGN6kg/dMmqk/nAy0Nkj8rbGBXmbj72Au6Q7VjSjYwCHvK/ERx4qics/d307TchHJJ4sDmZIxh
8ivdW5tsAtkM7f9iBn59hPraG6qGFoZ27GtOPs99GtYUQ79lGoge+XKLMiJ4uFNxZZtzOnrlXI+h
S/+KTHpFWwBV+eL7KzV3THu5RT6hiTTolROU/mOOrHI2RmnX5PKlxcMRWcLMrRB5ypxs7kzjiTmW
zOZM3ZqQpwXwmf5ExIM2AWgGAzRqzDxL2qWGGpk0EcEnzPUZbAcK81GyWVGPD8iH63YyOrgybOd+
NKiIHUyrcCLPQA2HC58ItXiEOEUY97Y6cXd1GG215Tbgpt6fTNgLtTXgL3GJ7jG9RaMXayAaCjGV
idpoDBvgS3fAGgmmIkJDx2601vPg3kyC+EJN00MER47/c3DczTjRHmqn2n1MmEwuDBfYxP6AJnxX
nme+t6GsLUzu3uFiKqJsQbhyWuBzdcpz9EM5i27hvBnUKnDT1YpNEOEK9RfW9m+DH6Zlx6lqpGpV
XkCMmG6Ra5LdGGC3m1Xe9v0ixuuEmLyaWJhcQymF5NH0vOV98WItBMaK59t/LoOOGvcehavcguh/
r4EebNqpNwwPBLjKJPn1yGOsPBfsvfsDFS+fwRRHqyVfv/xrL6w4ypxwWzE4wL/WHZK6aS929brd
vkOoCEneYbpaTmE6ZMLt1e/+qYuPpgoenkJFJp2AmqfuSCt9dvFXNd+Ub62IxpBWi895Q611qtXF
DyoS0syp2WJ4sA1/i5aRGIXraQ/vQagO0Gv3vupOtIiQu53mhntZnh8M7zn8fwlWyIDjBLg/rFi6
EsaBhgP3reINC/4LOtzZyaeB5JcRE+n2S6gW+lSkkoY0bKRzH4EWrMWw7stQzhJgeDetZqJWwWhl
Uzmu9TfPpF8MnnJPf8aFL0s+Qq7vDMqg+c1jwqwHVlZPGVq4pTqjo5p8eAvqGhb5Ign7biVU1Ftc
NnLqy/5Rl06uW1J9y5w3Lpf/Oat/bEnsTzWuPDEE8n/8zLWhX+UqTgPv8I/E3iXfNhbOUXuKHktk
P3OcmmZ8cP0RyemnWXrXuRqW+HImtbTV8P6EGz9R/yzbUa2HjPYXayR+HLIkkcX2jBf8Lw86+GMA
DQ6NjeOXdo4BqIxvMyhvXeYxWpZkfUfTNeYsb+1qISflqDzbjmdUYHjh6MoFygHcCs5VZgjcPwOC
TFFMZd/uz+NsVlIJruKwfGKkbYrrPwFAA6GcEAVqjf5CRrmCs7gE86tu8s8hTcdF2/kyrIE34+9i
+y+Ukil8LWMaf7/Fnro12RT5tE52q0JcJ98rqxCGIq0F63ZQ09CqUTbyvwwq87uMHpUc2avQa6VB
6sPlWtldTpicgoQhK8/Vg05WzYdn3Eboi4wSfBQ6S+q3xdQhhb3if4o2Nlp+DK1L+jUZf/dKH7kV
BoljaOiHvRhaVrlHrNp3a1nxRGBO0CwG4bNI5l9RwPq1G+NtoogPEGDOaDuqAyaPXciAxFM8qP+p
FboTDOfzLE4Q47TuhQ32cJxE8fOqTcYQJKPZEHbZ2gIcliuFDUH/Kb0oU8KVq3xzV4rghV3/aMUA
FGBqxC00BlCQo/dHE1BNwQg9VrNTcgNb4JMp//7iKs/g0N4NOuPdQfRJaQSZmzB7CtGXiJelTw0A
Aja/aj4wPArS8msBkW3D3LHadmtTPT5sHRF6AORYJq9uIlVVgMhH1XZJnUsnaJuQZaVdK4FaZME/
LScWhzEwga3d2onxgzGu4D5NUWnQyUDAPG7t3TMGMdgP27Kq0qVYfmFX6MTenumMdtsEYqsOYiUP
61jIVxf/1eXLtQJVRVmh7zp4RlRjZV5hvsLTAwf9VNYm2nopM1MXVOdc5gwBRZdqB7Qfhouz5UBV
Dp1DeV+BOJweiu4WLXWZi+empZX/Gq3dNMFZ4PQjjhOweGqbFpw9Dz2RUWqDTPh7B8bWZs8nHZUL
yFueIuzFuu4PzQyRlDz8AoAC5VGKeLc1im/2JuLfYI6PKQjvY765RynOXZDrQgGKLJFEVXClFads
9oRgiflbCh7maOseIruai1bzNt6aHAkk0SwP+pJAEQl7GNWHTOFiarZf8jV2DYd6hOSsIzxCG11D
bSgzA0skZbrJ3jkCLBMZqWWrL7sKqknQuhtIvE0759aIUY4L3a/C+w533OMDoBXMV3S/pjLl5GO6
V9RxGkRivPJeYoCR+fugx923Dj4Zy0dvnxYCXgFBEUapDMgEq/ELTvV4R7niKm2ni/Kp1DlxeMJq
PwqMk3L9uy/7yEG1yKJY4btv5QdkPQm4BMPYjF4jvzxG7IcjVVoTG1N/0OV+dopN6ZM1gnfueuH1
OmST7Hwov1e48+ctN9CuzvHjTujqreTlQZ0bgT6QUgspflc5t63soDV05hlDCFmBDaaDIAeDEhWZ
C7779OwdTcMz67RVSEekoqndO3YpCmpFGRoMsjFxqG1ijclc+15j3aMkhtpraS8u0FiTmRIQM/Ka
Y2lJgQvs44UUiCaQ4jwf73iELPo7fIHj7BRyTadXv6G3EJ94nACDXM+as9y0UB2H/hNoZqXO3rIc
qOcgP6PbswkVv3sjSwUqOnS5x6IXNudD9jcXaCOVQXGdxqg35MlPDii7Ab3VG2i7QBRPD8dzPuKl
cRdg6A/c+hpgPN/ghhSs2esUDjBCqD5j9zazmaO81dJi88l1wInjmdvhC8Fdf0T/3SrzGTkELqQf
jaxdHfkT3+LBxDNHIaqdS0K4BQXFCLu0InmLXuOMJsOgUqqc5Hx8JalM96viEuMsZnjmeI0L7tYQ
gLlBtES7hNV6qfcmFdglmGu+AXYIYZwdJEHP1EU2hB5CMVuXmzsRp/YT62aS79Slzoxw1sjqRLX2
NyQhmqLF9AQLy8usXHdOYWYUWuSH3J9SyXanDFkDCm19VChNHV2l1+p1Z2YgxbrklWRhafE/mEhb
NpEoCx6IkiKMV6BCLNwOSQwcK8St6/To59C5o7XYCY93SrKpSvud8lXzOh3lrDGcqD8Mrw/xCwfC
JoEmqvimBgGWkFpIcGGC/NOnFlxd+BgKpJS8N6A3NHbiLEggk4kTZBeUY+DKAnWMnsiaMESHPofi
fDoUrXk9cOAPZ0aS/i3u6tb2ZhVRbQLrCriwfHd0Z1lVdxtPCy0AhtCPoqrTfQd0Ya7oPrMjHtj2
TvXKcLahHvipIHbWzeulN5Im+pJDDECMIZUTfhu4uOddjsyzk13l23ktFwaqPQKlZpHluVj4suqk
omvcYwBy799AfzAfBHYg9cQr+H9B6KI7G8t46Ptidq3rvNT5p/5VlpfEBYwmMg5e+6S7GIHkjCxZ
tBWrJ1E0Fm8R3FtbXSQ5lqz40a9b9VG09lNDUnuL2qywdf6Q76cBoigVUMHryConWsdjgxJns2ep
WZFyvgON57cHQmOI0jhYgRX5PH43s8sGWfQEDIhNe8eZbDHMLD+fIvZcvM2m9syE2F2vsLx1HQwW
6FAlk7Sp5MkshoapD2BITp79Dk6B/vCy9J2ftE/HKkqq0E3nNZBchX9/aM5Bsr5WZCkyFugkFDmd
1AaT97o1qjYuACjwSKGK9/dnbBZncwoC443MKELfIXcQ9GE1zJQhLr5+8qAMj7RanUiUVB8bxbu1
xreaW9LIokLxgvQyqsKaI3FczZuvRaFJLH5ZgbKdlG3RLLnXf4LebJlAyGIZWFeF+e2QOZKor2r2
o0B+XAxQtrZc8InGJnQnnP018oQEI88RINECv3V7+dNOOHl2OGJ8ZoFBc9ltroKGdmu89GLjco7x
TIO6EAgpb3PjzVs/kbTbaiYTnu54ZBYw7ndQgviLTaCZ71aJy8GzWXsLpsg2gIKixZfvFPrJwThm
6G4TTc6gw5AuauSK3gk6kKu7iFdr13kFo6eZA0bq8geAWrUAZTlRBICfyazHQz+bhHYcdTBTn9J8
fvd/ljVWB8tdMas5JH/WfcEYOqDyazJntaDlNStMvmWwETuqwuFoNDHFXf2/C+PKElczB1KI4XQb
GK0qTjqVIQ0mEHViEM1XpdLMuofC47An/0adZNlUkuXACDjBMmB+AmoOdFirkZffxcg/yU4pf46F
kfYN0kI0onzsfXqXLjg3/D9guCNF6PjxsSwjlzVxM/RYAZoEBWc/uearhyQtXUvKDiqnWVHl9RPY
y9qqG5HyUJl1fp7XLu9ZoNDVlKlmGhROoTrADNv/VvMI2Nt2Vkh3rg8kisWzL79G4BeZes/DO/qA
A5/KqPIJszc7kfIHA8ctG1JCIx2yphU9AHHPrcioyLbuW7if9m6t3ItgMbRo7XNq0TYaiwYx9Xvg
P+hW8WCmx8QcEpTERnI7O/d/U6+/S7TKlRXPoU+8UHAkvU3SC7Qz3Px5vjXgsyEJzW4PNii3aQVX
unT+wKI6GHZ26wawmBUTQ0I8sEMka9+0zHHQaWoPLapIf+ij/W9d19F5sg89/zh8g5rEDZilTIVW
nn9c9wK4lTvyjr1J5aiQH/vv5CIcUXXNKXlDR7ywkyPfkiLIhqAsDRFRrBIDnpgxsSRkROa+gB22
ApGw88ZkGBdrzqxwFNzMHxs+xEvRzNfsYrGvZ3FvT7aqZA+lGYst4uWdcaHa08V7zLY5sdeM3JgD
Z34xti4rvcSeQIdS11TwihI1zCn2VFbiyeVRVERaWvss+ThEfYW7+YZURc7ybbM2+SpHlUt9RNnu
2Ii/A2XUQSAf7Ooxp409bNZOhuL1Je8/2hNTPe0QPBliBN8l1CiYQWOq76OXhz18b0UPFV3oJlmt
xtl62RwKtcZv1rz1cs1Saz1qSQng00D+UFMyZJS854iSXLChlj7bRMqVse4eKDOzRYEbIVPdHLYT
mg4lLqVIynGLk0JVQWb5sf7zpqMKbXvpfwhBKYj4fT/XeI29JcB40IA1OUnIxN+6GyuzkOMAVmO0
85jE0bWtV43sygTyn0hUJizM2ztMlDgxSy2hsg40odcrL1VoqBCDoqYWWP6qrL3vMePyiAzE9041
3J/Y4dAXIcDZzIJXRCoC8d/vPWhm6JcrZKEbP3Bs9+IBHSDzB5uKxEe8Q9TuXMZppTuo3a6kzh0y
eva6ndpndQC1ifbZwWNBPZDIySsCgJHXGls/XOLFVkcdt5LJIdwlDjNclpghatYslyS4XZMQS5Hw
Gjl9Iyl7y+KA0AEQT4vIRXFVqWKWeT4fURVmzFPMyOQ4Qvei05+nOPxZdjKMPjcojrFjlQwjPXPP
mt7HLSgB/yWK8nCTb3xbUX5XzukTvkdCW0cmn1qEPgnZ3EL6zwbwjF5faEJie6erCQJvbqo5zyUP
UQX0z7aMZRpw/kBwo/p9K7JOPVlFRkMxZ2Gr57LEmEgkVHRBGJrJg+HEPnWE5TTbLPcE2lMHApWC
byw9cMCoDoazsWaPrLgco09jS84EITw3ditFTuYToZ21aQbVd/xkPjzaJ/U1QsX4AgqPUWBvUROR
McKVcXb3B0LHlsHt4B0drobzvmgFGJz2shQW/xW8UKh7HGijIRWfU+pU5JIqfZIJAYbGZBgv2knp
sT0gTVWcoQcaZ675r9iOJny0XkDkVUadsVZP59kVr1gQGT3+ilClqIxY4Mgt/ZR8N0N06vwcLFiM
BBA6EX9UVfCmGH9nHCHePHMk2NbWlAXtCn60czD5hr23IQoE9wm1S6+iYTyqI3LxXnJd4vY09BuD
MNiAJarQ5RvD1I3p0tCY2Fjgp6zYtCiegjDZLoLU8wmNQ8h6utsytASz4QeJwzYcP/sKWw5XbMgC
CmXpgTFkzx7A4t1PD5hKRsh5/Oxo2gVUJwrRzgwF0iOIPVJznZZHC8jFZ5HDqwRAJTZW97E7qSeS
8vAfWKzR5QPB051JKtLt+BnSXnzjko4bnuAVV1p/NE5kk6iRCf3n39zerKBr6YtmBXcZjhNcqC4m
dC7nsp++xXPZmnNLdzeM8PdG58kr6hdI6fYnNnYDuNLoVQl4kR4Gax3UreoBXpWt9MGNyuDR/P1f
7t+1zhFB7AZMYkZZs1hoIDSydX7KD1rIv8o0NvDkVsvAaQGg+bnvpthiavNbeWdhD/HgEVAHee//
DxawZc0gxphBMphC+NzqQD7ZJYxfCSsQgaNik8xMQZc/1/bW4/qm3A7Q8geSjzHG0Hpr1yTkJ1Sd
JG5XULCQIAenqWUhoCqFXpZvDngCklDAwtqVLUdnUkNxBGC0BF+wAogHpyXv+HWSar+QBfh8oJZn
hzG1YIoCwgJUNQ/EFCwEbVgfc04rCb/wUISMgTHXx4mfLLt6nDhtOTb4bH9HSZdHhIaUPSSvqaA0
rzzpZrJilTL5LxHI3crzwmoKwPxZwk4GsYgZCJ+hZa9FhqDR+FT3AAUD7LgldZqi127v2yu3Fxg8
9vNfdYuKZXRVBL+/59TPna+BS6aYgoPLZMEIpeLOw5gr+2CIScu0/HnimmIAWr8+1cxT6ai9ovIa
CcaHtwc0xlzxlQAVehTTJiSmqZgyshhV679x0p/Delrg1zOy40pTkICpAflpfvQvVsFYj8cuSpx8
MZEEn/X5My7rw+FnWQJLpcnsGfKnvX2lzo9TWPl8qF9xMIiqsu2VPWL8VDHM10mbJXK5bfygSnwM
urznkDmdzLOQNJOrWybVTkuIgoGiKmI5qIMmOv9EtG/cnytHEu1C1BU64DYqUaHFnbF1RnvoAiJ2
n95Q02Bv1T+wJmQE3GazgOqR5Qgz86GWEUO2GGgkErNfIs7Vd2oxP8UVLQySyYRZQYhkOu6qhxbI
UvlyPQfD882rSiOfFjVv3YkRqIT4o0fNHNVDwk55cd0bxh7ev4l3YOmRujqrav8XxTiSas3svChs
BIl+PXC2V8GlUY7Ayd1WjKmX246NSbP1sCabvDIMxiEXCWUV7a6QNdk7uijuy4KLZ1YIeql54N4z
ETb/I5AzfwFpagAtdN5n+NNZk1YjGQZajOez4cGy7qN+WNDFCb4hYHa+Otfiu4iKCdoCaFWc0s7p
eI37vhE6SU1DgGZlVn2c4IeZubjtvi6RCOJqDAV08BgsuY6rd79OCtwwIMSf9iv0y/qP8QoOTDHM
gcKIN0lRKVSjlsdgvTCZbXzpXEbveYFw7Rows9ZJRnW3PcnPsIHY43xHmXZcVMWpflajCeaWP+Aw
pHlk4ICKFgZ38+/lhqsKXDp4cMZB2U1Dq0KQnVLquTIb8uRcR07trf/fvtnGru/apLZWP042s/az
KETSW1qhZjrMI3vdmQw76J0UNwvBxSW4k9ghaSB+pe+qh+rJ6z8KTEeVqsYC3e2CDCnUg0pWQRS3
bjFCuSHvhgMA5Xf5ncQ2DA4LXAWfA4xAuH3fYUKhDCNIiNpb2OoAWtt7E7SBYszN+WHXfcbkjInQ
Eod3z1peatzdsXX9us1jPwr/112y45D+389GuxYAlJHgRT5YLuyhEAGgvNlM94HBI1AKJhER1aWc
BZdhnrFaigW+agYmyR8F9KnLhWVbRKxW8Vg/VCSwavtedN6o74q3Im4rHb/1+oLhErIKTCqOFcfI
6D82GF5UaOv8lYOHXdPnC1WHW6NaN1hco7ieb72XvKOXyT3MbsGuzrCYDUXa2ucNwjL9234jtDOg
O0XaNGe5x2K2+bboskGx46qawVVlW4r9QLRrKgdQEmn9V/eVU3GkxzsFr9fzvVlURQtJghj/s8aw
U3ZcM+AsbzFsKz76ff2z5m2PiY67UgZoh88dcO2p7IIsJrqhI8J/kDGZ+P7iTk1o36w6AS6Aa7ES
xhpVId5iHc0mGWyRpKTULvY/IRH6D/oYeXiYLlKU8rQbhjVCV+7yiNCuS3qzs+YuLvLTSNUSSebP
vXlndV9riDHBDUXgQ7bAIckRx3NTjJ2ZociYG/Gd5xQFRHh1xqoVi/ZDDaSTFY+Tek5NaV/NGXTv
CAsxboCgaNDRZQyLXC897q7jLQjEpktBbsudX2r5GqMy9YeTfLI09nW+7VRTuZVCILKVxE5FjvwF
0vN9MP4iGLlIzf4wYHWHMHCIGC4C4hlIimghzpvqhwRC5nnJk7h0klfGku97jYJ0Rf4VbhqMfW8s
JuEYpE2gz+xw90VwnTJwd+R6o4AQD+a3xGmemDBal1HP1lwiG9whThAjqAiNflnpL/rRoQzgl8Dn
uYfdKTJif76mOjQLrjU5dMPlHi07diSpxFnVIWOThYCZUM2qzmHKaLQx7buDC7zDnwy4kKu+jZ/1
Nd+OCiOfmZpxtwKfRGMrFEJAbGG0DO1/0ZZcP9ybD3/R4LF4WjXZk0K+KwIGApTL5bkgD4FfDNgY
w5tsnsvjXBPKv1tJaGsWylTABac5UnEA3tDTD/n/rQwsP1V3KN/QbB/tI0Sdj2ijyjlXI3MYZumB
wUtv2ejTp/8NCELIdLEekSgTwERHr5ID9mNiiK5QyeR9FYqhusNI31IV1ysGllRhSUw+LQgc0KUq
v5/w5TkPWz4OuYc1NF4qNl6IeZnZ5pY3hZHMxPzdEhZ2qYwOnpFbMYEL3noQaMz43tViqeZI06xO
t1O9h4r7KjzXhY7oEVpNqvfRmIrAOTql6x3mEt+fntpDdhG7URs7whiDDZTCiDAjQG9iC4VBmJrh
IH60csKlGnZeZGCMtQZa0XffvdHrvrfCYwQBaVDX1pmx/k9RG8GueeLnFV+1gdbPOPRdVNAd/HJq
PBNs1J9jOI+SMEwr8jAIfk1+mXKWFt25Zfef5BY+i5mZANnirL7E4O/t6t0yFezP6zl9FCz1Y7i5
OLDhvs0xUczsGBojTjvwIpIcVJsdi2gLx78B7tDOnh+CxGTTnYXGu2HWL+mC+TEg5sKfkJ9dwsqO
uazC+jxLhDHI4KtSZLzr43DwNVn0QRMvBIcNOUvie5Q8lHyomXnmcDTkm0Wfg0QotOUN04lCxEnu
fq2ledcr88mOf0ft5lRzxOkoo+MPGipCxs8gpDL5rhYSuACpK4XPTf2xoVUZzYu+Ke2zkmDUlP/t
F+vj2KpGfRGabpt8o/jjaGeWlsejkUk23sQvhSBVPNR7BotLyeBq91XmpNnbQJa1EjhzqvY3JQPX
MwsR9QTnqoaHCdxkPvplpbz48JGcSX7gXmolIINvSKqLqtzdt28WQGdQDlbn2JkUha68G0M4tNvy
aD0Vn7nHueUBKz/30KUbdqCXfdKGTAiaRioQXleDDvNhBeqtk4+d0OonbNJ3fBudc4mxg5r9VR+D
xwuubAuFkAC2LQoRZRyDonOyeDm7Odhyk0edN1kXOm6BcnSYfxMw9Z4suraQS71hUFO1tYVIH6W6
US9DKO2WdVVoFbBuedYoINy2Cqz2A9sH3ThNyv/nnzC/9LT9jfJNuQSTmmXY0gsU0/60tpK4b6KO
a2Ykfx4fheLgrUnjoCHZdITrD8h7UhJ3aPuuXXr9p3vEwd0Wn4N0oqs/nACyW6KydrdX8JqjV8zy
hzMb4wZg8yXodPF1ahgyJXcclSxKAYnpZDvXMyBaNQs9e0E1e9QJai5YG2vjYPm+dlJmXye1yJjz
+a6p5zGCO7p8EAw8T/lRZSLYW35a6uxYwuN1wijU3HFZlj6/9NgvY7vimX6/xX90ObUKfy0NL39c
nX8biW3j/7EZEMXwd7gXYkpRVSbG0vp7DzqYQl3Fr+HTWy37r4wF9APKcO93lmt6B1KXqVMuoUgq
gWxTIph7O9nf7WXglozjY5SFv84AcCl8yv1V/528Ce6bP7KMDjmRs46mm3UsK2B1fkocu/jHYkSw
XcbNS27rXmaIi9bSXDMg+03YY+xgo+qtGcYyJ34xhYC1LMOPAb5b6tjmVCgm8ck5NMe651zauW80
lVKG9wHsrsZl502NdguByt+3/8GljxuW+QSPGMZQoFJvqtDZXz5bxmbWfGVzVgs4Q1+U6XITWJ7P
5WXtkSFYki9QPWJYpIneDrWfZZC1wXG/vaAxeNd2pDrrhDKRmQyTuDh1Ku+uO+W7ix0wpq0KlCW/
Sgz0WhwYms8aMhu4RWh2uv+BYglqluW6ezZrUfXIGWZ0a8yto9pWWVZ5u2eWqNyPa1MENlanBEKd
AFa9nHM+Hg01h9dcOd6zRUsqGzTlUbHoDYM0TKdQK2ejRjazgSURUnxERxEi01BeZHfsceeATtEn
6ukdIwy4NtpMp5S4l4YxUkA8naDjI+N8BsCAFsTvwr2ogi8EQ5qib+6JsWtElVtB6Z3eR9t8MhZZ
e2nPABIyhx0cU0ZKYEbusI1QdskpnlzaFKdlMCz5QXXNYQ4LC7AkOspMi3gd59XE0Vk4OCdx5AKe
ybSBsfMoCy6LumqyifxGIw3L4fMcfXwoM1G8dsSAo+/ms5hugXjHNeq2vLBc6iLDeMuPfv1EUPf4
pMsKUqDqa15nFKk8eZUunzk9JS6vzksCwTSs0fNOL92Zg57MFJk32lyqbFPeik1bqz3QaUvRw+9j
ZmevFNPcr5y3zzTJKx8E6qm2A0sO2UAB/Eg4tSPD1rc8Lzmfr5jH4v//VRuSHMwHCNUoJ0My6zCF
aM+tuosj1oL9fJMS1ExJWMORiNJbTqJjDRzGC/wuVjP3X8dnJgfPcDdLjhY2aDZlg9fxWQQYZtiS
1y62WD4Z0k8lelevqX0GnLUBZY3gi0Dzd8mc5L7HwsoBGru8Lq+b6PtdRbu75+JRAYTJFze+rg2y
Uae3zyGVThzNEql9504ZXk58lkuCzfWFJAj18wpyZbvBaX+Pe+WXgPc42XeYCvpsGwhKm+dSzT52
WrxNkO4N/FAdSSqo6Ez6lekbLWjf/CW5zFoz/HijI/bkMnBrAtdZU03OQnRXIAmoxxGmv1/P0+Y9
7CkPauOxyUwO4knQxMBozVd+W7EwTK1/WuC1eB6Tfmk/IyU1QWDPi+s10uRH0eqVIFm0DbKeUsy4
dFNy2vEViDY8Gvhy6Tam1dV4RrmypjnN6sMI0mAh+nSx+6iEFzkSE+i6k8Bjs6qBH2s9lJ5cbEdE
tVjkwNUH6Jntm5Ky9pLFVscd24+6ClhYN+4e5ryHTV7MKi2gI5uAp7ymzOqLLcXG70I2N5Q3IBQR
Z8jum63o5yQ2CZFwGA7TVBBx7C1/rJGzRxA5GpEb5Kd4Z/maldRLY1iK/LEuHDfabve+FZaYC5Ky
twOtDtIpVVRreSTUHju7cr2SK66MJrc+FqEMyT1hnU+5TKvZb6bN/8EUJIrxkwZ9+Uz6445X8qaJ
lni2TISR8HtiXJUYX2LiMhSulCi8kgaAcNJEzZGejBrXNifmu2EU2SvCZzGQDZKhQl7fSi/PulJJ
TgGAvEji7JkJAozeTxvFbGn6hB8YQ6ghWLVQYlAyT1sG8FrSXkAzp59BinS3Z63MequlrAupR13g
ozGQvyWNHddhA6STUfDbkQNPp8sV2XgJoSGMWdcO9Cgrsdqs3EeYTjPKTgRVDa1U5aMKhQA4UkFu
SWco9YRXvmSkFFP7vj2FKm7FOzsRubshfJywl8M5zVJ+47IPEe0vF45+EPBdaTvVon7Wic3wYQce
He06DtYGlstX+WkWQMDqkFpb0KMNEGIzghsJfo4sPVXQmlUbJ0KQJj8lu6ZgLwdSBpGd7daPSpNb
oIlhquYx+VrSlMRs0CUUk+eF2tgzQgX9fkW/2jvGtG5rBg80ckPukPNR+Y8OKLbfLEh5gDHh74B7
nwwjkC9skSaMXgGPGkjYjS0Cwj1a3TEQOGLbWIvxLC+VFgCa8/glhzKD8b03SC4XPf8KM4Xy8hSH
tT2mubkI0X1veLzAk4Deh3VWjxxmrPFMbjUUnHJiCDOauLmkkAbAFZ9p7J/M7d7aOwjatvvSw39V
6dcEY8qu7+DZ4maG3dJ8sXvzEzvEsixt/fUPAFi+e3mO0SMxZz3K1KGjtlZypO548cO8Mlc74e+W
W7ou/1tqQVsr+Yj3jgDXAVFK7Htktavv/5knk7iH6xnKOQu7UjkpNZ7318ya4h2KzL3BFYap9VT7
dHhyY0i1HH1bJFFZ3qpxiJSZJGlMMB6TtgouRf8yQaMW+9o0NbYpgehHspjKBZJAIxRPcblwNuut
OVFW0/JTwWG0v8hWa/IpsJxh3dTqy+miL77xdXzm0c9wKNtkRRO4ltYsv99MH6b3GI8CYkht4SAE
nUzDau5R5Z32G3OsTtWvKqDtGOyIBeC55NjN192W9qcWNdYcKiPd7SMfXz2YYlpla2+xGpU7jzFF
D05BNzHZWYjqktd0bFN/0Cr6NSHe9g/0Db95qC46RICA9h78I90/T2gm+a/GWLB1H3Zz+b+zoDhU
xLud73BhOb09tMnNFTATVw+0acPkubJ8HXm73Xedglrp6sWOAbkPuBUpclt70S5QIYE4JdrTKYAl
0GyjodrE4yciQT6cKncSnf6ajRfXdrEccMJDeWIRIqxJ4pSUQAuBiWx7zijSjV2q+pCYGNzAfl8I
TJJy7yVT+YunPhghSnDmgXA48XrGgP4k59AtA+s+VF93MOt448NnAwCGEiHU+53Gna6KTRJ6Qnpu
wA/YV05YQx7F/R7IHv0LVOOOD2fLoJ8QRBWew/FgG6PD9xKOC7fbR/BMjPwZq1XsEVgr0xiRvPoi
cFdBzxehyaqgvzu6nnjA7RbUqWDAFpJ85wzS5EuOsXGpu/7GiMx+AzIl8RQlzco1wmvZou+7xOBH
dYuKWUuoNgwAso1c310ZBPryr6KpDI75V2oeMM0/Au/RSpxcNVaTWWjO5hM2bMdH+UhvvUPoPlc+
vnD7QEvz7mMTnAqizzu011WdtDHzdEwOixhKHfY3Lqd/t2j4ITmmz0s0b+42ttPSFZuiZgM48Bxi
Dgg4yVX3YFpfpMvZmhLalspehfeUrihns+0tTmZdyeG3Pn8rVH9XmDHuqHYnTEdXTapDz95raL3h
kqXhKhhwFLJ8HHdnj22oVHW075fXMcMlZdJLN7ZDc0qfT+eoxKqYlcNSOUiDb+njeinhUJmxTsZy
jL4jhgUgARGeS6clzxaTUWdLzoBYBqRkyHVacYE8aLEUJgTCEsHUJuPMVl0hKJOgGZZV4gU9gi2k
1MvAyNtVc34uvU9Wdndx5nl2GMFUC8evdqaFF/iXD1LU54qMNfmu93auc3yiDJnoSzPxsj3iKcf+
wXcc8DOp6UfcFM+qhfdbRAo/mvHaRmvuePlqfTECHWCfhUx8qOQtxzs0iepIXlKE1f9zmYh87OKB
/0b0ev8wk7zcnMbUnpqmVcjEZxlK2N7ViUrhg7/9ULL3uTzed3EPG89fy3iGZWV8c2KzswkfBqhy
y61QqQeN2AxBYtzPpxZDTTWXouPtEXizMBOePPoY59k1FTDvfPkI2MFrhYELTZbQqBRVi8atZARx
6KGVya91u1R1CyPXF7vk0KNhsOZ7NNt6FUJXF8V271pxInvkHa67VnOONjhxtgC89OfYe9C9vH7a
FcfcmmzcW7G0B0hS1+0Ub7u+uvD9WoAFXV23xtIwYXQyq4OsNpxgQgWQ0omvSXS36VfkAyGvtHbI
UyVmQPhWhzBaeXT2pIP9CwdRImglCjK4Ahd3g/sOWfkxlej3r6BGWVqPhaBurmN2YekpAxBMYdMu
rkO/EAW2rPAudaLzXvL0vlyrZg1OG6zAWDERnp6vyIVeKlbFEC/wG4Hw7j4eVydyAeEO2LHODIxP
rojDoinFrhAohY3h2R+EkqlZa4IztmPUrjdL4zWiSZQeRUXgnm3VEVPfEMx7efUXivr4DaVb+h5v
/dlDXYAD6M17FAivrN0cr5DQpnPL1ESbqxilgcM2cwik6vN8H6nQV082QXnmp+mJsd3qu2jaD1Kw
2WAuZ3uJFe2HmNazOytQ3MAyy8aNIcGWb3T4zBfatpL3ImdpflW1jr1VmgghUFwCq9fIYi3C6Ac9
A/+56n5BpX4vVnoyr3Y5ujfP4duYL50GjEQ16tCdIRKBNDTqNBAn0EGQB2JWwXLWDkaQEZrKFcAP
ZPRbCIk7EZc/pLt7mW5//Qhyrsu31wF94M4jB+l+Mtypu7mLxnUXn51IuVjZNZVHArb3WtxJFSSi
jqwkRbwgs8UIZpkgOttv0iyVtQRd88iLHrJinNwNYk6qsmUD/SmCCCEJE1SMr4epPYJpAnP1Ba03
cAH/fDVOuBtHnHmf8njopkhWv0w9FY28LvLBafc8iZbCyI7ifdOmOt3Z3bc6C1MLMtefsW0AIiUY
4IAR2k8mtK24D3Lf/rJhUlc/4s/32HgtbN3GUl18JvyKdjjO73rUp7Roko2FHBcRm9/6N3lKBwSr
xAP0LTMhq1YWgKkKHoGntSKbnWBU1bxDddw72jlsZkx+my3LYa9/YuYTg24GVUb8+rWr7lRYDlSW
sVtWWa6eSoXVmxxtZqKObJOLdHPtToTvbJXOKWnj7nKzzERgH3aGWhfCN8vtVc1Krm7901/SpG47
OuhDHIjwovkrbReu0J/73K3nC+onmydcaAnqS79kw7uv3SewsZ+4S9lg8nGN87NvYQMmJJ2tZGfm
KkP6eJvEJR4ICjUArD0n0ZUxKbNNE6HnkppHmfUUfnZ8FKmGSFIQ/uCT3zlc4MhLhMz4bcRVW4nW
HBHQUHRvzhUH3y1DnxVL6Qmfx+4wShVc/2QxKo1UaTLMQw9ki12KAP+8o6WVKnmvubAjd8UhB746
z6Jz5WJugoxPDvvzgTPAQVUlNZYHDj55hEs/Y31JFP4i0BwMQF10KQqx+JPPFoCArN9kgBKZQH0i
E3xXVJF6JQd2rDmSoWAi3yPbubwiTy5EXhaLSTVhlW7yKEZRDMvviea0bFlwopwOa4gF1YKpDho6
JwSDUwAdjrNp1/VQG3CAJMrMlWV3QBpZc6PY62D8NvgQeKjg8v7/p6hTR/j99YvC6N0V0uPpb5Ys
ImQGgS3GHwMM/h3TkkKF4hxHRy1iZVb6dS92ll/2e5rHpKLq6oSosvsP7SAxzIp/NkWrj64hBfYu
HyPiSBwQrTW0MesoU5U4AcbXi2gKZDvb6wD3moUNY1u5N0nZywZLBz9mhW8/1KHNBFXrFfYMDkdi
pxKP/x6WDdIykjs9VeXI6c/gjTvRqPHV052anvKEspSJTm2ZJTkYn1k4tUo1EqDrzu8bqcvXKo7+
djM16OXvDcjUB9Jqly+VUhMQLd3t5Y9E0lNmGIvTg3yx+9MyeOUCJtws5wZDsCGLUuJS6fJcL02Q
HFSrjow+duQ337tPeXb3XAuJHw1zt+L0CC2WyXv+w62Q+BJ6bLHR1UBcrvWXfbLyYVdTK4mPOwgl
LhPH9xsoT9TWiCQcDDHBZWhdDlIolIvzdG+ky1Sp4W/I3AKmWBEqS9imaviQzPMOAMR0U69p6aEP
pVXfD5ClQR6cC1okHNlyw65LCYxZlGVafWTV+O8ytXOYzCxdcl9iXaRVPhM5GHFo1CAdaTTkQwgT
z1dM5Osx1K3ayb4lQ2u2KQ3Qa1eQ49+uCaKINzkArQmzrf8MDJK9TqRq2UZ3YZYOsK4umB0mbXq7
xSL8FENzvau2zmuKkk538+zUmaZ6t9FtlstQu+thmzg7L6MFPMhX4wtsHFDuA8mAPmqaZfRJAtEl
n6IXJLBu76Z1d/013w06Ry9lIYUzxJF1OKjUMyeOPIAHFz9Ee6rqUm0US5KUFUYmut9xybnproFM
tefI1cBhnhuLgi+PZwdHAgnw9hbiW9u789pgvbqizhzZiSC5mHQ5Kp3i+cnzePpdOh/Uw8oXr8QF
2g4e+rwImO9MnUvhnpAo+nhhMLwBcQ/SMgglUW4QMKrGIqZiuJuiopIWu6kJKSRRMT235lSe7q4+
9IHfvA287mAbtZl2lKD+z7/Fy/1C+NATBW1KU1FOGgRnW6JGhZKdEOXfJQs6tZqBa1JCoxj5ZEIA
FxiopH5iQcle2uXiHGaEpSv+r3g09DLCslaYgDpybWlX3CGOP805LnApfTq6YubaeQOiaSwv8lzz
rHB2eX/xt5z1+xe10Aq629ySk5R+8x9SbYZGeBNQE2Eez0qEtlvZqFWdOz/xjRUM8Fzm0y/DhWQ7
SYQe1E11oZB2l78y+O7o0Ng8EoagqY/pcbWs92lq8PQv7fsTvWskgEbOV6f98juVUy9q0GtijCJO
9aTtZXGOvKc1gKZOBivl1MW6MakDh6fn+YHeNbPXMSkxE6zxrMuENPnnQfvL/Y0u7dQtVW8GvxmK
Kqo6BeL3eWiCxtYR3J+zrV6cP22yXR7zo8+eRwyaIPod90gRLXr+zzqUHcdGMvKvWw51yteWZMdA
cIHK7H7moLWXSo/jKn/2Qq4Ya1fTuG5KsDtgtPUIez/RwRNrjKSC1f7KJuHUyMkkMV4Dh/49QVgD
I3XSokWtAMTItzm4p/ePkzkmhK1POZUk064q5tYaBcDVBI2YMNTjnPc3FamI7E+OG4f/+jssDXLR
d8i9Wt5jO696WHqQreZzTRhr6zfNPfjWy3YupEQznKOC2SBk64jdQsZ0VSBO8sRGzeKy+TIBDCAh
c6tHWsG+ZXb+PkZpYQG/dCptJz2irE7XOl4ENS2NKLFVb9UbJZYcVcAk7kq94lxZMZ3HLZBUzQg4
bQIycb7wtBKAKim42c7G6wY0PnZ9KhcHL4JOmYHfDzTVaijBMeCFq8QVeskGrBIvEgmS8qt+4Uja
rknhHtCEb9ijfskM49fbTAQkB/8x2fdlyxim12lYLU5riT/9imHjkgz8ig77YeB0kSa0v+LuIsnX
gRqjYiEOM0Ura3e8o5Ehcft29RdKpi0EebdyrXaBlHtkW0TJNpwRljN4Ne00TzMaTKb99UP4oNYI
mvnSh2KbULz/vLy6dd6y1CrM0rqgESX3xrermRWojo4slU4lNrD8Wh9Ts3U6m8fVE9xm9AzCMph/
jhOcDwCMY9Eju26Mpt6gVf8iBArcmGSCDG7mxM2jeSt8sNnV3zP35mywyhXaE34jPTD8QCuBsxwO
E05UGxtoxKKM8blkr4PmesqbIN2nueeNjbPzrXvYCKPt9pEch1segGEQ7EOkHH9G2Yj7VCidU7iU
Sp+QWSQArd39mUwzWjwep06SXkF0/0ea/i9dq4t/+57B9DoZp0mFoy5BSBQmMW2Vi8NSUF56ScsW
qRsQq+s0C+LsCMFjcYqqvsY1TkvpP61tFlPeBDFQ9q9NQsm+0i+xO4kmtMGgY7ZUaB8UYUk4XhYa
V+n3fuyzzmgcBR2kbt0rA0OPVol/uxL36RXqyjP0oZWeMh9ZGlQYzuUSJMV63StU2dWpVrUd1IIf
ozEgG8YTNW5bmRkDV5BZjzXKL2ObQHSNoGCKChn67tJoeMC3VFWint/pUjtsKbYz5fhApkeGt+JX
D+yelW499fNmZhJ7qc0tsegg3OXHRKee3vCuDLjlujlaZ3oCEav45DJ4sPodPQrUn1IM5LVXV0sT
BvNHQtpOOjALQcj1YZCPXJSeiwIJReWpfIOetiGklaH17xSi6zrsq9PFBZfn1k+ESHcwX9m1Dqfw
MQjBSCI9z//HZ4zHL2CCQ4EDwWISEtLpXrm9eZ7cq1AMCVXmFLmotaLAgdoxriIOD7XT38lMpoFc
78L2ePHJUvOFXx/mPOz9108FSwDgWINapf2sPJeqYkdKSj7NIYubHBb7e9l2qaYpOgXcV5Z3fuAa
lwqpNgNYJEj7NBuZfkXqSH85cfQK/oks3jS6Zs83WPsgHsskZta8AvRZFY7atHifh9eegjkWtbos
JJiWHwRPpfB73XEP/AJcQO69TinGmW/zEZWiYcDdX6qatFHE/bMWfY4obUZ6MgyiQMF59tbHzGon
bAipVkJwpsS7noHcPK6gG4kkwOZ2S37U6QETBU9jXV3I1q9F50xdeOEaVpkl0YAyo21w34JRoASE
zM059ViTtf6sJT5qxxRgCy6AgEnIiVST0Cg3pdZElg73/OZHSyw7+5+52vnJ8ZIdN25BVBr1MGf7
gux07TANreBdDq76kYyElSIC9SI0OhAQ+/Kx9dVtZGGH44B7ylETMDe7S8YZdC0v2rLnjqrTHTNr
HrHRn9xKFI3W+KKMMgzQ227LcsmzfLYVXT2ufBdIARpA1wbHSROnmvMyU4gVNMGfT2WTfOfYZlK+
jKPtcP6jPkYYIvOSf6i9qLAdbUn8VUycA7SAv54GWlB1oVcTBfTagT6FDqKHIX7/SsCYszaEvvh2
OmKoIa7fqi0ELz2owza7MUgZC1O4TKqpc0A24wVmejexywHmHov5QMKXtx34QvjQ47N289GzvGlc
QzIrfwOe7yjWltXzbu6TG1QCSyhhNhPSnMHzDinC6hJpILo0lSPUqqi18TbhbExcTd6NkDFfdeGS
Pge34IY6WHiVQ/kGUezC9ceoF4afVAdtKOpVXyvLABFKzhfgZXCy00vxDin7lbqnIyBfe+ahdBTE
IN0YwaN6l+uz1ac7I0NFPwXWg9QGohtjri9jkWBfW7ADuILU8l+TpQgNu3PGv/apczPMeP+ngA+W
7mmjhQf9nkBQMYLPG4fCEct5KJPuTU532c6dh9kVsYCgqFhRmQ2JhToDgl2deLiXYGUU5na20t/t
l/Ixd5aOyCMMO1lT3WaKgI/o3OUJoj8xnj+yoW06W48DDPxNt5BaWau/2EX1owHJMwvtHAQHczj9
R7ia9pmKOaLXUnSPXNJGlA6M10A/ME+YaSloprKFokR/OQLdVvYiq+3pfczugDVJSTcOjbJDXsEb
RovF6mISLznOAE6v8UboSNvmCpjdHmLM3FGyGgA8XXOEPHn/fNLXx12EgjkGQaIlCRO8eCy1ptok
ePwNRVlSyT1XsMHaf7YQZC9qDfw9H/PSN9yq/H/NfTm99WfbrJgVuzd2sUvt4f3Xjgpcnr9u531P
8SDaOWFOkQu4FGKYed7AsAudKH6Vn3ateShK7AOM6LAKPJC7Wz0k1BK3ZmpO6ZuZBMD6+vXg89Jp
ywHvp+UIkDGu/n4qhg7wnV05SzWarCeIGjSLF1PM+BOnodZMJri93sddWw3+Tr5HxK9qKEMzFTAC
dVqHa9YuQ9ZLFax5LUPu/HQhhTGNqZtyxxHfLuq++2vL5gi6jSWleTJNFSy+W6qRDo28fwAhkJ97
Ob/e1ntNsFaOAmXvq64ZC3CaCQwM35QNd2TUnMfqk94cIglIxw4noE8kpxVOEIjoRvj/n1tYfPoq
ZqAWefkDE8/WrH/cN/KFvY1ZGhzlcTq5/q4WWlZgpKjKR5N5BqgVmVy/cdupeCV+qXE6fk0ZIz5V
PvNTdiTYKjFfRpmD0zfhWWKLf06Ukd5opN0X7Ktk8FaFK4K2djvBJ7UUhFS1VQkNvgfqQNp99ZV0
BR5r0mThupdHrGrfUJEM3rBl9+v5reALbw4XiwIu6PPiBubrQkSymACO+ot/K5nIziTKGDn2L7fj
sJ+pvBwnfXVBraJqo533zlzQyB6Az7wn5fksHfE1bRUeiLaVD+7uSG9vhcmzuBYX1abQcpmyZV6h
1Gytpq9FjcVll/0ZHHSjEAiuteBYBu2BVu2npjjHcnbQipItypoO4TK6vXlGBdcTmmNsO4+6EW9t
bawMX3HxMBaoUe2DagDHSwHjXl12mpNUivPezBIM0qo3YFYERCaaRD2zZDKeySkphGXrDyODVJaN
Fo1KrRV86zBw7F3Lp8ztEOExMjT4ff+eCAZfnVbFflBVdSJd6ZuTznCOUqgxdhWZWGvPhOJzAKt4
0AjAeFFSLZ7AFazHnA37xW3tslw928tH88fwYcIEhF3JQZksSsq+mFeBh8iyRbazRj4O5DYwvwRa
Xs36emclnHECMOHvyPnyrMUyoKYVg89Zr0e9wRsbU8YY3JS3anvYKqHTZ5PoYHTppzTNNv6JoMGU
sl2buMJyJ0pbqlOcCCTQgHGWYpKqz44Y9nPeyavRVP0oOkP8CLQcBkk5RXteGNfcLp0QIG1yRp55
RpfbIn/f8g61hylJ0pt+UQh9PBg5bMd/a1atYGnQsyC4Afd0GB+3/vO0q62FGXQpULmbfcxWP5E1
HRxfkVG29Jxl3PuYlFAGdJZr+fMhnv0RpbwjswoxwiPZXGrUxjF0igmt/mLZeNqi6tqq4CCAs764
WMlc8PHrLCpFvfWKPn230ten5GhroiJj1V3BeCadSqXOo5aRE1uNYzRWiCCofHZPlSdjPkIxy+he
yMBAdsTY8P4YKz7t+l967QfmQG2Arg8QV2oB5PWhvLcuXveciVY3aSGM8YaGnrC5PQkW9ETtnlIx
jf9vxbtMEvd/N2kuN5W9IX5TU0sbCTh4R9q8soLmtrSzyM34hqufZZkLtC8IXHrafig21sh+wREL
smID5ewl3lzAAqnEeJpDMAcuwd7pDHTEasu1o+75QQm4czsVd7KWYr9WRaEBMFEvCtElArQX9689
yBd5TDvN4WqbkBCoHpCX4DKtTjcAft+gdQSBNnYZQyWF0fxNf5ZL7qWaPm6r9sarImzl3ynrTY4N
T2jiRgW3oYKNbRLaAeNzUzRzKWB7waVQn1wuUtLB/M2hfWiPBNfFsbX63VKODwYfelb8f+NW0mf7
w+V3aBXZB9Hl1UHAu4ynSHU6COoGPWrbqtg8jYdVx8i+oe7gKn3Byx/N9hGwiE9bi3g1v/Zsy4hY
mC6BC8WejLfyvJnoDC99A1qjSkzomJhqLibC4POOnqXmdAKpl/VYV9YGSPeo/1BAEC4nmBygMy9c
IIa44xLXQ+0CwYtvwyJHl4H0X7CneUP5ZjQdFfoJgkK2CXCyYrr3Obx8kWWDL1V4aL+3GDHgW+y0
8dBldHX5zhGQSGh6Bg23b3yw0AJIyT5uoRAUyv6iAV76mlUcKqHxwS6aJrOW07IPWB7uRe8QVpni
zW1/+Zemwcogzi9ubGfhZ8CxrwCn+p/sxA5/xIT4w5xlmj/aAj9SYVbkZy0TDcgCB5UnrD8IFi6+
kGGiVqYBTOkvynVh76/6+tIvW7c2dlPxu0VA8GJhFdWZezGozZWscpv71XlOp+Zpru8mu5LSvE1g
hpnCgrncZVr9fROgb90WaZ84LU/X0FkDge4FKWlXnmsUQMHnXFCxMHeK6YIG7xgC7lDW+otQbOmJ
ilEqf54CosoHJLw9WUoLG5+L551CD3JWhSirF3WtCL3c7UXIHrS2C5WQv9ZGOgfxjNaAXsmQia1Y
bpulicNngp5v4tmaKdwlkIDXFtsVRpHp/X2A0oz2WjU5jDe9JJ1yC2xTBm7ucHxozrK0tqmFu6rf
x5CW+YhqCwsUOcFaONWc1MGDyei5Lh6c9EdFW3TglW6ENC8XrUOG590Pg/bSYVcp7EzHJQdUFOkA
LsCDMUcXEbBYu6EcWuXs872jzs1DOj1KbAwJT2fBXan1m69Z9zzVxLVe5n64CPIcjHNrWdkm/zKP
IKCwqvMuRtWjTJDIkGHk/EXN7OzlPiLD9vf5+B7hyy6WNKkEgYznrpQXeThXcE6Hw8OeMsG3LwB1
mhw39KN3m/WksI8zqsjtKF61dvI8C7Hw5yNpm2P0GEFK2iokJUUCsGp91squv4kv90Fp3hXgMh9k
epqIMdmMBzs/tyEniuInmvIniPMI4wPOZJgJTHcDiOBc4R7ukKe1lLjrGl99DY6qhU7pW1H6hiA9
OIE2wEURC0KmiNCyP3uJ83g5bkemxBrsk75xnFCvFHVJpA2Qsi9lhGlW0xOclaGNLN2p9i2E0qAq
6Kyc7HpCphiYropRNsdbzQpWSNgaLBK7iC7DOcG77bm423pp0uweta+5AeTMBknYwLX47vwSGJ09
A1E2rlo50SO6jULlP5aCwIc0nJojUMhJQezr7egXpnH3PE+dJL65Xnts0qy8sPr6uHOBBop8qsyO
5m+rCogYiLIe4+VRSLj5d3h53W7NONdr1F4HFwMlXN0C/rEeu2R2LJCWWoMO1a3AwY24pZ/xt9IK
A7DYkUixS+wq2gQBktiT3ovAh3IUFbJim60xXwv6UE+tD78BGrsaOtiv99FiNXFHLxzOvHI0xu0O
o1X2yl3PKfBNnbO0rAS43XCQYpAHu/aMeUa2a2G6I+78/7emqvPHsMrBfUgp3o6/4k3eZKWh/ZIR
M6oR8XglOQssBqyVM6gTf92ODAXBTPVf159UxWM1L+ai97ctl7IxoDlaN67VAsLZvgb5UoR0CglB
qYiMAjsCTVP5QPZpUf9YwWasoBc8kKOI+fUR4yH3BSzCkUIZxD6RWleTR+k9BJf4/2ioZzPDykjn
3NRX8LmgSCiODDVtEU4u/BU9qzErYCtP1993bqOreGrlH0MGIRhfFuLmbRcazCZZ2AGwVl2RlWHC
2Wwb9T4mgfPK5s4pDXyB2/fa/2RfVMdEvjX9Do/aGBl+L/wG/wHAX9qgRleJ0X1YDt9b4HWAXt9d
gCpaPkiTf9LfkXqTNCDRt+IXHFHq/4NhuAAb+KpYokR+IDZyqCMZn45Mpa3eyQ40K8OfsPwqZ87i
0Qnxb0ew3HlmLaf7Oy+9GhUTYhpeAWZ3WU3/EM7tQ8JjpOHDjqN+J2ex63FOfbnoxZKxQ1tsy4yu
TZczrPtdq2975figqBAusi5jVIEpnjuw2E/UhiMDHoiGq8NFvlN5PMegM5HGs8//IYrJKyxnDbc5
TD1AaUoXYSy5e3/6UimisCUI8/yQ3WwjqwQnuTp2xUmvS6rjhvYMHbAJ3nz7snn96V6bt1EgwHMl
lbLN2s0MghT5ERWD4tAM6Ep0W44UytXnutx0wXbwZmI4dZbxjCjhzEgbAlXCawfxtgSeLJ1i1jo/
k9087woROgwMn3GPBWZijggT8zD8VAcMWD+YhkjArWZunKYFyv4SwSWaWmqEoqiVMA37brOE9BsZ
aPipGSADz8y9YWoDAiZ1kDSp+3axjDr5FHszRntCRTD3AIpRQcdbqAU77LA0EPWEALDYnOo8o5JB
CyjwE9y1eOq2QATHToFumsmUdrsvbolFI3uC2EJpU8llQvaYqDMGqWohVBWcMnpnHUw4/2hTFsH9
+s1VB1qFVSPufcN9P9jzifYEiIvindatB5wWu6E44n7/Oe4lGOLiN5stXYLeEkLmZJe9xi4b2eQg
JEg4r+cldFSIDXV6md5gnqm8RxEdyPXrYRpMbslcjoLTvkNokCTQP8eN2Fj0dypKKIM7upu3Ds7e
JIZhpe5rrLCvdjxXidRkuioaA/5yK97s0cLre1BxpdGSB/+9zZaEJ7bxbYqPmMQq77GaD+D3sZfz
P7Rf853FArusNaPMQnIY2hcVfUM66CbTgivmBDkme9Vr8fZw2lE07dWYvRpeiywHxM7pcI9FF73U
AgQmL7GziHg+/1BHIg9guuFjEqBmNq89FB2fXZPKD5A0RaNWTCXLCcIUdGvtcooT8UI0oB5MPXuM
g7KJsz1pgVDoIiS3W2XvNllizZIeoGQvzOOtH7xXZ5v2ynGsWoICa17M/mYkK52wHSV0HdKCrt6l
CBGC1RCtsNn86tsQIRHdjiGdQ/OPQZSIFRXciM8ft/tk2eUekf+D05un2Q1vjcPh/VtnrNJkfa7Z
oMEuBzbiS1hDS0Sy/7UQ/dKHxpeEtcCfp1VQva/JDArSoe+cnD/nY7K4zKOodzKNrntrAXoohI68
LmYAWHAAO8jeQmjdLhArPNYRrbDsojeQ5B2YgAo1obOS3vz9QDmTyy7aSUC/5xtsUEJdOE/K20kg
oX7ZAMhzgFMOwSbI8uZKn/0q7Wk97G8jUdQrwU0H7behFyzaEud2eb/8QUGA5Rnjsg3ECziuCcT8
TiniUSNxpEmJ37xhkegcFeFXM3Wh7S+4bzeDQsGoXE4C9JXNhZyopY6FToZUA65QxsAXWLwAHGuc
GJozr6I5MxyrJeBn3yx4cqKBZ2LIFjRBuSC7PJT4pgAOG25JrIA1LAJu9yZlWyb71IojbBx6VUhw
cmrTGc7xkIbR4aXWcu5PrOQeo8oyz/rHj4ceZ5Zuxg/dZDK5aFhtvwRgfcphzXMHDxLpWo6XYFvA
wMZ4z84wxvK7Ro7vipWQj/VOrbIr1LaaR37Z2D3LTGXXVwIsKx6WzyQtwGITvuJhwml3TTUtNTdd
Vmv7Xxib4Vsl5xvzuV8BFlKiMjFF8K01JGMT9/Lcdb70k0MK2Aisq6pQv8y9gsQWN5Qb3eF43S/h
VTN8UZe6wVk1+o5l5h2JeVH7zV4I7oKiuLjwsWViy8PkhNpNYuuDhBsSOlbF69s44ZchrbBNDPz/
yy0gmCyFbZGcwHkiVM0+1NIZm0SK20fZwBSi7LwK83igMuIqrwCDEgqOrNNYSFE2Rp3Ci2HOAxt1
SXxW3XZId13pexovoSH1TwZsu94NBTZJSMrI+bOL+s6Gl/k3ucBnMiMga1gdHjatb57IfpU84mD7
ionpCHNMk4TyMKjCG7iTifxPMBx9u8gYt96urSHHVUqO2DzG6L3fn63wU3I+YFqK2iVbrv61X6c1
84gISRU5Kgj8J3wx5Wm3j4dJn2k6dwDt6Drxktci0WMHdmKz+B0rhkLmJ29++lwvdh7BlLDVzmuc
laAxsd9ZJpjDJoufT5Ou8R2PD2pSXD1lFHCwUXNWtjY293vZ9FG9gQyMks3C752z0WARex3MG57N
UZxZYgs2+FsmB7deVWb1gN39gYyhzrOCIcPj5UhDqrkz+BORWf9Pt4vho05uaJfhNBW3YeXLbDUD
Kl5cL7/I8UiguKsDcTa5QKi3/F69iviygXI8p2am5i55+XdM7Qum2bbDcOtFlK6PmxUyQdqxrEKx
scePLdocg5jF1e+niwEJ0UDEl/tBQqhVkvKMmyC60cl3OmDUjVkPhSwcC5diWvrGEA205DBS2PtZ
Zk+MjEaAJ4ynWMojW1Mt5AkYbu0UU9gi0Fe25fzGD+vz/Tvp2EaDiWfS6S7BL0cWSc9C8tZQkFUT
7rfvRGFXkhtYB1/S3VPxLDyqLOD+z1TKQf1ru1iiThVRsxpIYCJKdIl57U7v3ybgmKDARZhSMldX
YhUKZyjpXC/LuEl7WI0OGnA0CLyULpaPx+makmmIzLK+YSdTtxedlPh9J3+AQM8P3jo0y2zBl++8
5arybzYsYpHgudO6hPckFLt87FZelVyfV1qgGvTANkgTl0C950XE2Fkn8KJy80TiBgGdsjLlIrpA
TiZbR6Mf7ohsMBI9oARktVI+daqAx28K4JfM7eIP4mugWdr8VVMrYy71ewzHadn/N0mwcDyB7thj
u1sx+HNymgzDZiaL5H9SEVpkReVy/vlmXD71MyVYOBvK7gO5s1xXJWnUmyRA3GMdsmZQktFPKeJW
Zf/PNTlW7R5X26BqJG9gxiR4VzAcv8Vu500I1yQSKaLwJkEAlRLmT7yYJGCV/lgHrdAV3aexxFWM
HtSCHAI1F1aGNQ+OzdDpAswv/3Ac+HqsD3bcAU/5Oharb2BDkqJWVaJfajGl0uje1OZ/j6uXLLfq
kO9jo5MNzE3IHUz7H1C+O/iGbBN4CYy+kIjfBHHBo4EIIbvyAZtJ7UWsLA4b8ltvlxJB9Kbp+T47
bfVxR+gffP05916zSUmpWdTbbD4pTOUynalpR9FfsJGhB71RKNRhePmFVZDHA6+G7OAnRb7ql7PH
ApDczkNNcICqvb6VJQWIdHY9XnbREtw7BV6IVClV+HpX1eO08KFzOKWd+i+KOF3rh+8zS/oYzeKi
IhafDsWmTNqpWZQZE+S7rgta+QmkX4jgvtcLbqyQqzna+AwWTSMN+VzxWYzVYbt1S+Od7/qRrpG7
d2AC6KljQHUm2eKp1JcWYmjJKrFpw8Wvepf6qvMJtWG3R+/6PMe/J0Mn+obj3mg9HIl6sdGHvnH/
1dI0ZgO1cwPkdcjUgiQlgM46CuNiVDiwGly1ascMGI6nDC2MK1qPUCnhbF6Ko11FjeT8sqSpfSDG
f+40gKnyzO9crd+Zd0on+RAPE8TWMWOEa0Wdvm97ppTeFksURVXsRKPiySrHEQ7Z1jW5wD1WReSm
rMRvlRdbvbhqTRRvJDzTS75owiVBE13A7UGD4OI+5QzCuc4cgwu4ra6T0yKp+n7nPr7+BpY9rxD7
3QdVn38CBdd6F4kIApa+8kJhL1BzhJPqf2ZXHiqbRuzqRZgPjJEKzqfPm56m/MeJ+qyku44q4VdD
LYkfSp9tn3WnQ+A+Trf8tDrbaatUJCAQn4qxAxeg1B+Q3+3yLBm1PplZSIAECUMxnytYDXIUakUp
4+Hu1MVWAfKpaXS+GDNJa75tgpHsW72iI1XFHj4wYcAbtHqsQ6jrLBskkibgzTk9GNnygMUKdDvE
o+LMuAJXEvGwrP/ErNjo5kB9COa4BV37CYmi3aOsoxaw2Tu2GVaubO2NPlg3Rp62/qwjucmC4SBv
FVU82bU9XQbqSTuNBFHp98FCYaLaR/Wt+1alsef7Mq5Ug0DRNvhEQObH1k7V/XYZB0G9pnZlfieP
tRp3eDEquQD9U8JjPqqND3XHK4VDpfnelTyWEBxOc1RuTHJk4nBFVBmjfmkJPdhgGk+GokErCC6M
Npq4n53dIOl0vn1vIOI6Ss6YPPwpAcPzjAbUe51lKOHuff+26j1UVgIxnXW8PnI/h5pZ/aCDkTBF
BbOSZNyv2C0m0YZFKu8w4uNffN1NAYAyWCP/PO4smJFsFM+1GWOADqetfNOoPNhRGZ6ZNzdTUyU+
lRCICkb3GpvPnjnMf/Tv6gfLzVcgJrDu/0myYa8ikQgpwSM1Z7b55kmjFWB9Lit/TDyDBN3RpolV
E10RUt9INZTfpxPGIDHMwbD1Lm9Jsx0YaRoXE+nFUbljI5/aUs/rmP7JeAIS1OiFIhHbGMbVavyo
lM/YXrBBt8EoQLZPBw9KcQ7j9uBa1JVEAQyeBeC8/mlKll1NLrMQSXPSj0dueEsqDdmrTtSUVR6x
PZLjc6FPFo6hYzFS66FLV7OUTFmapeNiOEmgWihpHyYhD94n0zXvy9HeS3fgrW+VMYz2mtYNGYM5
e9zTCwr04n+BMBhzLPdUVvMEmtf3xbHedWj+MryyYrrWumHseZId7szCAkzo+d1Iy7dNAK7SBLI6
dwy2dCXH9EsAmxQgYw4y4lgkQ6O+Kcuss4a215+qr3f7RUKG4RQAT8167dy5V8clqtSqP/akNDTH
dqw8d6Bv8cuwkvHFl+eaxvRxWWKStg+9Uxy4qTCHy0qjZQ9avent9LFAg+iz5j2WUyz3VO5XAwdL
JPSqEkLq8sZk6IK+xlII/nHUOQvnoAwZ8ZXc4BcHiSKmimKJuPeXSHdRsItgEsbsm1ayin0kT0AN
OYiwIiN3JWjOxVJXr6cGR07D4CTz/eMXbkfamBSIt6fa0oNBhX3iQaQwwTpO0YesSsyeEbKLUzlF
fn5bbS0QRkeBzX1Kq53L+bHX/qNoeZC7i/Cwdw2oAAzPKJ5f70ibMszPaXwsVtMVFK+FyGFfWOjQ
7oX/xiIcjfX0Kr/84atQPcb2mt0t7hi+95lFlUM60w2UO1kAKiohjrtHlqLqHuF0zqtKqBDShPy+
aUsbm5krdHNJSgm/PG+aZOzQhmqZzgewOESuoQr8wkkyYCiWngvohnClqqVQj07h2OoFW+q8lOvh
xWcvKjX93AL+oLIkc3bhBzPpgixpGQWQkNW8D3cAdoNU2nm4eRoCs6jjhK/l705LMV0K1ks/Ev78
gcPXfdHRMm6oTQP+bqbMVllrplsY/SxaJTnmMvzLg6dCEkbtEkMAvQ4dQ5ks0k58OczXhgO/9xJ2
TbtfyOJALN4p/yNJBEMtOyJbQRFwDM5IYX6HZgaJnHDzWsPZ4Fm0CK6IsCurO2EzgR2lUHiUJYSn
h+rKE1uxJdcmGpRkLbRjOnRh0oq9cojLK3qXQKj4VxZD8NMR/ZDWaxquuA6enMyt9H/hl904MFM9
nrOdyPWLkLqpVoRnjPJ81UySUlB2juuNJBeS6mw0OrZUV0fLt5dutxvjmc1eR45uXj/0j9Q3sFhZ
hgaKyVPYSSc2OPu1Y5vSHNAlPP1NuGpulVjsnzM2eQqfCt7qenhL9LPyhUsTqHri/RXIKdBBqGmZ
HJ1V7OPP92kxFLgcsB28A+A+3jhBe6mtI0BlFx6+H9v0W76rq//OSgTpDbrY8KH5Lmuia9YrDCuX
1EJY7ybnF3pKmQkWpTtxrqzg6wpIiHX4HdQqACeBgUJQreVVD//i3lQ7DNJn9itG9oW/aqLg+FPw
O01PEtk5MlFOVz36B2Nnqmwzh/NfNhSuWlmRdvDT4DAicy4jk+6WPUyEb2hmq5FfOyQCDN/seoC6
s18ltoFOWLsn1dN2Zm6mup6yYd4EdF/z6/6lK7fbtLIeaD7zIQ0MjEkKYlYVoZjd4LwLOMtWscE+
Afe8o6I+MjRirq9FN4u7Be0avFGjjmpUIKU8puGkS/37tu6HYCe1rHnULpTKQdWmz7qcERBqqr+V
zzAk6hDlmJA4XiRUD+kp2B30VkaHVMeWN0YGtcsMP+vP4dq+AwFnmRv1UPjzo0iq2R+8j28zbNAt
xJopkFm6Fc3R8aH9PeE//clC47jSM76H1/iisas6P9kIL6qFjS+nOZIe1kUVbUMnUT8HzbELB+CE
0I6r4tcs3sBO9w2Qw7zh3WJCG0Yho+kESDKIMv/wzExS4W0mcT3OwgHbP2ZyhT28bNwQbqfCx7of
F5eSBPJkn4tRe5xO76onreq+UzUVj7/+aNWb9AAQIVIoYx72KcorRH8v++yEAVP6Uqot9DyFjJms
0In9AG1Zt2VHB0wKatiMBvtKk8EVPX6dntWLPRmyahOzZrSuIJ7fATFO41pXFUQCFXngEHHZSKE8
RyW0VnbeRoiiaMA/cnPCz0yJ5l7c+Qct4i+HLDbCD/y2LGlStFCc1+qZH184kTgAfszVjAWRlPXq
5CLu8UFkEF2gJe7V78RrFfhYl4//wLX43/eS1nSDkUUSv1aEANGjme6mBzafiNn7H1SXTN536BWc
Nu9riRBW/Hu6Him3M20CXxYIkeyeHoSusgry2tlWLJp43L+gF8ZzYr2Hf6H7amAUw3cmcxpc1RjD
RNW64YL88fLj/6cW18opI/Y5zU9vDDhOrzDhJ2vb/HHkP8H2AaKOW/JHEh9jhxccGvHBFoF4cuyP
SheRYxTIYym8es11ZG8NYHojle0BvvW4/6KV4jVEzxuBv+QrO8RggUIWrH4leQYbEqevd4RygV90
NjwEwSqCHIAPwQesDFIRNmPc+KN+SYEoHry1ItZYvlBj24suHlBbA5AQD2du6yZoQe7fmBeQMHri
IJP0S/K+wn/0s0dOdoUIJ4BWhAcQzI6w+plNZ0Lk0Mnaxq9X8cX9ugQJG1adjPJLhnlAEyzQG7WA
PgsGhUqDYZd5NIomyoa7ZlU/RzqxyB5K7WWmF/okKCNtAR051CJyO3AvSbEc2v9fOT3dQOC6Hu2S
giFEx2kEEZnGLThAUQdKkln11XnLWv34gZXQ7uOOPRM7P5837JQIRPaLulIM+JEQUm2XXe7gfH25
eiKby4x93C1TxfB2VwzAbKFSPQUlUbS6Dz3yBCxXiHiS2m8mw6rue66ld5uZPI5aYxEOyQYS7OsH
gywkz19ALZf1+aeMRX5plbFsUnZ3Y55ZlWHAmC7NSL0azsh3qEEGr8JGGo7yApyo91QvIkWz4rBQ
7yG+XjnGunC57tzhZ/LDseHsiN6mtW5riGgZILGjiiIL7MGXSaQJJqIKEd6I9D4zv7YRTXZOT6CH
A1vuZnKEoZoG45FELIuvi5Ww8IfUn2ZBJaLLU1ja9pgYeJdYj0DiVa+dcHSB/B6GlaoLQ6bu/DcF
ZKEOi1nVDs5gOSn/oMrekvF8PlKizqGfWEJS/kcm4zYPi/tkRl9Hw0MXMqVefV718HMRiX64UjGc
rby7TMeD6sTzlPnNKXvbIYKtulvRRY6FSLzycAkzzsKKxxkhCg4dfwHafkm9Zp4ur3ngYKT0MI9X
33pJ4SYC8tuE6T8BTzZEnvBTPgsCGKdsnm61/GFXYFYLEX9MEyaMdAop6Zu2SvLtjd1yxpJchhge
2Dmk68zBRbO4Zy8yh+xv+GASB91CQdVppNmiNo4X17OV5oGllmUmhrn1lcNHKRe+rzItqUMDXp1r
MJjpAEJBFr4EnQZRiThclEWlwpYaT4DpBpSkmSLvkLHIrWdeVX/KjzpHClyMaUSRlXZy+Ug/b8od
zD+xejrugjLErbGRpVq86ZAnndiXolI18UvueQYIV9UnzSTZoJ2P/Wr3sFc5aN4RkZ8MZpHiQQFY
WWGnp6cMl0F7f9lrtNBlyAwro1mzRjviIwf0vEp+s39WG4zCxGTQYIr0PUSeJlSadZZwttbzfm/Z
h4tcG81EWIt63mL6eMuls2a7FJ0jFVM2NXrSSWGOFpi73USp+3FLMCUjcbZuPkzv5lbORFF6nhyj
DYemoxNAhhHw1ZfGqAzT6AdsBFOLPWaKbZB8scVfDInLnuc0Z6ZtSkab02T/RIpiqad4dlMU23An
F0xLKcdK2ewb9aHR/zx4hRn9HJ5fHvzAx5lukT38V6R0t+KKYZA5ANOGwNAZAZIGxwlWES1fPrBa
vcgx4HVf6iJ9BtOaDWhUD2hN+tTD5GmhhN9wxfVnvCtTTLqncSOQPruCatXu/YSppvHVIA4g4Ni4
HRxtDlkTZ68+Ze4qDGonLVzlaJGIfaKUeXIJJ+vNvUpnfEmvgh0CWTylkd8USjtynFiaOoQOJVkH
xc85gum9qoBGMGIhBX3EDaGooF7TbkQ4+CkNk7hYJHAImyp6ADFQo3zs2Xx+WCwwWJQNU78CRKn7
L2wror2egCYoWglYFc+3WtlIYoqiLHEGt/bpazPnKTP22MhNYFcXnYKIgRhfW38NiTFtj5Iso2dK
aHDF7+SSA/Mp0TTcikAdLWlk5gy68EMIqBd0aCUJvVGD6cFlaaCAG4++u4JJzJq8Y/gVwEHgUfN3
mH1hbm/MSTITdOBSvSeYOIk0q7OaRAETHkYgMqvLb0mEuiRp8S+15cw67zMQu7FPcpYvR1dC8pMJ
ftwYh8t/ps252+CJCIb6Ta78CvAgi/m3buKdTmLYkg1D2Oci9HOAZX5sQqO4EKFe5pxebynx7osB
zoWpZGqLYoV4BV3ywX7XC+xVGfp54PoAcysu0Cl9OOiskKsoO3WaXixvg//jNOFkQyZGc5QGdxtT
5ACNA58ECLB3FYZLb17irQ9HaxvftgxvNjG6pntkTFA147FA4X9MlYBiTChabESrhf0GT6fUT5U5
1UI0rnRiIowy16siA8QBrlB1lTRZvxCagVIaNuu1Ax/ekjNbWPoYGiPZ4rzhfuyxXh1/w2XJnVtP
rku7eKsaFB9YI/TJRyrGDfIuqfZZKmTJRv/lWnoXScTMYmo42UvZnaRuPjPsUtFjRTSkepY4/wyi
a9YK4treBjTEgdXJrwarczcBIh6gqFks9CivePwfz25sl3rcJ1eYTzs9Eq6XVXVcNwu2wmL9B7ld
ZkgHm8e+xygUkpDaWP8yvtQqnK4Ugqlcr2nbuRRkbyoOFKYjBFIPe4llxxKfzInwEvrwScdMYmtG
cywu4P/Y00gigvScf+nHIJnil4YXXvP2+wIg/raaRB+49KCLjqu41b3rwzKs6a1m5nXJLdyUikVn
Q5e5lqATXrFpOeCBRYmuyjWm+Oa3JDXCmQh8YHVfhShY8QymjV6dtXmFcop+SB2emUCpHocAQY/t
INaw7tVR+rrEew/FrxlrB0UK8vRbM00V8XV8HZFBcEkjTOGGPrLkXHqG1wN26sdYKEm0NJywriy3
NgGYBI+T2qWDsgKsT/XHsjn7Ql4KYEOBkvzlzS6svNVfl1SWmxD+JrVv6EOXtqXOM1gAveMsQK1Y
sJ7tpT/ICxeLVYEXc1NKGpw6H+KteShDUNmZHCvl8jAainhiaHe9u3C+q7Eis5QOkmzviAlDj9sc
nKFTdDIv/vr8YiAuLge5dLnutphsVRmpAka9UykEpozoQ77No1gkMp/Y6BXHQSQMXYzeq/AT3xFq
huOIdszDZibR9fSO0gsNs6B27jK5+U4qLSO1IZiAB6aEErrN16nAJzbx7Q6LAW0S+vHav6eZdK5+
PvJ338pU6HdnQTtrdgtxkibuaKHPRDoGFw6qjWeynexfBAQG5khau7wKER3UQqA7E+YhUcsBVBfq
fm/9YdXov5Dt1b+TvCd2x0sdkY+d+vEohgOjwK1YO5yjtpMCL8vPb29c6J8hdTAf3NvYmyPy2Hhy
rESySSWSvRvmePH9lib6P6TLYZnnu8k8NrAG4nxDfmuNvsmWjF07P6DjAvJyquXl+RFu8sgrCJg4
hlkJciPQlzWItqhftxK+bReHtXYsU2MOJrNEGRMi+SZ2hH2xwtIKvUWAI6PVPp7U5IVlJ9rb0rM/
b0Os+RTU6uMnWgiKVTV68MJQlhtxzN+CGu+K32yi2mQ+1QvdY990vbwf64n18thCmtwg3GJLcYVB
A1INzpCrsSnsdd0Nt9T4vBZxDqA8RXWjEqpAgfcSLpquEPgIxLlTR4+xd+I27N1R0rY8OohFSozw
WCPISeLVriwlHDOxvN5Ay6UB5JoiafllvWiFByteQlSHxQdqGRojQKZUeA+bXy/fXZTtBKaCnpls
Ntu2N0cGanI0TcIF3ygQuannqIEiUrwJzXycHccNcNpCfwWK9rNvoDY2H8PrUBGGssGers5vvUb9
v01FWXVCzeo4i3hSBQKDXTFrc/nQ8U1/QlgYQhrBInzJft8y5MgTN6e3+pu+EadpeuZe6QI/rz+J
6xa8qOJkl0FjpqhtpRF9hysWB/8xmjyHI0llVAj5bOjDXA9C38zIUneqdY5uqUvrJeWluRev06GO
cXz4LUG/8rGokgG+3tgWzteE109n7GoZvU+3/Z3nGC13gxs4ZbfRbWhuUQC4S0Q1rY8X7V7pKD68
hOihSXqlii3a7gpehApIyGq1MoYAHMFV1pXQqfU02oETienbp5vtzbedblry4gJ8QQ10z1GpYdl6
0E1M0iUaAzVzxWO/NZqt3iNEQhBlFMN7F8LUk4/kOc3LL+lfhAp5NhlvMvc+28JQrxu3L30VcGds
3MwscC3U354zlkiBkMfTjG3N95CIR7z56UBkex+XXRt8yc4gmSqTfnhOCD2QcrkAK+udt0aW3FTG
MomWH22A92yYRq9S1PmJY7qfPgDk3Lsl3rp4dZblyRbbqONZ17sjOuZG+f4xySaMPmEz7WV1tvIG
ULhj6xeXsLsauu90lkUUfItn3H3OpfUBdU4G6ngfiIBP8JWLF7kZ+TeNg+jEqwECXkB5UiF5xJEw
D6+xN3j9WsWL86sP3PLrUM0c7QK4bxoYGJ7HO98SLRsnUz+uftxIeElybPcHFJ5LzIVI5bl4OyhP
fqQenU5mpzMCjBTtMTcnF2b0Ts4qhICrscCLTYicmKDuSKxHC41JDd2ZnqnYGGROifwmyhHFEWCH
3UGnGBFURCEubmYTMV52hvVp1BPFWHktq+uES1/KKSDAARCAFzDNU9cFMS6U034dE+bhuzzZCRdL
ZcnddbC43U50K/85NI2/EEcxd/vwAbKn4YWmFYsJlBDxYPgQu0AzPiH6MVraZIZDdw4P62IyXnnt
d79JdSDWeoXxfOPjzY6ZbcyIB6l01MfXXhKpjRrqlvS0sAIr4QvOSRVZGwIROHfWdNszsH2JJ1sV
DhV8PwBJ4plYvNfltZa/SI5zNjyx5scvroTvaVSK1zn7M4woEVY5zsWtcEuAxAhegA9zX4C/BJof
TlPbn/eLcY3jumwroWa0aQAbLiqGgfh2KTmYibpNDHR9EaDS+YDb1R2wh99yxq+YGTQ55/1UJ9uJ
15aRj7DVZIZvXLL/HKCM8CU8ERxnmAMmDlGDTVLrvE0jAw5uX7Zn0IeoPGmvJkYYPsHbeXt/e8Sw
EoANl9/YypnGDHo4ifU+I0HNMjTTHgIhrzMMffeH4Eocgf/wpdB1GAikDu1uEPVciKQlnpfYWw8Q
xFeT5RPlFknvUNBkQxh4s55Lx2N30p8gkcVAf5vrW/0MG0QsXWK8nn552omHLQ1QOLyZ5HM8wbwB
GRNlzOZqcpLKUr+/53rBZ/EgWwGAlZjsSzeVqhTztDf76CnAUb86pfm7IXZIF9wM4PiF7g698sMO
FsbbQ0JxzTk1qzRHB3qsU61VZg3KDpZ9gIlK7qHQ26uamzY4Vz5MR+GA98kU7XfbbKzdtiMGoIbG
smLjb2k5EbV1yzGnW4AVllhSdPAqggc0k2UdZ9MvfGfrvWErv6TRlgA8BYTVrR8QOKggKyAw7piM
8/RM4XsiFozgEZ20S9m+TXKgbnv90tK8oQisJpseaH1clgSHx7KLmYYJRWu0vcenfKaMKbkX+Z0M
9E1UdXArVc1VEiqrPaw2H87wM0tzFvwuOq0nP9Lo/mb0GIsPfEojcg53opFnBsFex78QafAxtQ+f
Ad7fWu5lmfeE6Ks7ZzOWtOZjBLoJfmcwTlL8zyJ3FB6CmDlflzuJDm3jFmSO16nFzuLAZg76OG8f
yp0ndbWOzBQ6+jSzcAZmn3eUgvy7ikTkoG3htaTXe5wEVHzzrO3ET4E94TS1f29Twq+Z/734SJVR
Qm5NfqApWEtHtrzlkj1GBTAnMcuUAIQt0IEtwpJBS9rGfBLDuZRWaGxYNp24plD2kcPaOQf7Z4Ur
0Xd+H8UJXM8s1hC+4+RxPBQ9gSRPGeWXzihwuec5e6ys0HMX8gkU3fx+tGU9PrnTLcqyseDYSm1Q
GhYVz2eW0YuRlxovZruooi3VSOnfpzxAt5GqF3dlDhDrTtJnA9WpCchYj3UvDNL7cTskXLjoxwsB
4yLOIzmPcpPSFeLN+e5imHTt4XOdlgzs9DVUayj7sg77LQk2K4JGzwKZIxsV/LBYksgbAkRTpMAm
SvaSAqzuWquR5z//WGM7z/7JRfoByNco1wywS6O2cNv91oMrftdWSuo2wroFXWqm5OUglYCwdwah
jBjozsD++nLjx5ozIC2Rz73pV4uXavRNzk2YtM+uH6UMJsAihb9ET5Oj85Ej4zYEZPe/KDWaTYwE
pDDehC/dRQ7/e1tlVxRVIa1PoRujCoEIWurKNRJvorIRoHNm5KjIQ4JnwVOPDI3d6/wXaOdwsZsf
ZbpZ1h0vw81ejcFZnyI+hK7s9t6oAYRqf3hXapvHHSbVVbtsytP6CsscPgcWlRUVw5X2tB1Zi1R7
G87g/La6mwmQQ2dvEe12SvhYsEr/7zgzDuS3+aRLr3qKFmSx6LGfMDGUwTZ2Wx4HHamV3S+mmYR4
h+WOilJ7Y6hEjWpks2ym5Hha2Xo9AtwOn3/0OAVhXiNo4soOQyH3bVjhmnWGhoyHxrawIrURJMwH
D8u2o5z7l+NXdBBgh6uXcDuFyEJIz65jLiGnq8KcARHRxzlbm/xVl1xioYAVD6x9s9mL0HPKboCs
2MDRySLZrmdCfwz3eP+qj2BWvgeFON5ev3eIWH4uPF5fPQHYfV1wZMfjpN81vVg7nKr12ZRlixcR
V5ht1IrXECEoQuLg3BnAIzc4kxR+mp1iaPcqXKRfvz/5xom8gjI8UlZLB72wzbYcGR9iJDeZYFRF
rR4QRHJqFaA7zeLDRw316SbilstN9V7OG/dJbfEWU9bbcCUL9JOW4Egv6pobrGKTUlrhVob/2qSP
XmV5ck6ZNi+eZ+2LOKb7qQY1e9DlgsxGnDKwWQB+7Q7GGbcXkqW56CBsK1CV8dtVjxkKQMdhgONu
JK8644Wm+ougVGwC0cTUpg6gHLtvpT/tVNWBLo/aCxYHwQCRdRvnlyY0bwF0Sndo7ELd/hLZ11ng
b6yBrBW7pRf32HlUAl8VWzbdu/5hRLlcyONoN7XcP2nMrFYY7fKaW6uGfs2aA+Eedgx8chJ/4o+4
ehjeRTifT3OuNImdweQ767qWgWjpYGaXPx5LNi/6FYzW7XfWD0ZI5NTW4D8EHGH8MxkcTKxcL20O
cSMH0SW0d9elPRPVSSonrNlKI0TIA75Fe4rcy4OcLA0dr4Z2RUxH1v0aySXd0tt6RACCKKh0jDbr
OpvDln12Hl5bnTlx1TWy0lEvuargqPbpcT81uzpQ4LR5UQg3p4OzdCK5P0OcvYHYzsAJ9BEefv9F
kvW0MJhJq2xlt07JPhFsToU0k8b71s9wxtENCtltloUu+PJfAWeBZ6hnGqy9zqg4gOHkIvJtLglH
HY8jI2mUYVSCSx6t1mpat5FjY8lj1N3i9KJTWhIE0Srn5noIA6s1r5ck+WRJhGj7EoPPulDtOZs0
/qjV6VHzjDiNaSnvRwZcEZpDr7G5DXz5bsTZ2zl4Y5Gxso53JCLDYsJddwtV4qgyWpMYloE+syIc
CX2wvkeG16sjhtcWsqjschrU4pkVhJAqalXherEveMm68VRIzEfzCP7aOEF30YRKLzLRMYBzriL5
UhZydx7I3u65pDHtjktvLbyRGmMJoacI3nEO+Ct1Zzc+eRrrVszAR1HI6RAq3yhNlKjYN1jQcKTr
hTUZLb5UGWN0Bl7bapx9zsn7BlkJWPXYEz9akKxko9FRMYF/a9hYuxxoPTrvRfDZVEbIi20//ENb
7WXe55NBkOpv4krOgYMOZAKkgB+CrQA0n2pHGiNagS7MYIwq5Qc/jRkLF2odK3G33UvdyBJjwbo/
SzIeTVDYp7RbrUYXexvy8mhfN4N/mOQ4LXZvdZdfOVYicGKHrKI7TlAY0kavv6iCXNWT0jAxHCkV
4U5BACiP+PZbqUXr4y1Ycsv8s2aTJLhzT74/UKOgq8Z6vd7jkAEAX2tcOfBFfnga5qVGLJ3JHKRA
sm3e8t9LDC6Wr5nnP+cUkox1e5hKTTyPymtt3tHgdNcI++PVZ7dV1hcl6rYszI69bjOg8vRC7Iws
2sQ4+aOgKtSmkXJosl+5gGw6og7Z1nt+dPL9liHrGtNnf/T1hZW+OB424MedyDOQhi9xiWQY+blh
uIBdb8Ax/qga/u3QuI6ZnCfQGjsj81MG5g0CEXehIkAbavfGpwH2nQKt9DieQnkmZLpvMLNRQLim
LJqu4Jc7Y5yAMMmZflf7i6U4OjtOoScTZTVeOqnPoAYjh22fGMDBjyITYfsD5ch1rl4Z4R77Be1V
mhDjXGeUkKX1315qPUpzE+/JXv+oQHbXiR/UnlAUq4Tljv5LFRpBLKqZo5dFZJCzOcpva2JuWQ+z
Zw2GTLxAdOGC0wLgw8UfjwASOS054THh685rPF0L7tWga0QSMVCN6mcBaIv0OnPN4MoToCB+hST4
JewHyW4InUHQ6F528HCrGfjnmiDyTkp29Ube0viGxEYw/2U/dO3LK4cLjlCvOghdDihvcmBGEIkv
1JMhdvDdTCIOt+ZFtxjH9FjISWUBMSzeoxxrqjAWDcG8xAM+2lXSJtXOrqTZGDZzi1lAdIKXWfDz
mvsx1EQDVyfpWs1QBpzrDrcXw7AySTsKXCRk/RhDGq4VI8QpU/Zt5A0cvn9pkADmnHeOCj1hDLB1
oHNdtNUS2/ML9gAsrbVRVJVx7onM0nVEo2ZvJIjWfMgA7wjYsupgHamTh5Nb5tdo1ZyDj8qRSWmE
URFRZjagvLEsLs0mxk2gcA/QqbFNLyP7l/8ZiiJipBncrQcTVKZSRwXUDrGulLvDxHbUpCR8suP5
fP6wpy+Rj82zgu0TD1gXdmbTnViXZShKBF+eMlSdKtMsxUBOmFbhr05nnmdzMFUWs1c34QvTYhdr
308fUVaxRyF8GWh9JM7g2hUS3ln8q+IAt1mdufbKtniSWru28d5ursyJfDSyUFdpxvkm3pDuFEpG
+zOnkztGhzXnpawfAFsx5v+9HWMJKE0iRJTlxYwZlRFWAOeC9aGgWNmlbCDLoJfY5M2QV/4Rasqq
kLsUJrxM0Zn+MxgY4VUTwoKPfKow3RWi4+Ojh8KU6KKvJAcRA/UyD0AFmi3tBsb1A+ySp6RjaSj9
9q4U6mCtRXYpfl7PNs5dTc2YZcIrxycxSTN/ACAK7wczngprbNPVzE4v7/+M0FuAOlsgCRvecrDX
FNY5J9y24LbKrOFg+hivA/fMLyJHSBHZu5oGjjcYiatzY71paYcMTC8/slbl82HEdAZ1I5Ut5YXw
Z8TOUnZRDW7BR8iPfMgLHUJPpUwcmpIiBHfk/foDPU4PAiRlHUfB26zZRPj6ud3TTyNY0uik8bAN
g0DOXT+7Tk50Hn86iz8fvxCniyTaxkuNEVmp+d4xU1J51BDcimkNxH0dodD7Osow1wovJY9bfVIa
aARs7uuBD7tyGYlJR/AkEgyorZIYQOg7A8+3V5pyubnc+rgysAt/emrn3oLiM/DqLZ7BTo4lV2mv
C0jfxi6BKQjcl7vfk7gzkYHpKE8iVot0bLx30PGqdE1y5t6UbN3GIv7/JWPJVxYti7zefFZKiuut
LW6tLJKr136lbLZbwW/R/abt2+CBDA7L7ro6ZdtFVsm4sveF29h5M/qxfyw8Lf/KrcW5DxLCAbct
BS19GrGobuUZqhDttMVk0BTAglseCW5pjCWyMVOQqFNch2F1QgytLIHGICE+7zSgsIEz+ZQn0/Md
eRfCJYdVaqFtnLAL6qz84+GEuaoh69lIjT+Nx55zVZRRELhP6kK++iOaxmRIekJhBUugrEvJR63q
qDMLWzJ3h4dx3llK4ZvbcJwxXAALSNIptzlezeLVBDGpwlxRLHjYwJKlacwC6Sb1VGflQifDiynp
QPHbmYDCfyB4e0hexdDl5xkZ8CvGUKCNb7JqsGD0+dDG7NRlD2DPWRD1BbzCibPgoD3R97yodPd8
biJXS6Hqzmf70zBkCcrhgttf3jCRk6Cerv2240T94GO1dAdXOMAJWee1AGAVrOq6MNf7ELssrFXB
4dzC626pSitjiPrjNga+Zmr6uOMdqZYly6kLOwCKGSfNbgrN+f1+nRf58v8v+WT9C2Uf40Z8pTHw
UBhk7sZwrKKN7hxmKnx3418QoePEepk94nSLHGqvgVV6KJ2NSlSp27Diu48m2GLhyCMmAVgJ5+cZ
m5R6CJLdlm7M8hRHkA99rtxhuXEbx1zjnb8cqYueisW5jZrdqkOERJrLOKH7KXjnCfB72zm7fkUv
2e+PCE/H8CRpcf8RGaDxtHrx1CGNY9uC9IhKpqcztyQwZR9UmXruQqFLjsj+j7DxnkHviy4/FSw9
YMpG1XS/OZKjkP+9xwTtRInhEaHvv8YU9lAzPoAJnNxhRwD+hx2+n0OdB8GcTSUWmfv/rxMUXkpL
QwP3MUOilKJFwydOdP0v1HCAUSEXzvRCKRg19/+z0fsEdINc9snG1EUrVCcVq/3DpdvcqUm6dyTH
ZzdibBQHmLOjaKokKh6UcFI7X2avWoC5SnM3G1BQ64rTwYBMcIdjXU0lsvp6uCv45DI5uWQoRZkH
yEoYuO39I+GatMHydOSun30PCm7S48xmhKV7PdHOlxGCfiYBLE2tG1ZdMn4Qa9hzqMpN8ng3XU/0
d/cmM56CAg9SElJFNawXpcnrPLU4dSd8ustrF2+kdm4vcWa3F40vgeqarrXjtQM0Il7WVRYsXBlz
vVNsNgKhdUdJmxk6ajr4GTZCttZoTFJoQ5nMDQmdxGDq5ElF7Wv0V/ukdZXyB4O/mtmBeflp2Gey
19VCO7cUCuKt2lIG7Sv4ylKKfqIALtnn81IrVGNQQqp9rLEkFlVCs9481n9H3jL7NNDePvqy/YN5
u0BPfWB3i3/pquzzR4GabTsuvW0r/S9ZnQshE75jodF34Ozk+VVkVFaFQlNn/rwutRid0U5+0YzV
/X0mQhTwmU6kbmvRgNQLlXCEIv2UZJYyfNZhnpvLayjTLQE8NaivMRxVWYhh7MxA8kxSB3WS5zxi
V9sbeVyn5aEy7eFknCLancMMw4xrFcYHydXCFV/1uozYE3R9aQ99EwOPHGgRhTjnxXt3pHzWKu2G
yLsQZ0vNAVEYBsXhzuc/Lh8qqtgocTA8Z//2qzL0mx5zSOD5x5b1eq74h6mYEEvp11zhRdIwzbmf
WcTv8238r6VXm6P1igxYo3NRrPftt+ZTuFYY8JxpmvcZi/cVk7MExzTWBPssIkAC/SuB9kQOZljN
O/QogEeuq8fjsuoxMATSNDnJsEZL/x9kXZwzaORs3XcdQpM72poXQ7RuDB1MlzNTdtm3HGthAH6R
ETdqrK85eduMsb0kgY+joVJN+s/2iX3mtRq+0izmBIhAdr8WSDW4fc/EeGG5O2K/w3oVdE4UIanb
+KaVeWpS/14DLFTSEDXl3V3ahD12XPWwwTZyK5+srf5F/Wupc/7YWY5FBmv17DkdUUdf4uKiZ57d
b/uyLnRFH4HuaEEz/KZ15T/QYO15LXvo1cZDYRCJHpjUM7U1xiGqK4yQEF7/QJRFpe4yQWS8VHbH
iZqhtNjySM9VUd4p3nYlPfUVKyyDDIO0VVq86/0T5hzkvogiVdEI+TSLo4fp+bvLntP79W6LXh53
Qt18BfDHZbRhBBm+xGvSyZTKHOGSaddUt26avVTIjasJFBd+19tGV20S3KknNbNkR42f9xlBCtvf
ot8qxulT8SK8gDGCaHKRuA+VQRx42zbHyLdEZSYxZE7HF+PYJN9l6ixPSHUd1oy0sVFFqRLNw3qw
ni7Zz/5M8uaOmYxa36GXEI88ai6BETQagZdA7hdP75QdTiJ50UunoXKjGVS++8OdoWeJaGKyuQIJ
ffUUBizWsPSEANVqd6dMNRxAV9hzTSNLXBDELcSx22oOzzEVH309yTiGNXnFPTnBoXohPfK+AhtW
ei/aY5fmAl31zKNnuuHKu/XTt1Az/4JzaUsrWRly/l/3XtDRemOf2CxwuRF992gfS/ehHUuy+A5R
9CBQSnGrywW9VinLCT/fF1wL26tzg/Y+NbFRz1FS7gvLq6/knB0TPGuIEYjeKgwpS74d7CoQbIYJ
DQFcgH4zpPh2RhsZNiG/oGLYpVZegSvsPSbgTuodJO1uEC4vT9bzJPdXywuJtjzkVfKmEBGK0pA4
MMihkDgur4+Wn6ldQ+0siqx3gg0S8YFhyx99MSk4VLSuZ8jucAVeQRGfjRR/oFjdzoNJhRY8jefm
CtsdQaq2SYkdFghFy29K0RINzptZnJ4h/9tR9PSsa+7iMvimmcKOXznb07IgCeAok2EGSujLB1E6
d8v0NVMI+sTgrXVgB4d9TiROfZ3pQioohbb41fA5qYL3YitVU9CmCUXd/t5MpHJb/YuWlHwUThq8
Um+T1JFIfiKsLB7RBI4vxnN2ueKX/Pb5zQ8R6JyCvB/RzByEQ8cn3JuNtaK9B9zfy7c102Mmxic1
HyX/PZ51J1qHE09lT3WAk4PfUtKdzWJDmNcvfgGsWa1phepTvuAjXrZ2atk2xy0SHbWMdYo4aZOM
0JEF2V+MF3pLoICz498wN0O+b6TDIv5yAGM1IBHQqUm0rfni/aGbLEQHBdDvhhHq/zeNF01tUtF2
VFAyV5Dmgv6eMSMxTwhyeOlOnJwq1M8RsO6Re+LhQt/3h1HwRIaxQLBpYuGQ1kmfeBMCFx3xehXG
QvoNMIGOcH3mdJHDTl+kC8Ctd9IbwwXMPQkZiIHTXoUv5hErrO6QNCDiVP1B/HBKXWpPIjOqdFZm
5ksGgrrgJR/jqHaIETWh+RGIDIiXhFi0SIPvIbZDVexi0LMnI/hoP+AT1T0OSUJlVSgjgk1qmqv6
Z2qGEPqdFEIscMqnaZmJ6sQultdhJTIGOPs9SJFzJojWH/zvEriXZcrMkl9CuKPxdP4Bp/Dzh0ZI
E6Nn8ZtqcRbLoIMU31ys5i0/LN+gpuTSg+PYH86cKLJVpb5LG34tbKLK68xFCTIqOHU/XG0gDlJp
O+fPjAu8JbJm5O1Hy6qlMzGowtaxnlWc0CAYz5HsVw+TR1p88CddgiHXvYWNJ6CRZ7Vdsny81ycs
WaQJzo1bchsGaywNtNIZXZFTSFGQfLjoRSAn3eoqruWmyrqzwm++eG87zpv+J+2/TCvh9hxZXhbE
pUPnCQQEQ5RSv2hXC1563TyBNvPqyCMRsfppj/6jZMQ6Ewn6WK7MQNyQ4IQmmDYG8hOjsRdenFQm
1x29Ig6Fjw3ULSWcCKEUkJg+Mjdfrxr2GcNtbyJkZoXq7wpw4s9BFzr5pFg5UYWP87sIeVt4tRfN
Zi0WVE4XIb7pi7dhpvGUh5x/DOYjBU01pn6r7n1jCE0OnmWSOiSItoOE6P7/n6FhZ1stGYQ49Xza
EKHIwc3mAAtaVn9fCRj+76COsLy15OZEjlvnhfmN2972lwgWwmY96OkYN8qvvyC+fOgCXM4r3ueV
qQy94q/HdageKsl5gS2J2i7u8kaGtdjorWCdF8TjfEoJZ0XUk4cAdTy5vSZuzigEaHbB1xrMRwoC
88qD/ZYu289Nxg1RFvn7ezIxYa4w0KiMYYSVruHLL2itET1uw0cImzJBjrwO9Hy2TToFh8dEjbw1
w3aSKsL6rUgiFPAAHXBYqOxxoeXPzRYvyXgjXhs5vWxqXmNacYxnvBhE9rGwWkBhGuGbt0pCowYe
HZhm/H5dADpzJ/c4dXrinqKR0ug3JgCvlXa2d4B+4oJnBle3dZO9ZXlF+Q6ddS3VUrCOVKNu1ViC
47I8R1p1LqLHnrWwCnrKiOAuB7XkXODFDt925NL2VwHjdIEk2CrP9Rfi93nWF7UJoQ3DYP2x7Wju
oVanMViXmjf4cFOqyib4WKLi1XfwcRxi0zw8HKL65mZKPdXBp4MZExAThWfdqFiN/Rii8yB9hZth
F4UIwpeAALlUNZteEljdA2YwdCqI5I8Zalu00bMPg99DPBIWBlmy433QwELUEVIsD+AgxdrKNZQZ
2FNuM56vRFew26PYzvp0gZCsZ6vAdG32bbCpllh1vmS7gJQ5ykAMAvehy588wiYNSaqwdktWlUfW
y0/CIg4UHEnf/TX1Kgdu06p2yYJckkp94Cw6qcPlcg4HEXBasqHx7s2Kw8cQudL0a0mDgBQVcbtf
kK7BxpS3f2qaFx/hdtInBeUHyL7DgeYZRloa6cEIYOwotZOBnyzJ+cuM56IzGev7ul7K1VALCoYW
63wwzBylvwsseEsF4tBv4Kqp684QrwSySrK+/vxZ9xgJqEPH4aJqeRZPonrHrpittUFY9IBoZCfb
zQyQtSRpEUUVOkqN9dpniZf1dIVOVE6W8vewVtj+Y3I6iNmi7Sw1PhcaS7mfvE64KlOaLNduelsh
CWJHQZwbV87JgqVbik+0qv3C6GjFnLira0rr4w8uMEpvV5U+9IyCjWd5XcDWsZ+KphReBTVevOXT
MWFcOiyYp1q+HczMb7grpIa1vUOnDQhTB2pH/Ywqg7ORQq2XE7aeUt53bHmxdVJFyksg0ftPukfW
NZdkBv0b0YyF5XDkij64qlYqHBKUgqLOh54D/xCTiDMp41dSwSKD8lpNe74VNsBQz5/hYrGjJ8bh
/Ap1nL/6hJl5oYeq7u0O9DL+X9rMCQjAwwO5pQhMSaIZ6g+8j9VH1ixdFmaB5N5NJn9Mr4f5qrBe
8i5o7p0j/w9mNnJLBsOAMh4XTAo436X70ArdofOUOkcSDcEZSJ2+a4+uxUReguOZpf+92eikrwzu
59gZVlnwNEH3KXv/vrkPbsSiiAqbkfllLRlHqMq4heDOGXs66BdgQOHZenlbG/MTGnT6ehiIp0Cq
Ho3Xw+cpjLCL7IJqUKRTecruSFC4SwSC7XPcYIH8LBmscq8CyWLPuFHTMSriTabk72GnhRXXDr5S
aofappBU26Obi4B2tBu+TsGSuSOgjgvkdIm3dWn6HGUllOpgDt8pOZdet0IREjEjg/xX+cZCAuRP
0+tfOxCl41gAb3faBASFSq8GpfHhnuvBgtpr+H/dPntEbz3iwG+kwbVSlQMeS5zw2e7X146F9HKt
SYIab+Kn14vXLMgYikxJiHbeRvb/MoQrn5mUXd3a2BdXU8Pv4Zano1lHf/LopS1xyA1cPD9tu1xu
uGPL8mnwgjj01VxdD50i4R/P3IqbSM1Fq+BfsvPbn8Ufbkk79PmwlFAqSdecnmQ4jhp8YDLW5dZ2
NpHJbhTzUE+ekD3mqVXWPysMd3ahnC0+N+pN39KW8PAtBt0vFMSb2nw0YBWRGwHM6rZzhvNyIXzs
RnzU2VD1RNcoFy0O4/wuU42NfmTdfyEvmuVQjCPGnZjglCGTUtLXbpWr4GSTwxGoTdcELs0EN+UM
oMcFL6T/NOmJTGOrEj9pMAHjZK6jmebC3Sq986se/xkHeEPKD62CSN8I7ekBIJUbmXTqR7UAgMsF
4H97KneYD9ubBGOGQ0oC5mmqIrA9PP0rjXbWbAJhhjsd0hea9WZsiXAuVFioKys3apGXYgJ+nFCi
RK3gjRK5LQoL1ojOL2ySlg1BBC9F9LeEtNZswWajweJ2++czcOjBnX4S7dtPRaM46mwMcVkFb5dM
qRlXjEYhZ2JtY+FbNK1uCx902DCG6iNEmUTrWp1bMjILxAug7GZLqlPMlNjK4UQHAkA0tf+5qMf8
LOt4QCRCNz0fMmlCUfoObBUm0k2KzdetJaXzTh2BymPGeHEDiWbbyVG40geCwiCNIVdK4DGGBfYX
8oIyij+tKmLTP5Wgky3MKI7G+56nzWUWS81NDNS75aqYDHIbFyLPf/WvZnrbUfLkyp5dBauuPlHe
AfnM/8gykEgKxynvN0mqzB9uTThMMzaLTltIUiIWDuWSvvKdSeDKxdILiKiaaGJPGt025Qi0LpyV
rOzTYuM745BzuclzZR1pLZN20bmA33HIv9YHUiQPRO+0xcs4Bixx6Vazx45dlt8eLawSOWS6YLEr
JpIUIqVMwrq7nEjjveqWb5m0PX5KAjLabE0wxbIGDcP6H/lw/NuBzUOmetTf2vbehLUGNZdo6b8e
YrTRdj+nPioi626RFt7AeGStKzimM8T7mJKRlmSoUixpTqDBFoYtnfBk1tQaN2H7XjwS5r7KVSIG
lOfbgXfE7NyP1brAjGrq7x3LJhzsfoVwkRk/5DHCVO8P1i8fMODlD8qk5p36954HRNAS2nuSNDEm
z5Pz9nDum3EkDt+82Z56qUCbZT0hTbT40c+km03qcsDKP9Azm0SdiZcsfYj6Svl/zLUFpalxVSyg
wypP/Bbgxbs4MnSS50J4+EqsmayV3DMomt7zi2vIFVCW9T6Fgs5DHLk5ygoT9ZW+vb60ZHVizDgu
td0gNG/nHB9h/nkHA0gi0zjZK+qjQXg1drEFkmp4ZLeEwbPoe6g69XeMhojjTDMlG8GGm8X3bGp7
EzBpwlXZ/jjbBXcmVCjNEGu+/OJlN8Bfb6Qg8jyy1HXcqeQ+hXKapuAS+LCMMGKg/APMUreFmrzp
XFNS80tHEdgJV58456WBNXfSn6XR7BbmgA8BXDlFEFKZCuxqx9gU78vEh8R/8oz16ljFBG2aJDUk
n7U93BQ83W8dlDB1LrX/8BybGni/X2HijOfFtEDuC8C4y+hUkDPMh75pvXjkLP+unkTcA/KMLl4J
tm2rTBAFIup1fTsiMQj8FSdkdkmrxgduLaUMfmnjpp6NOT8olmlM41MG6TbfKHLll2mKldvnZg2c
4aBJGl1Sy0u8pLv0Uuf7+IvjXq2mwngB5c+LErLiDUFUEy6bu/qZUSenKLkXY5GQ8BYMojxFD2jo
7HauKdrGwOGJYRpFsrIO4F3MvOzQuZhEVYWbwfT/ruZB46VA7qOdRgp09Euq6s+Kdf/OB3rF6Iie
XQb1DwPHasLC/6C4kmpubZ6rbhXJ6BpXtfkNAP+d7TYEvp7TTBqLNInfVahR32x2+e6ayACRWqm2
7qZqZZVIkbNvGemlZofaag193wFFUT8yYfq/V+g9qYyk7WEhp8JYtWC/OZDO8MwkRbLhvhDK1vKq
87PG+xon8J5I2mIeSK/50lMnFi8ukerR//DQeVLfdSLPJGhprf/a7uUMoabC2KPayMLJigqsbTBE
KS2zoRrZMHpX6ED2zUnIzzjTElMMdyYoUvQDj2olL18yLLm4+8C77Wfk9C4B+hs1ym0v1sDpnULG
tukGUT7/XRF8ysKtsUvMZdtPqI4bnuBel2lJiZwVi3YF1zv0lA2MRdrbE9/FCEtfZoVVnPkBkpam
sZUF9+T74ndd56hKHhFNn0/rZBT0NU7R9Z+EGTq2Uc4ICnYggo3FUUvzn2qyIwJYlfirprVbzVEa
OA1VtpMz3rNu6ccovJ6ZWegG3oij91uO7LAAd/775PfEUVD05ityUjbUizu6Fgua39jO8GTTcnlf
dlyCr7br2yrneFnGbVczocRDUYyeOnHkRb10ldtQeGvQUkP4ptpoiKwyyUAh/Wc8X6yyGxhv3Ynr
wYf0HHPEpDQjv9p9IBZ1IGG7+Wka/828N+AAHgC+353rCfUxgKeOIAi3eCjYi2XhUHU/hAIulZSL
53NJAHd7cxorNS6ZCKSxTMa2du6QwUguhRK6BeV59palfsN+kmDVqwr1zdTil5ZvSflXeqs8SYbs
3v4fMKWO7qveneHjcwiHDmOyGcEolsH94RMX8zAEfDS6e2M3SXZnZ0lUe6Er45bAx8bEhcv7ksIp
L1uNYMWa1j1kHHYzKIugM6lnFoPqWYL/E9UqOOXXYVHL839y8I42iy327oyRlQR4EFDp8H+rJP+x
tNZgK6wdMb6joPowFN+j3q5QrG7bSyPZnnRhk5FnOKiyR0uS9Vmh3PCRjJdybBptQqx7Ho5Mk+e+
kX2usiq5lsiXHx+MsIupBDixBQCT9xH8MgYmIPqbZ+UQyNV6tL3oUEjgBlBET63h7xx7jOJmOfnH
qZVZFHk/YsO5pcBOPgHWIP3vQSypVZ5kT0y3jBKq99j+YuQN+aus9d/XwMQrGw7ILvAGU0G0E/HI
M7Lute5RuYbpkexE0/8LjLT+Lwd+ZJszFjoEXajO1dRl/4mng78SSoYYE6kg6sY3hB0KHcWXkMI4
X8rTOdFCvjm4HYwnVvVo3rgM/1Nj5u7biIYsYL0EBu9EjyDTpl6DE12Evt+hWmsTaU/qhGieL6KG
tp1d7N3Slj/qsgHtQ9mc3o8lmnGzynzSfWj7MW1L+vFW0y9nRXoETUIEPK4za3/f/ksLoPj22Ee+
QILVvyLRuKCN0uwUcvziygxxSF9zUvpUy77fstHaAFbGciZ/GtARStaHYqtEyZshDgPuefy4C0NB
woEfVuFgczxqGSnQcEjlKdR1MA0baTlAZhoziPM/5gd+s5QVjG9K6B6CjTwOyliQbw9QbVV8jeXr
EI6/DGxN4PTOjxr91jsiEaWOG8S8xkap2AyGow+idT4Bt5iWeTnEJsJ7/o9XlZboVt53Vu7RSQNY
iP7i2SOH032qlqzSY5BPZKnCSb/n5xs8EajpVFwvyuOSNOsj8oC1+k46eTvgLTmizKpTBLC9i5aB
R9l2Bt1u5zQW6tn069k6CdlUIQuXNCg6P0gbqq+fueIG1QWvy7H2X3b76hNZxuWmkt/78dncueLq
dboxDHWyqGzIMR9Nh4PuSwi+3iUYoUyZJ1EfBogIiKm5UTjvbzam+kLVQ0m0Qx5xSNBf8ugExwR0
cCUjk2lEmNum1RcnyKOgcLp+bmjHmdMjoQQYZLuUjAd0823jgyzxmSda47lmvxGURskYpF/fuLPP
8fY5GCKK+m0oVnmIcrfTxYzBC9Qtl20EpjPrRx7vSJb65973ddZ22yg8YAUfbfGzwa3n8zs+hBqs
k/XAjZmm4jTHfPo+qdyWChc6X9to+Sz27DRhI4wO0vQpOX/J84JVJPd0mwRfPUMcYscXB/VE2K/S
Ap8pFQ6UlsdDgpBByDQqLJbtriYz19fhufVdaRPWOGX/ZocNoefjut23UI75HeaAuM3o+4y/NP+0
Kz0wgNEc1HtZ88GQf1gpMPKoYP+IeB7z5WDFds2MdZwvHPx2FG8nRRGzKpkHycgCYgGFLfaqZBkH
CJ0RfnKao2J2OooHZKmgHQJsU7do1hHOBhAglZmxq/QJ5PvjhVza2AidqwohLcKkbjOEBROhaHUP
Fuvxf+UjRDv2mjhLC9oG4PB2wbtH7JdeLzOZoAY3W7a8Ac1lOjPbyBhvlWiBynYV77L2TuTBLBTq
iK4j/X+9Gu1aSc+zuWiPuqtTvZKDf5DNBjAf5ZA75hzmUBuFsD+ShUIDdSdJpDpkXm+RuRCKCCY+
ZKgB8MuBD1HdXy462q1M3L5oYUT8s6iR1toFnvcHVf39AbGIMDppPMmuQcmIyAKHLmLZ8mwzOzgO
WUbWdyvDlmE7EZl3Y5px60dWRPQSXSjJ7UbP7aoMh+Aq4y+VlKC188GPMAW/sZ9gZcg/A+anxtAZ
N6YWuawvFf+WZlTIvD3ET0/RzzOjvRE8bjDHPt4HoqzCtakEHkDuRIwdKk/oywR8HdkmQeLvDaTR
1/VGREOcKqwGEqQ11fPm3DBS6Sx4k+XT6YRvqXjX723MtsvJLzn3cuqccX/YuGI75Ti9crmphwiy
ny8mejlM4iQJf6aQbxZSTFLgI74/bfbWaiEMOwuOZ61QTJNvpOBBKpBASxhVGKyUNNDKyO2vijTU
Isut1xhW2KZXlJgnME33Rse/bZcF0j7WydShApilbZNt3qn17IsSnp+Wlc+CaVbJJUEpVMpyveLI
uqlhmUFNHy+DLndsOzRCKX/oRZ28bEtKGMARKBEyKar7VHP/VEq2IG+hufvf9r8PUUADeo4NaSPZ
km6zrF612dFGaK3z2R3gKZbXw1O89VBMYbikiUGFMulwyEs9LF8v4Nb0ZX7x/rk2xs+V6bfz7qfi
nNHXOYpI+bpfzY16uQFvC76d4BUUbIQzbenV1Su61oqhdd/d+e/VLUMMx6d1XzFHc7db15pgiSP4
F9kLdhz/Apr+uYOxiBBmJjOYFN7FqU5Jm82R9KRTeRGuFub4alb/V+5X3uRwYlxXAlqoMi4LAvo8
QkJcdRyM7w8ep6xCMaqkpkBca0rgs2vz5pRvRCq+huFqEnSloiuKK2cdfHAOBL87ZG2hQcPSgAaS
uAKVC3chhhkgBv+XN88zSuw0Z5BJxacxuwEIw09CkmrOg6G9CBoydI7BK7in+cjJs/zonYj5jQK9
m/MwzKGqL4A3Uq0N8TfxqadJRUBmBFO7zdHoWbZexI845EjLXEjN2XkPNW8TmxwSqWKUzh93J+Pc
6EjuJpekStmisy4mjSVIADEi5HVjXnETsoPF7VTGGpk3fBZnq9PHb9OkpNtmGmLV
`protect end_protected
